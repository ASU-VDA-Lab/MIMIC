module fake_netlist_6_1941_n_1614 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1614);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1614;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_148;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_147;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_145;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_146;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_144;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_143;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_54),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_57),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_77),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_109),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_51),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_86),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_70),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_49),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_4),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_62),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_82),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_29),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_2),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_96),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_8),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_55),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_58),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_18),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_142),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_69),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_92),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_126),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_37),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_44),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_13),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_103),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_23),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_13),
.Y(n_170)
);

BUFx10_ASAP7_75t_L g171 ( 
.A(n_16),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_129),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_101),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_72),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_76),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_115),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_25),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_31),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_40),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_75),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_43),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_27),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_41),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_121),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_136),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_38),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_127),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_123),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_63),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_61),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_122),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_106),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_67),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_47),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_74),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_81),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_113),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_88),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_79),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_44),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_105),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_78),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_120),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_22),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_100),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_25),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_52),
.Y(n_209)
);

BUFx10_ASAP7_75t_L g210 ( 
.A(n_133),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_83),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_59),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_117),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_139),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_18),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_91),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_138),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_21),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_66),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_1),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_68),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_56),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_43),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_108),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_16),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_29),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_73),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_128),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_60),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_141),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_99),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_89),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g233 ( 
.A(n_48),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_36),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_30),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_102),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_125),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_112),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_11),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g240 ( 
.A(n_21),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_132),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_104),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_93),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_22),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_38),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_35),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_35),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_0),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_42),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_116),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_107),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_114),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_4),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_118),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_65),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_7),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_90),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_98),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_41),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_27),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_10),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_85),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_71),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_111),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_46),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_64),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_8),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_50),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_28),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_137),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_94),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_12),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_1),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_24),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_9),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_53),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_11),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_36),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_80),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_140),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_24),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_6),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_31),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_130),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_2),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_97),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_14),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_7),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_9),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_39),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_131),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_253),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_240),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_240),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_240),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_195),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_240),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_240),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_240),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_162),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_240),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_240),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_164),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_253),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_206),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_153),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_171),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_273),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_177),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_181),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_273),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_181),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_177),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_168),
.Y(n_314)
);

INVxp33_ASAP7_75t_SL g315 ( 
.A(n_151),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_172),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_177),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_177),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_174),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_186),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_175),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_187),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_189),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_190),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_227),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_191),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_151),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_177),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_171),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_180),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_192),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_245),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_245),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_169),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_186),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_208),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_223),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_196),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_279),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_226),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_239),
.Y(n_341)
);

BUFx10_ASAP7_75t_L g342 ( 
.A(n_176),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_198),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_246),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_260),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_272),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_199),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_171),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_200),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_278),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_275),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_203),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_154),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_204),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_205),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_154),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_197),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_289),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_247),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_247),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_210),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_278),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_213),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_357),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_309),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_309),
.B(n_211),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_310),
.B(n_210),
.Y(n_367)
);

AND2x4_ASAP7_75t_L g368 ( 
.A(n_313),
.B(n_291),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_313),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_357),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_357),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_317),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_317),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_357),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_318),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_357),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_318),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_328),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_328),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_293),
.Y(n_380)
);

AND2x6_ASAP7_75t_L g381 ( 
.A(n_357),
.B(n_291),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_293),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_294),
.B(n_176),
.Y(n_383)
);

NAND2xp33_ASAP7_75t_L g384 ( 
.A(n_300),
.B(n_155),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_294),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_295),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_295),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_297),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_297),
.B(n_291),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_298),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_296),
.Y(n_391)
);

INVx5_ASAP7_75t_L g392 ( 
.A(n_342),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_298),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_299),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_299),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_305),
.B(n_361),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_327),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_301),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_303),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_301),
.B(n_302),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_302),
.B(n_212),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_314),
.B(n_212),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_332),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_330),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_337),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_332),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_316),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_333),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_310),
.B(n_229),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_337),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_312),
.B(n_229),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_333),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_334),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_334),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_306),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_312),
.B(n_263),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_353),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_319),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_336),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_336),
.Y(n_420)
);

OA22x2_ASAP7_75t_L g421 ( 
.A1(n_359),
.A2(n_263),
.B1(n_221),
.B2(n_182),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_321),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_320),
.B(n_143),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_320),
.B(n_335),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_335),
.B(n_210),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_340),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_340),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_341),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_424),
.B(n_341),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_385),
.Y(n_430)
);

OAI22xp33_ASAP7_75t_L g431 ( 
.A1(n_397),
.A2(n_361),
.B1(n_339),
.B2(n_305),
.Y(n_431)
);

NAND2xp33_ASAP7_75t_L g432 ( 
.A(n_381),
.B(n_197),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_424),
.B(n_322),
.Y(n_433)
);

BUFx10_ASAP7_75t_L g434 ( 
.A(n_399),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_380),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_385),
.Y(n_436)
);

INVx2_ASAP7_75t_SL g437 ( 
.A(n_367),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_380),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_385),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_382),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_424),
.B(n_323),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_382),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_386),
.Y(n_443)
);

INVx2_ASAP7_75t_SL g444 ( 
.A(n_367),
.Y(n_444)
);

INVx8_ASAP7_75t_L g445 ( 
.A(n_392),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_404),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_424),
.B(n_324),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_402),
.B(n_326),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_389),
.B(n_401),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_387),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_390),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_390),
.Y(n_452)
);

NOR2xp67_ASAP7_75t_L g453 ( 
.A(n_392),
.B(n_331),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_387),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_390),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_423),
.B(n_338),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_393),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_388),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_394),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_393),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_409),
.B(n_292),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_388),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_394),
.Y(n_463)
);

AOI21x1_ASAP7_75t_L g464 ( 
.A1(n_400),
.A2(n_182),
.B(n_163),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_393),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_394),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_393),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_397),
.B(n_327),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_398),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_393),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_395),
.Y(n_471)
);

BUFx4f_ASAP7_75t_L g472 ( 
.A(n_393),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_395),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_364),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_365),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_365),
.Y(n_476)
);

NAND2xp33_ASAP7_75t_L g477 ( 
.A(n_381),
.B(n_197),
.Y(n_477)
);

OA22x2_ASAP7_75t_L g478 ( 
.A1(n_409),
.A2(n_360),
.B1(n_359),
.B2(n_304),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_392),
.B(n_347),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_398),
.Y(n_480)
);

OR2x6_ASAP7_75t_L g481 ( 
.A(n_421),
.B(n_423),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_389),
.B(n_344),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_398),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_412),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_412),
.Y(n_485)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_414),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_412),
.Y(n_487)
);

NAND2x1p5_ASAP7_75t_L g488 ( 
.A(n_389),
.B(n_147),
.Y(n_488)
);

INVx2_ASAP7_75t_SL g489 ( 
.A(n_425),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_412),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_414),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_412),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_407),
.B(n_349),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_400),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_413),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_418),
.B(n_352),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_412),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_413),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_369),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_364),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_421),
.A2(n_401),
.B1(n_389),
.B2(n_409),
.Y(n_501)
);

INVxp33_ASAP7_75t_SL g502 ( 
.A(n_417),
.Y(n_502)
);

NAND3xp33_ASAP7_75t_L g503 ( 
.A(n_384),
.B(n_354),
.C(n_356),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_414),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_422),
.B(n_315),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_391),
.B(n_325),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_369),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_372),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_392),
.B(n_342),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_415),
.B(n_165),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_372),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_364),
.Y(n_512)
);

NAND2xp33_ASAP7_75t_SL g513 ( 
.A(n_425),
.B(n_282),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_370),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_409),
.B(n_363),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_373),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_411),
.B(n_343),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_373),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_414),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_375),
.Y(n_520)
);

OAI22xp33_ASAP7_75t_L g521 ( 
.A1(n_417),
.A2(n_277),
.B1(n_269),
.B2(n_225),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_404),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_419),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_411),
.B(n_355),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_366),
.B(n_292),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_366),
.B(n_307),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_411),
.B(n_392),
.Y(n_527)
);

AND2x6_ASAP7_75t_L g528 ( 
.A(n_401),
.B(n_163),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_419),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_416),
.B(n_329),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_415),
.Y(n_531)
);

AND2x6_ASAP7_75t_L g532 ( 
.A(n_401),
.B(n_221),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_414),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_375),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_377),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_421),
.A2(n_411),
.B1(n_368),
.B2(n_383),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_377),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_416),
.B(n_348),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_414),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_427),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_396),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_420),
.Y(n_542)
);

NAND2xp33_ASAP7_75t_L g543 ( 
.A(n_381),
.B(n_197),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_378),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_420),
.B(n_426),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_426),
.Y(n_546)
);

BUFx4f_ASAP7_75t_L g547 ( 
.A(n_427),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_428),
.B(n_304),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_368),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_392),
.B(n_350),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_392),
.B(n_342),
.Y(n_551)
);

INVx5_ASAP7_75t_L g552 ( 
.A(n_381),
.Y(n_552)
);

NAND3xp33_ASAP7_75t_L g553 ( 
.A(n_383),
.B(n_362),
.C(n_311),
.Y(n_553)
);

BUFx10_ASAP7_75t_L g554 ( 
.A(n_368),
.Y(n_554)
);

AND3x2_ASAP7_75t_L g555 ( 
.A(n_368),
.B(n_217),
.C(n_243),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_378),
.B(n_342),
.Y(n_556)
);

INVxp33_ASAP7_75t_L g557 ( 
.A(n_428),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_379),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_427),
.Y(n_559)
);

NAND3xp33_ASAP7_75t_L g560 ( 
.A(n_427),
.B(n_311),
.C(n_308),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_427),
.Y(n_561)
);

INVxp33_ASAP7_75t_L g562 ( 
.A(n_428),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_379),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_405),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_405),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_427),
.B(n_308),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_405),
.B(n_233),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_405),
.B(n_238),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_405),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_405),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_410),
.B(n_233),
.Y(n_571)
);

INVx1_ASAP7_75t_SL g572 ( 
.A(n_410),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_403),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_403),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_403),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_430),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_494),
.B(n_454),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_456),
.B(n_370),
.Y(n_578)
);

OAI22xp33_ASAP7_75t_L g579 ( 
.A1(n_481),
.A2(n_243),
.B1(n_201),
.B2(n_242),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_SL g580 ( 
.A1(n_448),
.A2(n_290),
.B1(n_233),
.B2(n_278),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_437),
.B(n_143),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_554),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_430),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_545),
.Y(n_584)
);

BUFx5_ASAP7_75t_L g585 ( 
.A(n_528),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_526),
.B(n_144),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_437),
.B(n_144),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_468),
.B(n_360),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_454),
.B(n_370),
.Y(n_589)
);

NAND2xp33_ASAP7_75t_SL g590 ( 
.A(n_468),
.B(n_155),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_458),
.B(n_371),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_530),
.B(n_145),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_538),
.B(n_145),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_458),
.B(n_371),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_462),
.B(n_371),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_436),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_462),
.B(n_374),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_481),
.A2(n_207),
.B1(n_150),
.B2(n_284),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_436),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_444),
.B(n_146),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_545),
.Y(n_601)
);

INVxp67_ASAP7_75t_L g602 ( 
.A(n_446),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_439),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_439),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_475),
.B(n_146),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_549),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_549),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_557),
.B(n_374),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_444),
.B(n_148),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_476),
.B(n_374),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_542),
.B(n_148),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_449),
.B(n_435),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_451),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_451),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_449),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_452),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_557),
.B(n_376),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_434),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_489),
.B(n_149),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_489),
.B(n_149),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_452),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_562),
.B(n_376),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_560),
.B(n_152),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_501),
.A2(n_536),
.B1(n_481),
.B2(n_478),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_522),
.B(n_502),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_455),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_562),
.B(n_376),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_431),
.B(n_152),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_566),
.B(n_438),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_461),
.B(n_156),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_440),
.B(n_159),
.Y(n_631)
);

NOR2xp67_ASAP7_75t_L g632 ( 
.A(n_505),
.B(n_214),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_449),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_495),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_442),
.B(n_406),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_481),
.A2(n_160),
.B1(n_157),
.B2(n_285),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_461),
.B(n_156),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_443),
.B(n_406),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_478),
.A2(n_160),
.B1(n_157),
.B2(n_285),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_450),
.B(n_408),
.Y(n_640)
);

NAND2xp33_ASAP7_75t_L g641 ( 
.A(n_528),
.B(n_219),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_572),
.B(n_158),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_498),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_523),
.Y(n_644)
);

INVx8_ASAP7_75t_L g645 ( 
.A(n_528),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_471),
.B(n_408),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_455),
.Y(n_647)
);

INVxp67_ASAP7_75t_L g648 ( 
.A(n_525),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_525),
.B(n_158),
.Y(n_649)
);

INVxp33_ASAP7_75t_L g650 ( 
.A(n_510),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_548),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_473),
.B(n_173),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_480),
.B(n_408),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_531),
.Y(n_654)
);

NAND3xp33_ASAP7_75t_L g655 ( 
.A(n_553),
.B(n_503),
.C(n_546),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_529),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_482),
.B(n_179),
.Y(n_657)
);

OR2x2_ASAP7_75t_L g658 ( 
.A(n_548),
.B(n_344),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_554),
.Y(n_659)
);

AO22x2_ASAP7_75t_L g660 ( 
.A1(n_541),
.A2(n_216),
.B1(n_193),
.B2(n_194),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_459),
.B(n_381),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_429),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_429),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_513),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_429),
.B(n_345),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_459),
.B(n_381),
.Y(n_666)
);

OAI22xp5_ASAP7_75t_SL g667 ( 
.A1(n_510),
.A2(n_506),
.B1(n_502),
.B2(n_288),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_482),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_434),
.B(n_515),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_463),
.B(n_381),
.Y(n_670)
);

O2A1O1Ixp33_ASAP7_75t_L g671 ( 
.A1(n_432),
.A2(n_477),
.B(n_543),
.C(n_567),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_499),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_499),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_463),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_554),
.Y(n_675)
);

AOI22x1_ASAP7_75t_L g676 ( 
.A1(n_488),
.A2(n_237),
.B1(n_231),
.B2(n_209),
.Y(n_676)
);

NAND2xp33_ASAP7_75t_L g677 ( 
.A(n_528),
.B(n_222),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_507),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_493),
.B(n_161),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_550),
.B(n_258),
.Y(n_680)
);

NOR2x1p5_ASAP7_75t_L g681 ( 
.A(n_556),
.B(n_287),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_568),
.B(n_264),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_569),
.B(n_381),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_466),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_466),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_508),
.Y(n_686)
);

OR2x6_ASAP7_75t_L g687 ( 
.A(n_478),
.B(n_345),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_555),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_433),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_472),
.A2(n_197),
.B(n_255),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_508),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_496),
.B(n_161),
.Y(n_692)
);

BUFx5_ASAP7_75t_L g693 ( 
.A(n_528),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_569),
.B(n_224),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_469),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_511),
.B(n_228),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_511),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_469),
.B(n_255),
.Y(n_698)
);

OR2x6_ASAP7_75t_L g699 ( 
.A(n_517),
.B(n_346),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_540),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_524),
.B(n_286),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_483),
.Y(n_702)
);

NOR2xp67_ASAP7_75t_L g703 ( 
.A(n_509),
.B(n_230),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_528),
.A2(n_255),
.B1(n_288),
.B2(n_287),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_441),
.B(n_286),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_513),
.B(n_232),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_483),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_447),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_516),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_571),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_516),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_518),
.Y(n_712)
);

NOR3xp33_ASAP7_75t_L g713 ( 
.A(n_521),
.B(n_358),
.C(n_351),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_506),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_518),
.B(n_255),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_488),
.B(n_166),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_SL g717 ( 
.A(n_434),
.B(n_236),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_520),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_520),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_534),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_534),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_488),
.B(n_167),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_552),
.B(n_241),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_552),
.B(n_250),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_540),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_535),
.B(n_251),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_535),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_552),
.B(n_252),
.Y(n_728)
);

OR2x6_ASAP7_75t_L g729 ( 
.A(n_479),
.B(n_346),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_537),
.B(n_254),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_544),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_544),
.B(n_257),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_558),
.B(n_351),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_552),
.B(n_262),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_552),
.B(n_265),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_563),
.B(n_266),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_575),
.B(n_268),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_573),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_582),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_633),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_577),
.B(n_532),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_672),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_586),
.A2(n_532),
.B1(n_527),
.B2(n_453),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_673),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_615),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_618),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_592),
.A2(n_532),
.B1(n_561),
.B2(n_559),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_593),
.B(n_532),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_662),
.B(n_358),
.Y(n_749)
);

BUFx12f_ASAP7_75t_L g750 ( 
.A(n_688),
.Y(n_750)
);

NOR2x2_ASAP7_75t_L g751 ( 
.A(n_699),
.B(n_687),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_624),
.A2(n_574),
.B1(n_573),
.B2(n_575),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_629),
.B(n_460),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_585),
.B(n_693),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_585),
.B(n_693),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_719),
.B(n_651),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_678),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_654),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_584),
.B(n_460),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_663),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_582),
.Y(n_761)
);

NAND2xp33_ASAP7_75t_L g762 ( 
.A(n_585),
.B(n_551),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_648),
.B(n_588),
.Y(n_763)
);

OR2x2_ASAP7_75t_SL g764 ( 
.A(n_655),
.B(n_170),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_615),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_668),
.B(n_564),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_601),
.B(n_460),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_686),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_691),
.Y(n_769)
);

OR2x4_ASAP7_75t_L g770 ( 
.A(n_625),
.B(n_178),
.Y(n_770)
);

OR2x6_ASAP7_75t_L g771 ( 
.A(n_687),
.B(n_464),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_606),
.B(n_465),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_611),
.B(n_465),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_697),
.Y(n_774)
);

INVxp67_ASAP7_75t_SL g775 ( 
.A(n_700),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_733),
.Y(n_776)
);

INVx2_ASAP7_75t_SL g777 ( 
.A(n_658),
.Y(n_777)
);

BUFx2_ASAP7_75t_L g778 ( 
.A(n_602),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_709),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_699),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_607),
.B(n_465),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_711),
.Y(n_782)
);

NAND3xp33_ASAP7_75t_SL g783 ( 
.A(n_580),
.B(n_701),
.C(n_705),
.Y(n_783)
);

INVx4_ASAP7_75t_L g784 ( 
.A(n_582),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_712),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_718),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_624),
.A2(n_574),
.B1(n_543),
.B2(n_477),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_L g788 ( 
.A1(n_598),
.A2(n_432),
.B1(n_234),
.B2(n_283),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_720),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_721),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_727),
.Y(n_791)
);

INVx1_ASAP7_75t_SL g792 ( 
.A(n_590),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_665),
.B(n_183),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_659),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_731),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_714),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_634),
.B(n_564),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_605),
.B(n_467),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_687),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_664),
.B(n_467),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_733),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_699),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_612),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_576),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_643),
.B(n_467),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_659),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_644),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_656),
.B(n_470),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_659),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_583),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_635),
.Y(n_811)
);

INVx5_ASAP7_75t_L g812 ( 
.A(n_645),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_578),
.B(n_470),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_635),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_585),
.B(n_547),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_608),
.B(n_470),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_596),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_649),
.B(n_491),
.Y(n_818)
);

BUFx2_ASAP7_75t_L g819 ( 
.A(n_729),
.Y(n_819)
);

AND2x2_ASAP7_75t_SL g820 ( 
.A(n_716),
.B(n_547),
.Y(n_820)
);

OR2x6_ASAP7_75t_L g821 ( 
.A(n_669),
.B(n_464),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_638),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_638),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_689),
.A2(n_472),
.B1(n_504),
.B2(n_561),
.Y(n_824)
);

NAND3xp33_ASAP7_75t_SL g825 ( 
.A(n_679),
.B(n_202),
.C(n_184),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_640),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_681),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_729),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_640),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_599),
.Y(n_830)
);

INVx5_ASAP7_75t_L g831 ( 
.A(n_645),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_729),
.A2(n_519),
.B1(n_491),
.B2(n_559),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_617),
.B(n_504),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_622),
.B(n_519),
.Y(n_834)
);

INVx5_ASAP7_75t_L g835 ( 
.A(n_645),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_675),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_585),
.B(n_693),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_700),
.Y(n_838)
);

NAND2x1p5_ASAP7_75t_L g839 ( 
.A(n_675),
.B(n_486),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_627),
.B(n_533),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_693),
.B(n_457),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_628),
.B(n_533),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_708),
.B(n_565),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_722),
.A2(n_539),
.B1(n_484),
.B2(n_485),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_692),
.B(n_185),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_675),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_646),
.Y(n_847)
);

AND2x2_ASAP7_75t_SL g848 ( 
.A(n_717),
.B(n_539),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_603),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_610),
.B(n_632),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_693),
.B(n_457),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_657),
.B(n_474),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_710),
.B(n_713),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_581),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_693),
.B(n_579),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_630),
.B(n_486),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_604),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_682),
.B(n_474),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_646),
.B(n_694),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_589),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_660),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_613),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_683),
.B(n_457),
.Y(n_863)
);

INVx1_ASAP7_75t_SL g864 ( 
.A(n_667),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_737),
.B(n_474),
.Y(n_865)
);

INVxp67_ASAP7_75t_L g866 ( 
.A(n_637),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_614),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_616),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_636),
.A2(n_188),
.B1(n_215),
.B2(n_218),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_737),
.B(n_500),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_660),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_589),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_587),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_660),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_591),
.Y(n_875)
);

NOR3xp33_ASAP7_75t_SL g876 ( 
.A(n_636),
.B(n_220),
.C(n_235),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_642),
.B(n_486),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_591),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_600),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_700),
.B(n_725),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_704),
.A2(n_244),
.B1(n_248),
.B2(n_249),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_609),
.B(n_256),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_594),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_594),
.Y(n_884)
);

A2O1A1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_671),
.A2(n_259),
.B(n_261),
.C(n_267),
.Y(n_885)
);

NAND3xp33_ASAP7_75t_L g886 ( 
.A(n_619),
.B(n_620),
.C(n_623),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_631),
.B(n_514),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_621),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_706),
.Y(n_889)
);

BUFx2_ASAP7_75t_L g890 ( 
.A(n_696),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_595),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_652),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_595),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_725),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_725),
.B(n_457),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_661),
.B(n_540),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_626),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_650),
.B(n_639),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_597),
.B(n_500),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_647),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_597),
.B(n_512),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_726),
.A2(n_485),
.B1(n_484),
.B2(n_487),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_730),
.B(n_512),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_661),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_732),
.B(n_512),
.Y(n_905)
);

NAND2x1p5_ASAP7_75t_L g906 ( 
.A(n_674),
.B(n_540),
.Y(n_906)
);

BUFx2_ASAP7_75t_L g907 ( 
.A(n_684),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_639),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_666),
.B(n_670),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_685),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_736),
.B(n_570),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_641),
.A2(n_445),
.B(n_677),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_695),
.Y(n_913)
);

OAI21xp5_ASAP7_75t_L g914 ( 
.A1(n_666),
.A2(n_570),
.B(n_565),
.Y(n_914)
);

INVx2_ASAP7_75t_SL g915 ( 
.A(n_715),
.Y(n_915)
);

INVx4_ASAP7_75t_L g916 ( 
.A(n_702),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_783),
.B(n_680),
.Y(n_917)
);

OAI21x1_ASAP7_75t_L g918 ( 
.A1(n_914),
.A2(n_653),
.B(n_670),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_739),
.Y(n_919)
);

NOR3xp33_ASAP7_75t_SL g920 ( 
.A(n_908),
.B(n_274),
.C(n_281),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_746),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_739),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_R g923 ( 
.A(n_796),
.B(n_653),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_803),
.B(n_738),
.Y(n_924)
);

O2A1O1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_825),
.A2(n_715),
.B(n_698),
.C(n_707),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_912),
.A2(n_445),
.B(n_540),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_804),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_777),
.B(n_270),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_811),
.A2(n_676),
.B1(n_698),
.B2(n_703),
.Y(n_929)
);

CKINVDCx6p67_ASAP7_75t_R g930 ( 
.A(n_750),
.Y(n_930)
);

CKINVDCx20_ASAP7_75t_R g931 ( 
.A(n_758),
.Y(n_931)
);

NOR3xp33_ASAP7_75t_SL g932 ( 
.A(n_886),
.B(n_271),
.C(n_276),
.Y(n_932)
);

INVx4_ASAP7_75t_L g933 ( 
.A(n_739),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_807),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_804),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_778),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_793),
.B(n_280),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_763),
.B(n_866),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_814),
.A2(n_487),
.B1(n_490),
.B2(n_492),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_853),
.B(n_492),
.Y(n_940)
);

O2A1O1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_898),
.A2(n_735),
.B(n_734),
.C(n_728),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_794),
.Y(n_942)
);

AND2x2_ASAP7_75t_SL g943 ( 
.A(n_848),
.B(n_497),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_R g944 ( 
.A(n_889),
.B(n_124),
.Y(n_944)
);

OAI21x1_ASAP7_75t_SL g945 ( 
.A1(n_859),
.A2(n_690),
.B(n_490),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_866),
.B(n_723),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_822),
.B(n_724),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_R g948 ( 
.A(n_761),
.B(n_119),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_878),
.B(n_0),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_845),
.B(n_3),
.Y(n_950)
);

OAI21xp33_ASAP7_75t_SL g951 ( 
.A1(n_855),
.A2(n_3),
.B(n_5),
.Y(n_951)
);

INVx2_ASAP7_75t_SL g952 ( 
.A(n_827),
.Y(n_952)
);

INVx3_ASAP7_75t_SL g953 ( 
.A(n_751),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_741),
.A2(n_445),
.B(n_110),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_817),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_884),
.B(n_5),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_884),
.B(n_6),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_876),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_R g959 ( 
.A(n_761),
.B(n_95),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_748),
.A2(n_87),
.B(n_84),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_854),
.A2(n_873),
.B1(n_879),
.B2(n_890),
.Y(n_961)
);

AO21x1_ASAP7_75t_L g962 ( 
.A1(n_855),
.A2(n_10),
.B(n_12),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_823),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_761),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_817),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_892),
.B(n_15),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_761),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_864),
.B(n_17),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_830),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_SL g970 ( 
.A1(n_773),
.A2(n_19),
.B(n_20),
.C(n_23),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_770),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_846),
.B(n_20),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_792),
.B(n_26),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_799),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_770),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_826),
.B(n_26),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_815),
.A2(n_28),
.B(n_30),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_815),
.A2(n_32),
.B(n_33),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_799),
.B(n_32),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_829),
.B(n_33),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_762),
.A2(n_34),
.B(n_37),
.Y(n_981)
);

NAND2xp33_ASAP7_75t_L g982 ( 
.A(n_846),
.B(n_34),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_742),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_754),
.A2(n_39),
.B(n_40),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_847),
.B(n_42),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_756),
.B(n_45),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_SL g987 ( 
.A(n_784),
.B(n_45),
.Y(n_987)
);

OAI22x1_ASAP7_75t_L g988 ( 
.A1(n_861),
.A2(n_874),
.B1(n_871),
.B2(n_780),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_794),
.Y(n_989)
);

OAI21xp33_ASAP7_75t_SL g990 ( 
.A1(n_787),
.A2(n_872),
.B(n_893),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_846),
.B(n_776),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_860),
.B(n_875),
.Y(n_992)
);

NAND3xp33_ASAP7_75t_L g993 ( 
.A(n_876),
.B(n_818),
.C(n_885),
.Y(n_993)
);

NOR3xp33_ASAP7_75t_L g994 ( 
.A(n_819),
.B(n_828),
.C(n_802),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_818),
.A2(n_842),
.B(n_856),
.C(n_877),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_883),
.B(n_891),
.Y(n_996)
);

INVx4_ASAP7_75t_L g997 ( 
.A(n_846),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_787),
.A2(n_861),
.B1(n_874),
.B2(n_871),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_806),
.B(n_809),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_806),
.Y(n_1000)
);

AOI21x1_ASAP7_75t_L g1001 ( 
.A1(n_863),
.A2(n_850),
.B(n_896),
.Y(n_1001)
);

INVx2_ASAP7_75t_SL g1002 ( 
.A(n_749),
.Y(n_1002)
);

NAND3xp33_ASAP7_75t_L g1003 ( 
.A(n_885),
.B(n_842),
.C(n_881),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_764),
.B(n_882),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_754),
.A2(n_837),
.B(n_755),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_848),
.A2(n_776),
.B1(n_740),
.B2(n_760),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_856),
.A2(n_877),
.B(n_773),
.C(n_800),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_755),
.A2(n_837),
.B(n_851),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_784),
.B(n_809),
.Y(n_1009)
);

NAND2x1p5_ASAP7_75t_L g1010 ( 
.A(n_812),
.B(n_831),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_836),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_SL g1012 ( 
.A1(n_841),
.A2(n_851),
.B(n_909),
.C(n_896),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_841),
.A2(n_865),
.B(n_870),
.Y(n_1013)
);

AOI21x1_ASAP7_75t_L g1014 ( 
.A1(n_863),
.A2(n_813),
.B(n_798),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_800),
.A2(n_786),
.B(n_744),
.C(n_785),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_760),
.B(n_907),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_843),
.B(n_753),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_745),
.Y(n_1018)
);

HB1xp67_ASAP7_75t_L g1019 ( 
.A(n_749),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_836),
.B(n_801),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_830),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_843),
.B(n_904),
.Y(n_1022)
);

OAI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_909),
.A2(n_752),
.B(n_899),
.Y(n_1023)
);

AOI221xp5_ASAP7_75t_L g1024 ( 
.A1(n_869),
.A2(n_881),
.B1(n_788),
.B2(n_779),
.C(n_795),
.Y(n_1024)
);

BUFx12f_ASAP7_75t_L g1025 ( 
.A(n_911),
.Y(n_1025)
);

O2A1O1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_757),
.A2(n_782),
.B(n_759),
.C(n_767),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_745),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_821),
.Y(n_1028)
);

AO32x2_ASAP7_75t_L g1029 ( 
.A1(n_824),
.A2(n_915),
.A3(n_916),
.B1(n_821),
.B2(n_771),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_838),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_867),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_765),
.B(n_835),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_838),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_821),
.Y(n_1034)
);

NAND3xp33_ASAP7_75t_L g1035 ( 
.A(n_788),
.B(n_869),
.C(n_832),
.Y(n_1035)
);

O2A1O1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_768),
.A2(n_791),
.B(n_790),
.C(n_769),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_904),
.B(n_820),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_867),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_903),
.A2(n_905),
.B(n_901),
.Y(n_1039)
);

NAND3xp33_ASAP7_75t_SL g1040 ( 
.A(n_743),
.B(n_747),
.C(n_844),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_904),
.B(n_840),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_805),
.A2(n_808),
.B(n_789),
.C(n_774),
.Y(n_1042)
);

HB1xp67_ASAP7_75t_L g1043 ( 
.A(n_797),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_833),
.B(n_834),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_789),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_765),
.B(n_835),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_888),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_810),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_797),
.B(n_775),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_916),
.B(n_913),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_934),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_1003),
.A2(n_752),
.B(n_852),
.Y(n_1052)
);

AO31x2_ASAP7_75t_L g1053 ( 
.A1(n_995),
.A2(n_858),
.A3(n_816),
.B(n_887),
.Y(n_1053)
);

INVx1_ASAP7_75t_SL g1054 ( 
.A(n_931),
.Y(n_1054)
);

OAI22x1_ASAP7_75t_L g1055 ( 
.A1(n_1035),
.A2(n_880),
.B1(n_911),
.B2(n_775),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_SL g1056 ( 
.A1(n_1007),
.A2(n_880),
.B(n_895),
.C(n_772),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_923),
.B(n_1048),
.Y(n_1057)
);

INVx3_ASAP7_75t_SL g1058 ( 
.A(n_921),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_992),
.B(n_868),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_938),
.B(n_913),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_936),
.Y(n_1061)
);

AOI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_1035),
.A2(n_766),
.B1(n_910),
.B2(n_771),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_996),
.B(n_862),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_1004),
.B(n_857),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_1044),
.A2(n_835),
.B(n_812),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_1013),
.A2(n_831),
.B(n_812),
.Y(n_1066)
);

CKINVDCx16_ASAP7_75t_R g1067 ( 
.A(n_944),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_926),
.A2(n_906),
.B(n_781),
.Y(n_1068)
);

AO21x2_ASAP7_75t_L g1069 ( 
.A1(n_1040),
.A2(n_895),
.B(n_902),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_1041),
.A2(n_831),
.B(n_839),
.Y(n_1070)
);

NAND3xp33_ASAP7_75t_L g1071 ( 
.A(n_950),
.B(n_771),
.C(n_766),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_942),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_930),
.Y(n_1073)
);

INVx1_ASAP7_75t_SL g1074 ( 
.A(n_974),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1022),
.B(n_849),
.Y(n_1075)
);

AOI221xp5_ASAP7_75t_L g1076 ( 
.A1(n_968),
.A2(n_897),
.B1(n_900),
.B2(n_888),
.C(n_894),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1016),
.B(n_839),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_R g1078 ( 
.A(n_1028),
.B(n_894),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_946),
.B(n_831),
.Y(n_1079)
);

AO32x2_ASAP7_75t_L g1080 ( 
.A1(n_998),
.A2(n_963),
.A3(n_939),
.B1(n_929),
.B2(n_1029),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_1008),
.A2(n_918),
.B(n_1001),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1024),
.B(n_1017),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_919),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_983),
.Y(n_1084)
);

AO31x2_ASAP7_75t_L g1085 ( 
.A1(n_929),
.A2(n_939),
.A3(n_917),
.B(n_962),
.Y(n_1085)
);

BUFx10_ASAP7_75t_L g1086 ( 
.A(n_973),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_L g1087 ( 
.A1(n_945),
.A2(n_1014),
.B(n_1042),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_925),
.A2(n_954),
.B(n_1023),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_919),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_999),
.B(n_1020),
.Y(n_1090)
);

BUFx2_ASAP7_75t_SL g1091 ( 
.A(n_999),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_1003),
.A2(n_943),
.B1(n_998),
.B2(n_1006),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_993),
.A2(n_990),
.B(n_941),
.C(n_1015),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_1000),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_1023),
.A2(n_1010),
.B(n_1036),
.Y(n_1095)
);

CKINVDCx11_ASAP7_75t_R g1096 ( 
.A(n_953),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1045),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_1010),
.A2(n_1026),
.B(n_960),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1047),
.Y(n_1099)
);

CKINVDCx6p67_ASAP7_75t_R g1100 ( 
.A(n_989),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_1012),
.A2(n_947),
.B(n_1050),
.Y(n_1101)
);

AOI21xp33_ASAP7_75t_L g1102 ( 
.A1(n_993),
.A2(n_970),
.B(n_951),
.Y(n_1102)
);

O2A1O1Ixp5_ASAP7_75t_L g1103 ( 
.A1(n_981),
.A2(n_985),
.B(n_976),
.C(n_980),
.Y(n_1103)
);

OAI22x1_ASAP7_75t_L g1104 ( 
.A1(n_958),
.A2(n_979),
.B1(n_1034),
.B2(n_961),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_1020),
.B(n_1002),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1049),
.A2(n_1037),
.B(n_1032),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_949),
.B(n_957),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_956),
.B(n_937),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_987),
.A2(n_986),
.B1(n_966),
.B2(n_982),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1043),
.B(n_924),
.Y(n_1110)
);

BUFx3_ASAP7_75t_L g1111 ( 
.A(n_1011),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1019),
.B(n_988),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_928),
.B(n_940),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_935),
.B(n_955),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1032),
.A2(n_1046),
.B(n_1018),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_963),
.A2(n_1025),
.B1(n_1038),
.B2(n_1031),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_965),
.B(n_969),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_920),
.B(n_994),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1046),
.A2(n_1027),
.B(n_991),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1009),
.A2(n_987),
.B(n_1021),
.Y(n_1120)
);

O2A1O1Ixp5_ASAP7_75t_L g1121 ( 
.A1(n_984),
.A2(n_977),
.B(n_978),
.C(n_972),
.Y(n_1121)
);

O2A1O1Ixp5_ASAP7_75t_SL g1122 ( 
.A1(n_1029),
.A2(n_932),
.B(n_971),
.C(n_975),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_933),
.A2(n_997),
.B(n_922),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1011),
.B(n_1033),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1011),
.B(n_1033),
.Y(n_1125)
);

INVxp67_ASAP7_75t_SL g1126 ( 
.A(n_919),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1030),
.B(n_1033),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_1030),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_922),
.Y(n_1129)
);

OAI21xp5_ASAP7_75t_SL g1130 ( 
.A1(n_952),
.A2(n_922),
.B(n_964),
.Y(n_1130)
);

AO31x2_ASAP7_75t_L g1131 ( 
.A1(n_1029),
.A2(n_948),
.A3(n_959),
.B(n_964),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_967),
.A2(n_950),
.B(n_917),
.C(n_783),
.Y(n_1132)
);

OR2x6_ASAP7_75t_L g1133 ( 
.A(n_967),
.B(n_1025),
.Y(n_1133)
);

A2O1A1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_967),
.A2(n_950),
.B(n_917),
.C(n_783),
.Y(n_1134)
);

A2O1A1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_950),
.A2(n_917),
.B(n_783),
.C(n_1003),
.Y(n_1135)
);

INVx1_ASAP7_75t_SL g1136 ( 
.A(n_931),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_992),
.B(n_996),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_936),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_992),
.B(n_996),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_992),
.B(n_996),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_927),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_992),
.B(n_996),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_934),
.Y(n_1143)
);

BUFx8_ASAP7_75t_L g1144 ( 
.A(n_1000),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_1032),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_992),
.B(n_996),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_936),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_926),
.A2(n_1005),
.B(n_1008),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_927),
.Y(n_1149)
);

OR2x2_ASAP7_75t_L g1150 ( 
.A(n_936),
.B(n_763),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_SL g1151 ( 
.A1(n_995),
.A2(n_1007),
.B(n_1032),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_926),
.A2(n_1005),
.B(n_1008),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_926),
.A2(n_1005),
.B(n_1008),
.Y(n_1153)
);

AO31x2_ASAP7_75t_L g1154 ( 
.A1(n_995),
.A2(n_1007),
.A3(n_929),
.B(n_939),
.Y(n_1154)
);

AO31x2_ASAP7_75t_L g1155 ( 
.A1(n_995),
.A2(n_1007),
.A3(n_929),
.B(n_939),
.Y(n_1155)
);

OA21x2_ASAP7_75t_L g1156 ( 
.A1(n_995),
.A2(n_1007),
.B(n_1013),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_992),
.B(n_996),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_995),
.A2(n_1007),
.A3(n_929),
.B(n_939),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_992),
.B(n_996),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1003),
.A2(n_995),
.B(n_1007),
.Y(n_1160)
);

OAI22x1_ASAP7_75t_L g1161 ( 
.A1(n_1035),
.A2(n_908),
.B1(n_861),
.B2(n_874),
.Y(n_1161)
);

OR2x6_ASAP7_75t_L g1162 ( 
.A(n_1025),
.B(n_739),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1039),
.A2(n_912),
.B(n_748),
.Y(n_1163)
);

INVx5_ASAP7_75t_L g1164 ( 
.A(n_919),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_938),
.B(n_777),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_926),
.A2(n_1005),
.B(n_1008),
.Y(n_1166)
);

INVxp67_ASAP7_75t_SL g1167 ( 
.A(n_1049),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1039),
.A2(n_912),
.B(n_748),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_992),
.B(n_996),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_992),
.B(n_996),
.Y(n_1170)
);

INVx5_ASAP7_75t_L g1171 ( 
.A(n_919),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_926),
.A2(n_1005),
.B(n_1008),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_938),
.B(n_296),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_926),
.A2(n_1005),
.B(n_1008),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1039),
.A2(n_912),
.B(n_748),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_931),
.Y(n_1176)
);

NOR2xp67_ASAP7_75t_L g1177 ( 
.A(n_993),
.B(n_886),
.Y(n_1177)
);

OR2x6_ASAP7_75t_L g1178 ( 
.A(n_1025),
.B(n_739),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_934),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1137),
.B(n_1139),
.Y(n_1180)
);

NOR2xp67_ASAP7_75t_L g1181 ( 
.A(n_1150),
.B(n_1147),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1068),
.A2(n_1066),
.B(n_1081),
.Y(n_1182)
);

AND2x2_ASAP7_75t_SL g1183 ( 
.A(n_1109),
.B(n_1156),
.Y(n_1183)
);

AOI222xp33_ASAP7_75t_L g1184 ( 
.A1(n_1092),
.A2(n_1173),
.B1(n_1160),
.B2(n_1135),
.C1(n_1177),
.C2(n_1108),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1141),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_1164),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1143),
.Y(n_1187)
);

NOR2xp67_ASAP7_75t_L g1188 ( 
.A(n_1064),
.B(n_1061),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1148),
.A2(n_1153),
.B(n_1152),
.Y(n_1189)
);

NAND2x1p5_ASAP7_75t_L g1190 ( 
.A(n_1164),
.B(n_1171),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1166),
.A2(n_1172),
.B(n_1174),
.Y(n_1191)
);

INVx3_ASAP7_75t_L g1192 ( 
.A(n_1145),
.Y(n_1192)
);

NOR2xp67_ASAP7_75t_L g1193 ( 
.A(n_1107),
.B(n_1128),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1165),
.B(n_1090),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_1072),
.Y(n_1195)
);

CKINVDCx20_ASAP7_75t_R g1196 ( 
.A(n_1096),
.Y(n_1196)
);

AO31x2_ASAP7_75t_L g1197 ( 
.A1(n_1093),
.A2(n_1055),
.A3(n_1092),
.B(n_1161),
.Y(n_1197)
);

NAND2x1p5_ASAP7_75t_L g1198 ( 
.A(n_1164),
.B(n_1171),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1109),
.B(n_1132),
.Y(n_1199)
);

NAND2xp33_ASAP7_75t_SL g1200 ( 
.A(n_1140),
.B(n_1142),
.Y(n_1200)
);

NAND2x1p5_ASAP7_75t_L g1201 ( 
.A(n_1171),
.B(n_1145),
.Y(n_1201)
);

CKINVDCx11_ASAP7_75t_R g1202 ( 
.A(n_1058),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1146),
.B(n_1157),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1103),
.A2(n_1134),
.B(n_1177),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1159),
.A2(n_1170),
.B(n_1169),
.C(n_1052),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1071),
.A2(n_1167),
.B1(n_1060),
.B2(n_1113),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_1144),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1179),
.Y(n_1208)
);

NAND2x1p5_ASAP7_75t_L g1209 ( 
.A(n_1074),
.B(n_1106),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1086),
.A2(n_1082),
.B1(n_1102),
.B2(n_1052),
.Y(n_1210)
);

NAND2x1p5_ASAP7_75t_L g1211 ( 
.A(n_1074),
.B(n_1095),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_SL g1212 ( 
.A(n_1067),
.B(n_1073),
.Y(n_1212)
);

OAI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1101),
.A2(n_1121),
.B(n_1071),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1102),
.A2(n_1062),
.B(n_1059),
.C(n_1063),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1084),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1149),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1110),
.B(n_1077),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_1105),
.B(n_1162),
.Y(n_1218)
);

O2A1O1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_1116),
.A2(n_1112),
.B(n_1079),
.C(n_1056),
.Y(n_1219)
);

AO31x2_ASAP7_75t_L g1220 ( 
.A1(n_1116),
.A2(n_1120),
.A3(n_1070),
.B(n_1065),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1085),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1097),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1098),
.A2(n_1122),
.B(n_1119),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1099),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1144),
.Y(n_1225)
);

INVx1_ASAP7_75t_SL g1226 ( 
.A(n_1054),
.Y(n_1226)
);

OA21x2_ASAP7_75t_L g1227 ( 
.A1(n_1062),
.A2(n_1114),
.B(n_1117),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1151),
.A2(n_1156),
.B(n_1115),
.Y(n_1228)
);

AOI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1118),
.A2(n_1075),
.B(n_1104),
.Y(n_1229)
);

BUFx2_ASAP7_75t_L g1230 ( 
.A(n_1094),
.Y(n_1230)
);

AND2x4_ASAP7_75t_L g1231 ( 
.A(n_1105),
.B(n_1178),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1057),
.B(n_1086),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1123),
.A2(n_1130),
.B(n_1127),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1076),
.B(n_1078),
.Y(n_1234)
);

OA21x2_ASAP7_75t_L g1235 ( 
.A1(n_1080),
.A2(n_1085),
.B(n_1158),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1129),
.A2(n_1128),
.B(n_1125),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1091),
.B(n_1136),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_L g1238 ( 
.A(n_1083),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1126),
.Y(n_1239)
);

AO21x2_ASAP7_75t_L g1240 ( 
.A1(n_1069),
.A2(n_1085),
.B(n_1053),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1124),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1162),
.A2(n_1178),
.B1(n_1133),
.B2(n_1136),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1053),
.A2(n_1158),
.B(n_1155),
.Y(n_1243)
);

NAND2x1_ASAP7_75t_L g1244 ( 
.A(n_1162),
.B(n_1178),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1054),
.B(n_1138),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1053),
.A2(n_1158),
.B(n_1155),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1154),
.A2(n_1155),
.B(n_1080),
.Y(n_1247)
);

BUFx2_ASAP7_75t_L g1248 ( 
.A(n_1176),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_SL g1249 ( 
.A1(n_1080),
.A2(n_1131),
.B1(n_1133),
.B2(n_1154),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1083),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1083),
.Y(n_1251)
);

BUFx4_ASAP7_75t_SL g1252 ( 
.A(n_1133),
.Y(n_1252)
);

NAND3xp33_ASAP7_75t_L g1253 ( 
.A(n_1089),
.B(n_1154),
.C(n_1100),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1089),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1131),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1089),
.A2(n_783),
.B1(n_1035),
.B2(n_950),
.Y(n_1256)
);

O2A1O1Ixp33_ASAP7_75t_SL g1257 ( 
.A1(n_1135),
.A2(n_995),
.B(n_783),
.C(n_1132),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1165),
.B(n_898),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_SL g1259 ( 
.A(n_1067),
.B(n_921),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_1090),
.B(n_1111),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1173),
.B(n_783),
.Y(n_1261)
);

INVx2_ASAP7_75t_SL g1262 ( 
.A(n_1144),
.Y(n_1262)
);

BUFx12f_ASAP7_75t_L g1263 ( 
.A(n_1096),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1109),
.A2(n_1139),
.B1(n_1140),
.B2(n_1137),
.Y(n_1264)
);

AO31x2_ASAP7_75t_L g1265 ( 
.A1(n_1093),
.A2(n_1135),
.A3(n_1055),
.B(n_995),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1163),
.A2(n_1175),
.B(n_1168),
.Y(n_1266)
);

OAI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1135),
.A2(n_586),
.B(n_592),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1068),
.A2(n_1066),
.B(n_1081),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1163),
.A2(n_1175),
.B(n_1168),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1051),
.Y(n_1270)
);

OA21x2_ASAP7_75t_L g1271 ( 
.A1(n_1160),
.A2(n_1087),
.B(n_1088),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1163),
.A2(n_1175),
.B(n_1168),
.Y(n_1272)
);

CKINVDCx6p67_ASAP7_75t_R g1273 ( 
.A(n_1058),
.Y(n_1273)
);

INVxp67_ASAP7_75t_L g1274 ( 
.A(n_1165),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1160),
.A2(n_783),
.B1(n_1035),
.B2(n_950),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1135),
.A2(n_586),
.B(n_592),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1137),
.B(n_1139),
.Y(n_1277)
);

OR2x2_ASAP7_75t_L g1278 ( 
.A(n_1054),
.B(n_1136),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1173),
.B(n_783),
.Y(n_1279)
);

OAI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1135),
.A2(n_586),
.B(n_592),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1147),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_1164),
.Y(n_1282)
);

OA21x2_ASAP7_75t_L g1283 ( 
.A1(n_1160),
.A2(n_1087),
.B(n_1088),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1163),
.A2(n_1175),
.B(n_1168),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1068),
.A2(n_1066),
.B(n_1081),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1137),
.B(n_1139),
.Y(n_1286)
);

BUFx4f_ASAP7_75t_L g1287 ( 
.A(n_1058),
.Y(n_1287)
);

O2A1O1Ixp5_ASAP7_75t_L g1288 ( 
.A1(n_1267),
.A2(n_1276),
.B(n_1280),
.C(n_1199),
.Y(n_1288)
);

OR2x2_ASAP7_75t_L g1289 ( 
.A(n_1278),
.B(n_1217),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_SL g1290 ( 
.A1(n_1205),
.A2(n_1203),
.B(n_1180),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1255),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1187),
.Y(n_1292)
);

OR2x2_ASAP7_75t_L g1293 ( 
.A(n_1258),
.B(n_1226),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_SL g1294 ( 
.A1(n_1205),
.A2(n_1286),
.B(n_1277),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1261),
.A2(n_1279),
.B1(n_1275),
.B2(n_1188),
.Y(n_1295)
);

O2A1O1Ixp5_ASAP7_75t_L g1296 ( 
.A1(n_1199),
.A2(n_1204),
.B(n_1213),
.C(n_1279),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1261),
.A2(n_1275),
.B1(n_1210),
.B2(n_1256),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1210),
.A2(n_1256),
.B1(n_1181),
.B2(n_1234),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1234),
.A2(n_1232),
.B1(n_1193),
.B2(n_1274),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1264),
.B(n_1184),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1274),
.A2(n_1237),
.B1(n_1209),
.B2(n_1242),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_SL g1302 ( 
.A1(n_1214),
.A2(n_1190),
.B(n_1198),
.Y(n_1302)
);

CKINVDCx14_ASAP7_75t_R g1303 ( 
.A(n_1196),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_SL g1304 ( 
.A1(n_1214),
.A2(n_1190),
.B(n_1198),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1241),
.B(n_1206),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1209),
.A2(n_1253),
.B1(n_1230),
.B2(n_1229),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1194),
.B(n_1218),
.Y(n_1307)
);

OA21x2_ASAP7_75t_L g1308 ( 
.A1(n_1223),
.A2(n_1243),
.B(n_1246),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1200),
.B(n_1281),
.Y(n_1309)
);

AND2x4_ASAP7_75t_L g1310 ( 
.A(n_1218),
.B(n_1231),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1231),
.B(n_1248),
.Y(n_1311)
);

AOI211xp5_ASAP7_75t_L g1312 ( 
.A1(n_1257),
.A2(n_1219),
.B(n_1245),
.C(n_1228),
.Y(n_1312)
);

OA21x2_ASAP7_75t_L g1313 ( 
.A1(n_1266),
.A2(n_1269),
.B(n_1284),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1185),
.B(n_1216),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1211),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1249),
.A2(n_1287),
.B1(n_1244),
.B2(n_1183),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1287),
.A2(n_1183),
.B1(n_1270),
.B2(n_1208),
.Y(n_1317)
);

OR2x2_ASAP7_75t_L g1318 ( 
.A(n_1197),
.B(n_1265),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1215),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_SL g1320 ( 
.A1(n_1186),
.A2(n_1282),
.B(n_1207),
.Y(n_1320)
);

O2A1O1Ixp5_ASAP7_75t_L g1321 ( 
.A1(n_1272),
.A2(n_1221),
.B(n_1239),
.C(n_1222),
.Y(n_1321)
);

BUFx10_ASAP7_75t_L g1322 ( 
.A(n_1262),
.Y(n_1322)
);

A2O1A1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1247),
.A2(n_1224),
.B(n_1265),
.C(n_1233),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1195),
.A2(n_1207),
.B1(n_1225),
.B2(n_1201),
.Y(n_1324)
);

OR2x2_ASAP7_75t_L g1325 ( 
.A(n_1197),
.B(n_1265),
.Y(n_1325)
);

OA21x2_ASAP7_75t_L g1326 ( 
.A1(n_1189),
.A2(n_1191),
.B(n_1182),
.Y(n_1326)
);

INVx1_ASAP7_75t_SL g1327 ( 
.A(n_1195),
.Y(n_1327)
);

O2A1O1Ixp5_ASAP7_75t_L g1328 ( 
.A1(n_1192),
.A2(n_1250),
.B(n_1251),
.C(n_1265),
.Y(n_1328)
);

INVx1_ASAP7_75t_SL g1329 ( 
.A(n_1260),
.Y(n_1329)
);

O2A1O1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1225),
.A2(n_1212),
.B(n_1259),
.C(n_1201),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1273),
.A2(n_1186),
.B1(n_1282),
.B2(n_1254),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1236),
.B(n_1238),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_SL g1333 ( 
.A1(n_1186),
.A2(n_1282),
.B(n_1227),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_SL g1334 ( 
.A1(n_1186),
.A2(n_1282),
.B(n_1227),
.Y(n_1334)
);

AND2x6_ASAP7_75t_L g1335 ( 
.A(n_1238),
.B(n_1252),
.Y(n_1335)
);

OR2x2_ASAP7_75t_L g1336 ( 
.A(n_1197),
.B(n_1220),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1197),
.B(n_1238),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1235),
.B(n_1240),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1235),
.B(n_1240),
.Y(n_1339)
);

NOR2xp67_ASAP7_75t_L g1340 ( 
.A(n_1263),
.B(n_1202),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1196),
.A2(n_1283),
.B1(n_1271),
.B2(n_1202),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1268),
.B(n_1285),
.Y(n_1342)
);

BUFx8_ASAP7_75t_SL g1343 ( 
.A(n_1196),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1278),
.B(n_1217),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1258),
.B(n_1194),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1217),
.B(n_1180),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1261),
.A2(n_1109),
.B1(n_1279),
.B2(n_1275),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1258),
.B(n_1194),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_1194),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1261),
.B(n_1279),
.Y(n_1350)
);

BUFx2_ASAP7_75t_R g1351 ( 
.A(n_1207),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_1230),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1217),
.B(n_1180),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1258),
.B(n_1194),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1261),
.A2(n_1109),
.B1(n_1279),
.B2(n_1275),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1217),
.B(n_1180),
.Y(n_1356)
);

NAND2x1p5_ASAP7_75t_L g1357 ( 
.A(n_1233),
.B(n_1228),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1336),
.B(n_1318),
.Y(n_1358)
);

CKINVDCx20_ASAP7_75t_R g1359 ( 
.A(n_1343),
.Y(n_1359)
);

INVx2_ASAP7_75t_SL g1360 ( 
.A(n_1332),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1337),
.B(n_1325),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_1332),
.B(n_1323),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1309),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1308),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1301),
.Y(n_1365)
);

BUFx2_ASAP7_75t_L g1366 ( 
.A(n_1315),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1305),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1291),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_1303),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1342),
.B(n_1292),
.Y(n_1370)
);

INVx4_ASAP7_75t_L g1371 ( 
.A(n_1335),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1357),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1341),
.B(n_1338),
.Y(n_1373)
);

OR2x6_ASAP7_75t_L g1374 ( 
.A(n_1333),
.B(n_1334),
.Y(n_1374)
);

AOI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1350),
.A2(n_1347),
.B1(n_1355),
.B2(n_1297),
.Y(n_1375)
);

INVx1_ASAP7_75t_SL g1376 ( 
.A(n_1352),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1339),
.B(n_1289),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1319),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1350),
.A2(n_1300),
.B1(n_1295),
.B2(n_1298),
.Y(n_1379)
);

OA21x2_ASAP7_75t_L g1380 ( 
.A1(n_1321),
.A2(n_1288),
.B(n_1328),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1306),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1290),
.B(n_1294),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1317),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1344),
.B(n_1293),
.Y(n_1384)
);

OR2x6_ASAP7_75t_L g1385 ( 
.A(n_1302),
.B(n_1304),
.Y(n_1385)
);

AO21x2_ASAP7_75t_L g1386 ( 
.A1(n_1316),
.A2(n_1299),
.B(n_1314),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1346),
.B(n_1356),
.Y(n_1387)
);

BUFx2_ASAP7_75t_L g1388 ( 
.A(n_1311),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1345),
.B(n_1354),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1328),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1296),
.Y(n_1391)
);

OR2x6_ASAP7_75t_L g1392 ( 
.A(n_1330),
.B(n_1320),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1367),
.B(n_1353),
.Y(n_1393)
);

AOI221xp5_ASAP7_75t_L g1394 ( 
.A1(n_1375),
.A2(n_1379),
.B1(n_1296),
.B2(n_1391),
.C(n_1382),
.Y(n_1394)
);

INVx4_ASAP7_75t_L g1395 ( 
.A(n_1385),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1362),
.B(n_1310),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1377),
.B(n_1313),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1370),
.B(n_1361),
.Y(n_1398)
);

INVxp67_ASAP7_75t_SL g1399 ( 
.A(n_1368),
.Y(n_1399)
);

AND2x4_ASAP7_75t_L g1400 ( 
.A(n_1362),
.B(n_1310),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1368),
.Y(n_1401)
);

BUFx3_ASAP7_75t_L g1402 ( 
.A(n_1366),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1370),
.B(n_1326),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1391),
.B(n_1312),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1378),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1370),
.B(n_1348),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1370),
.B(n_1349),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1361),
.B(n_1307),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1358),
.B(n_1324),
.Y(n_1409)
);

INVx4_ASAP7_75t_L g1410 ( 
.A(n_1385),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1358),
.B(n_1327),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1394),
.A2(n_1375),
.B1(n_1382),
.B2(n_1392),
.Y(n_1412)
);

AO21x2_ASAP7_75t_L g1413 ( 
.A1(n_1404),
.A2(n_1364),
.B(n_1390),
.Y(n_1413)
);

OAI21xp33_ASAP7_75t_L g1414 ( 
.A1(n_1394),
.A2(n_1381),
.B(n_1365),
.Y(n_1414)
);

HB1xp67_ASAP7_75t_L g1415 ( 
.A(n_1401),
.Y(n_1415)
);

INVx2_ASAP7_75t_SL g1416 ( 
.A(n_1402),
.Y(n_1416)
);

AOI221xp5_ASAP7_75t_L g1417 ( 
.A1(n_1404),
.A2(n_1381),
.B1(n_1363),
.B2(n_1387),
.C(n_1376),
.Y(n_1417)
);

AO21x1_ASAP7_75t_SL g1418 ( 
.A1(n_1409),
.A2(n_1373),
.B(n_1390),
.Y(n_1418)
);

INVxp67_ASAP7_75t_L g1419 ( 
.A(n_1411),
.Y(n_1419)
);

AOI222xp33_ASAP7_75t_L g1420 ( 
.A1(n_1393),
.A2(n_1383),
.B1(n_1387),
.B2(n_1340),
.C1(n_1369),
.C2(n_1376),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1398),
.B(n_1360),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1401),
.Y(n_1422)
);

NAND3xp33_ASAP7_75t_L g1423 ( 
.A(n_1393),
.B(n_1385),
.C(n_1392),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1395),
.A2(n_1383),
.B1(n_1385),
.B2(n_1386),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1399),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1398),
.B(n_1373),
.Y(n_1426)
);

INVx5_ASAP7_75t_L g1427 ( 
.A(n_1395),
.Y(n_1427)
);

OAI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1395),
.A2(n_1385),
.B1(n_1392),
.B2(n_1374),
.Y(n_1428)
);

OAI31xp33_ASAP7_75t_L g1429 ( 
.A1(n_1409),
.A2(n_1331),
.A3(n_1329),
.B(n_1384),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1395),
.A2(n_1386),
.B1(n_1392),
.B2(n_1374),
.Y(n_1430)
);

INVx2_ASAP7_75t_SL g1431 ( 
.A(n_1402),
.Y(n_1431)
);

INVx4_ASAP7_75t_L g1432 ( 
.A(n_1395),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1399),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1411),
.A2(n_1371),
.B1(n_1374),
.B2(n_1351),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1410),
.A2(n_1386),
.B1(n_1374),
.B2(n_1388),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1405),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1403),
.B(n_1372),
.Y(n_1437)
);

OAI221xp5_ASAP7_75t_L g1438 ( 
.A1(n_1410),
.A2(n_1409),
.B1(n_1384),
.B2(n_1411),
.C(n_1397),
.Y(n_1438)
);

INVx1_ASAP7_75t_SL g1439 ( 
.A(n_1415),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1422),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_SL g1441 ( 
.A(n_1417),
.B(n_1396),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1413),
.Y(n_1442)
);

INVxp67_ASAP7_75t_L g1443 ( 
.A(n_1418),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1413),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1418),
.B(n_1406),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1436),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1436),
.Y(n_1447)
);

OR2x6_ASAP7_75t_L g1448 ( 
.A(n_1423),
.B(n_1410),
.Y(n_1448)
);

INVxp33_ASAP7_75t_L g1449 ( 
.A(n_1434),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_1416),
.Y(n_1450)
);

NAND2x1p5_ASAP7_75t_SL g1451 ( 
.A(n_1416),
.B(n_1431),
.Y(n_1451)
);

INVx4_ASAP7_75t_SL g1452 ( 
.A(n_1431),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1419),
.B(n_1425),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1426),
.B(n_1403),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1426),
.B(n_1403),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_SL g1456 ( 
.A(n_1420),
.B(n_1396),
.Y(n_1456)
);

INVx4_ASAP7_75t_SL g1457 ( 
.A(n_1425),
.Y(n_1457)
);

OR2x6_ASAP7_75t_L g1458 ( 
.A(n_1423),
.B(n_1410),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1420),
.B(n_1396),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1414),
.B(n_1359),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1445),
.B(n_1437),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1452),
.B(n_1427),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1441),
.B(n_1414),
.Y(n_1463)
);

INVxp33_ASAP7_75t_L g1464 ( 
.A(n_1460),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1446),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1446),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1453),
.B(n_1433),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1445),
.B(n_1437),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1443),
.B(n_1437),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1451),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1443),
.B(n_1421),
.Y(n_1471)
);

OR2x6_ASAP7_75t_L g1472 ( 
.A(n_1448),
.B(n_1432),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1449),
.A2(n_1412),
.B1(n_1430),
.B2(n_1428),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_SL g1474 ( 
.A(n_1448),
.B(n_1429),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1439),
.B(n_1406),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1447),
.Y(n_1476)
);

NOR4xp25_ASAP7_75t_L g1477 ( 
.A(n_1456),
.B(n_1438),
.C(n_1424),
.D(n_1435),
.Y(n_1477)
);

NAND2x1p5_ASAP7_75t_L g1478 ( 
.A(n_1440),
.B(n_1427),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1439),
.B(n_1406),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1447),
.Y(n_1480)
);

NOR2x1p5_ASAP7_75t_L g1481 ( 
.A(n_1450),
.B(n_1432),
.Y(n_1481)
);

NAND4xp25_ASAP7_75t_L g1482 ( 
.A(n_1459),
.B(n_1429),
.C(n_1397),
.D(n_1407),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_L g1483 ( 
.A(n_1450),
.B(n_1322),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1440),
.B(n_1408),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1457),
.B(n_1450),
.Y(n_1485)
);

AND2x4_ASAP7_75t_SL g1486 ( 
.A(n_1448),
.B(n_1458),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1457),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1457),
.B(n_1448),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_SL g1489 ( 
.A1(n_1448),
.A2(n_1371),
.B1(n_1396),
.B2(n_1400),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1465),
.Y(n_1490)
);

OAI22xp33_ASAP7_75t_SL g1491 ( 
.A1(n_1474),
.A2(n_1458),
.B1(n_1448),
.B2(n_1444),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1488),
.B(n_1461),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1488),
.B(n_1454),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1463),
.B(n_1455),
.Y(n_1494)
);

OAI21xp33_ASAP7_75t_L g1495 ( 
.A1(n_1477),
.A2(n_1458),
.B(n_1444),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1465),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1466),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1466),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1476),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1483),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1488),
.B(n_1455),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1467),
.B(n_1451),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1461),
.B(n_1455),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1464),
.B(n_1322),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1468),
.B(n_1457),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1476),
.Y(n_1506)
);

NOR2xp67_ASAP7_75t_SL g1507 ( 
.A(n_1470),
.B(n_1371),
.Y(n_1507)
);

INVx1_ASAP7_75t_SL g1508 ( 
.A(n_1469),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1480),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1484),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1473),
.B(n_1408),
.Y(n_1511)
);

NAND2x1p5_ASAP7_75t_L g1512 ( 
.A(n_1470),
.B(n_1380),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1471),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1475),
.Y(n_1514)
);

OAI21xp33_ASAP7_75t_SL g1515 ( 
.A1(n_1481),
.A2(n_1458),
.B(n_1442),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1482),
.B(n_1389),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1468),
.B(n_1457),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1479),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1496),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1512),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1496),
.Y(n_1521)
);

INVx3_ASAP7_75t_L g1522 ( 
.A(n_1512),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1505),
.B(n_1485),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_1500),
.B(n_1487),
.Y(n_1524)
);

INVxp33_ASAP7_75t_L g1525 ( 
.A(n_1507),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1497),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1512),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1505),
.B(n_1485),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1517),
.B(n_1485),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1513),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1517),
.B(n_1478),
.Y(n_1531)
);

INVxp67_ASAP7_75t_SL g1532 ( 
.A(n_1502),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_1500),
.Y(n_1533)
);

NOR2xp67_ASAP7_75t_L g1534 ( 
.A(n_1515),
.B(n_1462),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1503),
.B(n_1478),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1513),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1495),
.A2(n_1458),
.B1(n_1486),
.B2(n_1472),
.Y(n_1537)
);

NOR2x1_ASAP7_75t_L g1538 ( 
.A(n_1502),
.B(n_1481),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1491),
.A2(n_1458),
.B1(n_1486),
.B2(n_1472),
.Y(n_1539)
);

CKINVDCx16_ASAP7_75t_R g1540 ( 
.A(n_1504),
.Y(n_1540)
);

INVx1_ASAP7_75t_SL g1541 ( 
.A(n_1508),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1497),
.Y(n_1542)
);

INVx4_ASAP7_75t_L g1543 ( 
.A(n_1492),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1541),
.B(n_1532),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1523),
.B(n_1492),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1523),
.B(n_1493),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1530),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1543),
.Y(n_1548)
);

AOI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1533),
.A2(n_1489),
.B1(n_1507),
.B2(n_1510),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1530),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1530),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1537),
.A2(n_1539),
.B1(n_1532),
.B2(n_1541),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1530),
.Y(n_1553)
);

AOI21xp5_ASAP7_75t_L g1554 ( 
.A1(n_1537),
.A2(n_1511),
.B(n_1494),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1524),
.B(n_1516),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1543),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1543),
.B(n_1493),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1524),
.B(n_1503),
.Y(n_1558)
);

OAI21xp33_ASAP7_75t_L g1559 ( 
.A1(n_1539),
.A2(n_1514),
.B(n_1518),
.Y(n_1559)
);

AOI221xp5_ASAP7_75t_L g1560 ( 
.A1(n_1525),
.A2(n_1518),
.B1(n_1498),
.B2(n_1499),
.C(n_1506),
.Y(n_1560)
);

INVxp67_ASAP7_75t_L g1561 ( 
.A(n_1523),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1536),
.Y(n_1562)
);

AOI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1528),
.A2(n_1472),
.B1(n_1501),
.B2(n_1469),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1544),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1561),
.B(n_1543),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1545),
.B(n_1543),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1546),
.B(n_1528),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1544),
.Y(n_1568)
);

INVx2_ASAP7_75t_SL g1569 ( 
.A(n_1557),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1558),
.B(n_1540),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1557),
.B(n_1540),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1556),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1560),
.B(n_1536),
.Y(n_1573)
);

AOI221xp5_ASAP7_75t_L g1574 ( 
.A1(n_1573),
.A2(n_1552),
.B1(n_1554),
.B2(n_1559),
.C(n_1555),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1567),
.B(n_1548),
.Y(n_1575)
);

AOI21xp33_ASAP7_75t_SL g1576 ( 
.A1(n_1571),
.A2(n_1552),
.B(n_1525),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1570),
.B(n_1528),
.Y(n_1577)
);

O2A1O1Ixp33_ASAP7_75t_L g1578 ( 
.A1(n_1573),
.A2(n_1538),
.B(n_1562),
.C(n_1553),
.Y(n_1578)
);

OA22x2_ASAP7_75t_L g1579 ( 
.A1(n_1569),
.A2(n_1549),
.B1(n_1563),
.B2(n_1529),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1564),
.A2(n_1568),
.B1(n_1529),
.B2(n_1534),
.Y(n_1580)
);

OAI221xp5_ASAP7_75t_L g1581 ( 
.A1(n_1566),
.A2(n_1538),
.B1(n_1565),
.B2(n_1534),
.C(n_1572),
.Y(n_1581)
);

AOI221xp5_ASAP7_75t_L g1582 ( 
.A1(n_1573),
.A2(n_1531),
.B1(n_1519),
.B2(n_1526),
.C(n_1542),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1575),
.Y(n_1583)
);

NAND5xp2_ASAP7_75t_L g1584 ( 
.A(n_1574),
.B(n_1551),
.C(n_1550),
.D(n_1547),
.E(n_1529),
.Y(n_1584)
);

OAI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1580),
.A2(n_1531),
.B1(n_1472),
.B2(n_1478),
.Y(n_1585)
);

NAND3x1_ASAP7_75t_L g1586 ( 
.A(n_1577),
.B(n_1531),
.C(n_1521),
.Y(n_1586)
);

OAI22xp33_ASAP7_75t_SL g1587 ( 
.A1(n_1581),
.A2(n_1536),
.B1(n_1522),
.B2(n_1520),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1584),
.B(n_1576),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1586),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1583),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1587),
.Y(n_1591)
);

AOI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1585),
.A2(n_1579),
.B1(n_1582),
.B2(n_1536),
.Y(n_1592)
);

INVx1_ASAP7_75t_SL g1593 ( 
.A(n_1586),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1588),
.A2(n_1578),
.B(n_1521),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1589),
.Y(n_1595)
);

NOR2x1_ASAP7_75t_L g1596 ( 
.A(n_1593),
.B(n_1519),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1591),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1592),
.B(n_1535),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1596),
.Y(n_1599)
);

NOR2x1_ASAP7_75t_L g1600 ( 
.A(n_1594),
.B(n_1590),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1598),
.B(n_1526),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1599),
.Y(n_1602)
);

INVx1_ASAP7_75t_SL g1603 ( 
.A(n_1602),
.Y(n_1603)
);

XOR2xp5_ASAP7_75t_L g1604 ( 
.A(n_1603),
.B(n_1597),
.Y(n_1604)
);

INVx3_ASAP7_75t_L g1605 ( 
.A(n_1604),
.Y(n_1605)
);

AOI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1605),
.A2(n_1595),
.B1(n_1600),
.B2(n_1601),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1606),
.A2(n_1605),
.B1(n_1542),
.B2(n_1527),
.Y(n_1607)
);

OR3x2_ASAP7_75t_L g1608 ( 
.A(n_1607),
.B(n_1509),
.C(n_1490),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1608),
.B(n_1535),
.Y(n_1609)
);

OAI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1608),
.A2(n_1527),
.B(n_1522),
.Y(n_1610)
);

OAI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1609),
.A2(n_1610),
.B(n_1527),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1609),
.A2(n_1527),
.B1(n_1520),
.B2(n_1522),
.Y(n_1612)
);

AOI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1612),
.A2(n_1522),
.B1(n_1520),
.B2(n_1535),
.Y(n_1613)
);

AOI211xp5_ASAP7_75t_L g1614 ( 
.A1(n_1613),
.A2(n_1611),
.B(n_1522),
.C(n_1520),
.Y(n_1614)
);


endmodule