module fake_jpeg_21268_n_135 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx13_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx5p33_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx4f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_29),
.Y(n_41)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_13),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_14),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_25),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_33),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_24),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_32),
.B1(n_29),
.B2(n_16),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_27),
.A2(n_22),
.B1(n_16),
.B2(n_14),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_22),
.B1(n_26),
.B2(n_20),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_29),
.Y(n_55)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_25),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_44),
.B(n_33),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_32),
.B(n_27),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_58),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_47),
.B(n_49),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_34),
.C(n_28),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_42),
.C(n_39),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

NOR3xp33_ASAP7_75t_SL g52 ( 
.A(n_36),
.B(n_30),
.C(n_34),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_52),
.B(n_60),
.Y(n_79)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_59),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_34),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_33),
.B(n_23),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_33),
.B1(n_30),
.B2(n_31),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_33),
.B1(n_43),
.B2(n_37),
.Y(n_64)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

AND2x6_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_31),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_20),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_61),
.B(n_21),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_12),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_64),
.A2(n_43),
.B1(n_37),
.B2(n_59),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_76),
.C(n_50),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_50),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_71),
.B(n_78),
.Y(n_89)
);

XNOR2x1_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_75),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_77),
.Y(n_88)
);

NOR2xp67_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_19),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_39),
.C(n_24),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_51),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_26),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_57),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_80),
.A2(n_84),
.B(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_83),
.Y(n_94)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_79),
.A2(n_52),
.B(n_57),
.Y(n_84)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_57),
.B(n_56),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_90),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_56),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_92),
.Y(n_100)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_63),
.B1(n_65),
.B2(n_70),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_69),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_95),
.B(n_98),
.Y(n_112)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_97),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_69),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_SL g101 ( 
.A1(n_87),
.A2(n_85),
.B(n_80),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_101),
.A2(n_80),
.B(n_84),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_68),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_103),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_103),
.A2(n_15),
.B1(n_19),
.B2(n_21),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_106),
.Y(n_115)
);

AO221x1_ASAP7_75t_L g106 ( 
.A1(n_101),
.A2(n_94),
.B1(n_53),
.B2(n_87),
.C(n_39),
.Y(n_106)
);

OAI322xp33_ASAP7_75t_L g107 ( 
.A1(n_99),
.A2(n_72),
.A3(n_91),
.B1(n_76),
.B2(n_77),
.C1(n_19),
.C2(n_21),
.Y(n_107)
);

NOR3xp33_ASAP7_75t_SL g117 ( 
.A(n_107),
.B(n_19),
.C(n_21),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_15),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_104),
.A2(n_53),
.B(n_2),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_111),
.A2(n_112),
.B1(n_104),
.B2(n_109),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_113),
.B(n_24),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_100),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_116),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_117),
.B(n_118),
.Y(n_120)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_114),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_123),
.Y(n_126)
);

OAI21x1_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_111),
.B(n_110),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_113),
.B1(n_108),
.B2(n_105),
.Y(n_125)
);

INVxp33_ASAP7_75t_L g131 ( 
.A(n_125),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_108),
.C(n_117),
.Y(n_127)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_127),
.A2(n_128),
.A3(n_120),
.B1(n_12),
.B2(n_15),
.C1(n_10),
.C2(n_7),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_124),
.A2(n_15),
.B1(n_8),
.B2(n_6),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_129),
.A2(n_127),
.B1(n_5),
.B2(n_3),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_L g130 ( 
.A1(n_126),
.A2(n_12),
.A3(n_10),
.B1(n_18),
.B2(n_5),
.C1(n_0),
.C2(n_4),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_130),
.Y(n_132)
);

OAI221xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_18),
.B1(n_24),
.B2(n_131),
.C(n_132),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_18),
.Y(n_135)
);


endmodule