module fake_jpeg_12560_n_437 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_437);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_437;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_3),
.B(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g112 ( 
.A(n_48),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_6),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_50),
.B(n_53),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_56),
.Y(n_127)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_57),
.Y(n_140)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_27),
.B(n_6),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_59),
.B(n_63),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_61),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_62),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_27),
.B(n_6),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_64),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_66),
.Y(n_143)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_27),
.B(n_7),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_68),
.B(n_70),
.Y(n_121)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_19),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_19),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_72),
.B(n_75),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_74),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_43),
.Y(n_75)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

BUFx10_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_77),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_23),
.Y(n_80)
);

NAND2xp33_ASAP7_75t_SL g139 ( 
.A(n_80),
.B(n_83),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_43),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_82),
.B(n_84),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_20),
.B(n_28),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_20),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_86),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_28),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_16),
.B(n_7),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_88),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_30),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_91),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_92),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_16),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_53),
.A2(n_38),
.B1(n_16),
.B2(n_42),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_95),
.A2(n_113),
.B1(n_114),
.B2(n_118),
.Y(n_165)
);

AOI221xp5_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_30),
.B1(n_45),
.B2(n_35),
.C(n_33),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_98),
.B(n_101),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_66),
.A2(n_38),
.B1(n_40),
.B2(n_39),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_99),
.A2(n_106),
.B1(n_111),
.B2(n_117),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_77),
.A2(n_38),
.B1(n_40),
.B2(n_39),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_70),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_73),
.A2(n_42),
.B1(n_32),
.B2(n_41),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_73),
.A2(n_32),
.B1(n_41),
.B2(n_36),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_81),
.A2(n_32),
.B1(n_41),
.B2(n_36),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_115),
.A2(n_76),
.B1(n_62),
.B2(n_56),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_72),
.A2(n_46),
.B1(n_31),
.B2(n_33),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_80),
.A2(n_41),
.B1(n_36),
.B2(n_32),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_80),
.A2(n_25),
.B(n_36),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_129),
.A2(n_136),
.B(n_48),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_74),
.A2(n_41),
.B1(n_36),
.B2(n_32),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_131),
.A2(n_132),
.B1(n_142),
.B2(n_48),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_54),
.A2(n_35),
.B1(n_31),
.B2(n_25),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_75),
.B(n_0),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_0),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_67),
.B(n_7),
.C(n_12),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_0),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_69),
.A2(n_7),
.B1(n_12),
.B2(n_2),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_57),
.A2(n_58),
.B1(n_64),
.B2(n_89),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_109),
.A2(n_92),
.B(n_82),
.C(n_86),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_146),
.B(n_174),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_147),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_148),
.B(n_168),
.Y(n_200)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_149),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_150),
.B(n_172),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_151),
.Y(n_201)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_152),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_71),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_L g202 ( 
.A1(n_153),
.A2(n_158),
.B(n_163),
.Y(n_202)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_107),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_161),
.Y(n_198)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_55),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_107),
.Y(n_159)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

BUFx24_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

INVx3_ASAP7_75t_SL g230 ( 
.A(n_160),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_128),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_162),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_52),
.Y(n_163)
);

OA22x2_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_139),
.B1(n_124),
.B2(n_108),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_164),
.A2(n_169),
.B1(n_186),
.B2(n_187),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_110),
.Y(n_166)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_166),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_56),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_104),
.C(n_115),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_88),
.Y(n_168)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_L g171 ( 
.A1(n_108),
.A2(n_90),
.B1(n_83),
.B2(n_61),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_171),
.A2(n_178),
.B1(n_112),
.B2(n_140),
.Y(n_216)
);

OR2x4_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_48),
.Y(n_173)
);

NAND2xp67_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_176),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_121),
.B(n_85),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_96),
.Y(n_175)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_175),
.Y(n_214)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_119),
.B(n_135),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_181),
.Y(n_215)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_136),
.A2(n_56),
.B(n_78),
.C(n_47),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_102),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_182),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_126),
.B(n_79),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_184),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_102),
.B(n_91),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_103),
.B(n_9),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_192),
.Y(n_226)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_130),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g187 ( 
.A(n_127),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_145),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_220)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_100),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_144),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_103),
.B(n_9),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_146),
.A2(n_143),
.B1(n_130),
.B2(n_100),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_197),
.A2(n_206),
.B1(n_211),
.B2(n_213),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_199),
.B(n_229),
.C(n_180),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_164),
.A2(n_143),
.B1(n_123),
.B2(n_126),
.Y(n_206)
);

NAND2xp67_ASAP7_75t_L g209 ( 
.A(n_164),
.B(n_173),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_209),
.B(n_1),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_165),
.A2(n_94),
.B1(n_137),
.B2(n_134),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_164),
.A2(n_65),
.B1(n_51),
.B2(n_60),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_216),
.A2(n_231),
.B1(n_186),
.B2(n_170),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_154),
.A2(n_123),
.B1(n_116),
.B2(n_137),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_219),
.A2(n_224),
.B1(n_232),
.B2(n_120),
.Y(n_242)
);

AOI32xp33_ASAP7_75t_L g221 ( 
.A1(n_176),
.A2(n_120),
.A3(n_140),
.B1(n_97),
.B2(n_127),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_221),
.A2(n_160),
.B(n_190),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_171),
.A2(n_153),
.B1(n_163),
.B2(n_167),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_150),
.B(n_104),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_150),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_153),
.B(n_116),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_178),
.A2(n_94),
.B1(n_134),
.B2(n_60),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_163),
.A2(n_97),
.B1(n_112),
.B2(n_120),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_233),
.Y(n_268)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_204),
.Y(n_234)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_234),
.Y(n_276)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_214),
.Y(n_235)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_235),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_237),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_167),
.Y(n_237)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_238),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_198),
.B(n_158),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_239),
.B(n_242),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_207),
.A2(n_181),
.B(n_158),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_241),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_243),
.A2(n_232),
.B1(n_202),
.B2(n_199),
.Y(n_284)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_214),
.Y(n_244)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_244),
.Y(n_294)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_195),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_245),
.Y(n_279)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_195),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_246),
.Y(n_290)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_247),
.B(n_251),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_212),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_248),
.B(n_254),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_215),
.A2(n_160),
.B(n_147),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_249),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_228),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_256),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_208),
.B(n_149),
.Y(n_252)
);

NOR2x1_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_253),
.Y(n_272)
);

OAI21x1_ASAP7_75t_L g253 ( 
.A1(n_208),
.A2(n_191),
.B(n_189),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_188),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_266),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_218),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_224),
.A2(n_155),
.B1(n_177),
.B2(n_166),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_257),
.A2(n_263),
.B1(n_264),
.B2(n_230),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_200),
.B(n_151),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_258),
.B(n_259),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_205),
.B(n_187),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_222),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_262),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_215),
.A2(n_187),
.B(n_2),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_227),
.C(n_193),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_205),
.B(n_8),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_213),
.A2(n_8),
.B1(n_3),
.B2(n_4),
.Y(n_263)
);

OR2x6_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_1),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_264),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_218),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_196),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_209),
.B(n_1),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_193),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_270),
.A2(n_201),
.B1(n_217),
.B2(n_203),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_281),
.B(n_256),
.Y(n_300)
);

XOR2x1_ASAP7_75t_L g312 ( 
.A(n_283),
.B(n_233),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_284),
.A2(n_264),
.B1(n_257),
.B2(n_263),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_286),
.A2(n_264),
.B(n_234),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_243),
.A2(n_225),
.B1(n_210),
.B2(n_216),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_288),
.A2(n_298),
.B1(n_299),
.B2(n_264),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_237),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_292),
.C(n_293),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_236),
.B(n_210),
.C(n_225),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_254),
.B(n_210),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_240),
.A2(n_220),
.B1(n_194),
.B2(n_230),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_296),
.A2(n_297),
.B1(n_248),
.B2(n_238),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_240),
.A2(n_194),
.B1(n_230),
.B2(n_223),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_266),
.A2(n_252),
.B1(n_251),
.B2(n_241),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_242),
.A2(n_264),
.B1(n_239),
.B2(n_253),
.Y(n_299)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_300),
.Y(n_337)
);

MAJx2_ASAP7_75t_L g301 ( 
.A(n_271),
.B(n_267),
.C(n_258),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_301),
.B(n_286),
.C(n_271),
.Y(n_331)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_274),
.Y(n_302)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_302),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_303),
.A2(n_307),
.B1(n_318),
.B2(n_323),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_275),
.A2(n_250),
.B1(n_248),
.B2(n_265),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_304),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_277),
.B(n_262),
.Y(n_305)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_305),
.Y(n_335)
);

NAND3xp33_ASAP7_75t_L g306 ( 
.A(n_269),
.B(n_261),
.C(n_259),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_306),
.B(n_321),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_270),
.A2(n_264),
.B1(n_249),
.B2(n_267),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_308),
.A2(n_309),
.B1(n_311),
.B2(n_317),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_310),
.B(n_276),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_287),
.A2(n_298),
.B1(n_299),
.B2(n_275),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_312),
.B(n_283),
.Y(n_328)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_277),
.Y(n_314)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_314),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_272),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_315),
.B(n_320),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_295),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_319),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_287),
.Y(n_317)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_317),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_297),
.A2(n_244),
.B1(n_235),
.B2(n_248),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_280),
.B(n_260),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_295),
.B(n_247),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_272),
.B(n_246),
.Y(n_321)
);

OAI22x1_ASAP7_75t_L g322 ( 
.A1(n_273),
.A2(n_217),
.B1(n_245),
.B2(n_238),
.Y(n_322)
);

A2O1A1Ixp33_ASAP7_75t_SL g348 ( 
.A1(n_322),
.A2(n_291),
.B(n_294),
.C(n_285),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_269),
.B(n_196),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_324),
.B(n_326),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_282),
.A2(n_223),
.B(n_201),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_325),
.B(n_327),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_268),
.B(n_203),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_279),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_328),
.B(n_342),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_331),
.B(n_336),
.C(n_345),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_313),
.B(n_289),
.C(n_293),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_338),
.A2(n_346),
.B1(n_303),
.B2(n_321),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_307),
.A2(n_288),
.B1(n_284),
.B2(n_278),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_340),
.A2(n_311),
.B1(n_330),
.B2(n_308),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_320),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_341),
.B(n_302),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_313),
.B(n_312),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_327),
.B(n_290),
.Y(n_343)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_343),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_312),
.B(n_292),
.C(n_278),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_309),
.A2(n_296),
.B1(n_268),
.B2(n_276),
.Y(n_346)
);

OA22x2_ASAP7_75t_L g370 ( 
.A1(n_348),
.A2(n_318),
.B1(n_322),
.B2(n_291),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_301),
.B(n_294),
.C(n_285),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_349),
.B(n_325),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_351),
.B(n_324),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_353),
.B(n_362),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_356),
.A2(n_330),
.B1(n_340),
.B2(n_333),
.Y(n_375)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_357),
.Y(n_377)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_337),
.Y(n_358)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_358),
.Y(n_380)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_339),
.Y(n_359)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_359),
.Y(n_387)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_343),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_361),
.B(n_363),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_336),
.B(n_310),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_329),
.Y(n_364)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_364),
.B(n_365),
.Y(n_378)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_329),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_338),
.B(n_334),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_366),
.A2(n_368),
.B(n_369),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_331),
.B(n_301),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_367),
.B(n_371),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_332),
.B(n_316),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_352),
.A2(n_314),
.B1(n_300),
.B2(n_305),
.Y(n_369)
);

NAND2x1_ASAP7_75t_SL g388 ( 
.A(n_370),
.B(n_348),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_342),
.B(n_319),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_372),
.B(n_328),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_347),
.B(n_326),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_373),
.A2(n_335),
.B(n_349),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_374),
.A2(n_375),
.B1(n_379),
.B2(n_384),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_376),
.B(n_353),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_356),
.A2(n_333),
.B1(n_344),
.B2(n_335),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_366),
.A2(n_344),
.B1(n_334),
.B2(n_351),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_355),
.B(n_345),
.C(n_346),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_385),
.B(n_355),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_388),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_354),
.A2(n_350),
.B1(n_348),
.B2(n_322),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_389),
.B(n_370),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_390),
.B(n_393),
.C(n_395),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_391),
.B(n_392),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_385),
.B(n_362),
.C(n_367),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_382),
.B(n_372),
.C(n_371),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_382),
.B(n_360),
.C(n_363),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_381),
.A2(n_369),
.B(n_370),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_396),
.A2(n_402),
.B(n_388),
.Y(n_403)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_397),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_374),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_398),
.B(n_379),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_383),
.B(n_360),
.C(n_370),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_400),
.B(n_383),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_387),
.B(n_279),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_401),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_378),
.A2(n_348),
.B(n_290),
.Y(n_402)
);

AO21x2_ASAP7_75t_L g416 ( 
.A1(n_403),
.A2(n_386),
.B(n_384),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_399),
.A2(n_377),
.B1(n_378),
.B2(n_389),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_404),
.A2(n_412),
.B1(n_400),
.B2(n_395),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_392),
.B(n_380),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_405),
.B(n_406),
.Y(n_419)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_402),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_408),
.B(n_413),
.Y(n_414)
);

CKINVDCx14_ASAP7_75t_R g412 ( 
.A(n_394),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_408),
.A2(n_396),
.B(n_397),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_415),
.A2(n_420),
.B(n_407),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_416),
.B(n_417),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_409),
.A2(n_393),
.B(n_390),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_418),
.B(n_411),
.C(n_3),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_403),
.A2(n_376),
.B(n_375),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_410),
.B(n_9),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_421),
.B(n_410),
.Y(n_423)
);

NOR2x1_ASAP7_75t_L g422 ( 
.A(n_411),
.B(n_15),
.Y(n_422)
);

NOR2x1_ASAP7_75t_L g427 ( 
.A(n_422),
.B(n_414),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_423),
.Y(n_431)
);

OA21x2_ASAP7_75t_SL g425 ( 
.A1(n_419),
.A2(n_413),
.B(n_407),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_425),
.B(n_428),
.C(n_415),
.Y(n_429)
);

OAI211xp5_ASAP7_75t_L g430 ( 
.A1(n_426),
.A2(n_427),
.B(n_416),
.C(n_4),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_429),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_430),
.Y(n_433)
);

OAI321xp33_ASAP7_75t_L g434 ( 
.A1(n_432),
.A2(n_423),
.A3(n_431),
.B1(n_424),
.B2(n_12),
.C(n_15),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_434),
.A2(n_433),
.B(n_5),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_435),
.A2(n_11),
.B(n_1),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_436),
.B(n_11),
.Y(n_437)
);


endmodule