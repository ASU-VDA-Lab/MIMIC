module fake_ariane_1823_n_1926 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1926);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1926;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_590;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1860;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_177;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_28),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_149),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_108),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_31),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_22),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_65),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_25),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_34),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_39),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_77),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_166),
.Y(n_189)
);

BUFx10_ASAP7_75t_L g190 ( 
.A(n_6),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_129),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_47),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_54),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_133),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_29),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_29),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_97),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_117),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_87),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_142),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_32),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_5),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_96),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_37),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_7),
.Y(n_205)
);

BUFx10_ASAP7_75t_L g206 ( 
.A(n_79),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_123),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_163),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_46),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_127),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_100),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_35),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_7),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_154),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_21),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_146),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_34),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_173),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_111),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_159),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_151),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_103),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_86),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_42),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_128),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_10),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_155),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_32),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_35),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_110),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_136),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_131),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_90),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_75),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_28),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_83),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_176),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_8),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_175),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_168),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_41),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_167),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_73),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_2),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_42),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_38),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_98),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_104),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_25),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_174),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_121),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_74),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_48),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_19),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_105),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_24),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_170),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_20),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_125),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_1),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_1),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_130),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_116),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_160),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_39),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_135),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_69),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_54),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_120),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_58),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_158),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_139),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_141),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_41),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_102),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_78),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_113),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_36),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_85),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_48),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_18),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_106),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_61),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_148),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_20),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_153),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_55),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_122),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_72),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_26),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_150),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_107),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_99),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_8),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_57),
.Y(n_295)
);

BUFx10_ASAP7_75t_L g296 ( 
.A(n_134),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_36),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_94),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_70),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_13),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_30),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_19),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_52),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_52),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_15),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_30),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_114),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_118),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_64),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_76),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_66),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_13),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_112),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_164),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_26),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_0),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_60),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_165),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_44),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_169),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_92),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_15),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_144),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_49),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_0),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_143),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_88),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_65),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_115),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_18),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_40),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_59),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_24),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_81),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_132),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_16),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_59),
.Y(n_337)
);

BUFx10_ASAP7_75t_L g338 ( 
.A(n_157),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_2),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_56),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_66),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_60),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_57),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_11),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_40),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_101),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_44),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_61),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_49),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_126),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_67),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_37),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_203),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_253),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_210),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_234),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_322),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_210),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_272),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_177),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_274),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_220),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_220),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_182),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_183),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_222),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_184),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_185),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_202),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_222),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_303),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_193),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_253),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_195),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_233),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_310),
.B(n_3),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_221),
.Y(n_377)
);

NOR2xp67_ASAP7_75t_L g378 ( 
.A(n_336),
.B(n_3),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_311),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_233),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_236),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_336),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_236),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_240),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_202),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_201),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_310),
.B(n_4),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_313),
.B(n_4),
.Y(n_388)
);

INVxp67_ASAP7_75t_SL g389 ( 
.A(n_261),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_313),
.B(n_5),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_240),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_183),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_344),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_247),
.Y(n_394)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_261),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_212),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_192),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_247),
.Y(n_398)
);

NOR2xp67_ASAP7_75t_L g399 ( 
.A(n_192),
.B(n_6),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_309),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_213),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_263),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_226),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_228),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_263),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_347),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_309),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_264),
.Y(n_408)
);

NOR2xp67_ASAP7_75t_L g409 ( 
.A(n_215),
.B(n_9),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_264),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_L g411 ( 
.A(n_215),
.B(n_9),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_223),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_221),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_266),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_266),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_346),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_241),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_267),
.B(n_10),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_267),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_273),
.B(n_11),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_245),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_273),
.Y(n_422)
);

INVxp33_ASAP7_75t_SL g423 ( 
.A(n_246),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_346),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_249),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_276),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_254),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_256),
.Y(n_428)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_253),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g430 ( 
.A(n_253),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_276),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_279),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_191),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_191),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_265),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_191),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_191),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_279),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_206),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_206),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_354),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_429),
.B(n_180),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_430),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_355),
.B(n_260),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_355),
.B(n_282),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_421),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_358),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_416),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_354),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_376),
.B(n_253),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_358),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_362),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_354),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_373),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_373),
.Y(n_455)
);

CKINVDCx8_ASAP7_75t_R g456 ( 
.A(n_377),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_373),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_412),
.B(n_362),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_424),
.Y(n_459)
);

INVx6_ASAP7_75t_L g460 ( 
.A(n_412),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_363),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_363),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_366),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_366),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_370),
.Y(n_465)
);

BUFx8_ASAP7_75t_L g466 ( 
.A(n_412),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_377),
.A2(n_302),
.B1(n_332),
.B2(n_331),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_370),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_375),
.Y(n_469)
);

NAND2xp33_ASAP7_75t_L g470 ( 
.A(n_375),
.B(n_253),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_400),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_407),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_380),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_357),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_380),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_353),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_381),
.B(n_260),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_381),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_383),
.B(n_282),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_413),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_383),
.B(n_301),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_384),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_360),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_384),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_391),
.B(n_288),
.Y(n_485)
);

INVx6_ASAP7_75t_L g486 ( 
.A(n_391),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_394),
.B(n_288),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_394),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_398),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_398),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_402),
.Y(n_491)
);

AND3x2_ASAP7_75t_L g492 ( 
.A(n_387),
.B(n_337),
.C(n_301),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_402),
.B(n_337),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_405),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_405),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_408),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_408),
.Y(n_497)
);

NAND2x1_ASAP7_75t_L g498 ( 
.A(n_410),
.B(n_248),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_410),
.B(n_293),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_414),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_414),
.B(n_293),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_415),
.B(n_345),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_415),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_419),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_419),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_422),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_422),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_413),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_426),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_426),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_431),
.B(n_298),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_431),
.B(n_345),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_432),
.Y(n_513)
);

AND2x6_ASAP7_75t_L g514 ( 
.A(n_432),
.B(n_179),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_438),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_438),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_369),
.B(n_325),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_453),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_466),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_480),
.Y(n_520)
);

BUFx10_ASAP7_75t_L g521 ( 
.A(n_460),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_444),
.B(n_385),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_443),
.B(n_364),
.Y(n_523)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_464),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_453),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_464),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_449),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_464),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_464),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_460),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_464),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_466),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_483),
.B(n_367),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_464),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_453),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_458),
.B(n_389),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_453),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_474),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_467),
.A2(n_388),
.B1(n_390),
.B2(n_418),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_464),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_460),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_483),
.B(n_368),
.Y(n_542)
);

INVx5_ASAP7_75t_L g543 ( 
.A(n_514),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_464),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_510),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_510),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_460),
.Y(n_547)
);

BUFx4f_ASAP7_75t_L g548 ( 
.A(n_510),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_444),
.B(n_395),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_510),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_510),
.Y(n_551)
);

BUFx8_ASAP7_75t_SL g552 ( 
.A(n_476),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_476),
.B(n_361),
.Y(n_553)
);

OR2x6_ASAP7_75t_L g554 ( 
.A(n_498),
.B(n_378),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_443),
.B(n_372),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_510),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_466),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_442),
.B(n_423),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_483),
.B(n_374),
.Y(n_559)
);

INVxp67_ASAP7_75t_SL g560 ( 
.A(n_466),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_446),
.B(n_386),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_453),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_454),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_446),
.B(n_396),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_454),
.Y(n_565)
);

INVx8_ASAP7_75t_L g566 ( 
.A(n_517),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_444),
.B(n_397),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_481),
.B(n_397),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_458),
.B(n_365),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_510),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_474),
.B(n_356),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_510),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_480),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_454),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_508),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_466),
.Y(n_576)
);

NOR2x1p5_ASAP7_75t_L g577 ( 
.A(n_498),
.B(n_401),
.Y(n_577)
);

INVx5_ASAP7_75t_L g578 ( 
.A(n_514),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_516),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_458),
.B(n_403),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_458),
.B(n_404),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_458),
.B(n_417),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_449),
.Y(n_583)
);

AOI21x1_ASAP7_75t_L g584 ( 
.A1(n_498),
.A2(n_307),
.B(n_298),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_481),
.B(n_382),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_516),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_516),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_517),
.B(n_425),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_516),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_516),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_449),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_516),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_516),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_517),
.B(n_392),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_454),
.Y(n_595)
);

INVx1_ASAP7_75t_SL g596 ( 
.A(n_459),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_442),
.B(n_427),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_516),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_503),
.Y(n_599)
);

AND2x2_ASAP7_75t_SL g600 ( 
.A(n_470),
.B(n_194),
.Y(n_600)
);

OR2x6_ASAP7_75t_L g601 ( 
.A(n_477),
.B(n_378),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_517),
.B(n_428),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_441),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_467),
.A2(n_420),
.B1(n_409),
.B2(n_411),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_L g605 ( 
.A1(n_456),
.A2(n_305),
.B1(n_304),
.B2(n_300),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_456),
.B(n_435),
.Y(n_606)
);

AND2x6_ASAP7_75t_L g607 ( 
.A(n_463),
.B(n_307),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_454),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_455),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_456),
.B(n_359),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_504),
.B(n_433),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_450),
.A2(n_399),
.B1(n_409),
.B2(n_411),
.Y(n_612)
);

INVxp33_ASAP7_75t_SL g613 ( 
.A(n_508),
.Y(n_613)
);

NAND2xp33_ASAP7_75t_R g614 ( 
.A(n_448),
.B(n_434),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_449),
.Y(n_615)
);

INVx8_ASAP7_75t_L g616 ( 
.A(n_517),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_455),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_455),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_455),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_455),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_503),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_459),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_503),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_503),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_463),
.Y(n_625)
);

BUFx10_ASAP7_75t_L g626 ( 
.A(n_460),
.Y(n_626)
);

CKINVDCx14_ASAP7_75t_R g627 ( 
.A(n_448),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_441),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_504),
.B(n_382),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_504),
.B(n_436),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_450),
.A2(n_399),
.B1(n_439),
.B2(n_437),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_460),
.B(n_440),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_504),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_441),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_503),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_506),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_471),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_509),
.B(n_513),
.Y(n_638)
);

BUFx10_ASAP7_75t_L g639 ( 
.A(n_486),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_463),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_463),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_471),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_509),
.B(n_513),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_481),
.B(n_190),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_506),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_509),
.B(n_199),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_506),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_506),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_465),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_509),
.A2(n_209),
.B1(n_217),
.B2(n_205),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_441),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_465),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_465),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_506),
.Y(n_654)
);

CKINVDCx16_ASAP7_75t_R g655 ( 
.A(n_448),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_513),
.B(n_200),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_441),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_513),
.B(n_190),
.Y(n_658)
);

OAI22xp33_ASAP7_75t_L g659 ( 
.A1(n_472),
.A2(n_290),
.B1(n_268),
.B2(n_270),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_465),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_484),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_472),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_484),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_484),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_484),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_488),
.Y(n_666)
);

INVx4_ASAP7_75t_L g667 ( 
.A(n_486),
.Y(n_667)
);

NOR3xp33_ASAP7_75t_L g668 ( 
.A(n_445),
.B(n_187),
.C(n_186),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_447),
.B(n_326),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_447),
.B(n_248),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_624),
.B(n_451),
.Y(n_671)
);

NAND2x1_ASAP7_75t_L g672 ( 
.A(n_667),
.B(n_486),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_599),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_597),
.B(n_451),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_558),
.B(n_486),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_644),
.B(n_452),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_644),
.B(n_452),
.Y(n_677)
);

O2A1O1Ixp5_ASAP7_75t_L g678 ( 
.A1(n_638),
.A2(n_473),
.B(n_461),
.C(n_462),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_527),
.Y(n_679)
);

BUFx6f_ASAP7_75t_SL g680 ( 
.A(n_627),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_523),
.B(n_486),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_637),
.B(n_571),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_637),
.B(n_493),
.Y(n_683)
);

OAI22xp33_ASAP7_75t_L g684 ( 
.A1(n_539),
.A2(n_485),
.B1(n_445),
.B2(n_511),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_594),
.B(n_461),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_594),
.B(n_462),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_594),
.B(n_468),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_566),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_624),
.B(n_468),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_594),
.B(n_469),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_599),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_555),
.B(n_486),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_571),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_539),
.A2(n_491),
.B1(n_478),
.B2(n_482),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_527),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_583),
.Y(n_696)
);

BUFx5_ASAP7_75t_L g697 ( 
.A(n_521),
.Y(n_697)
);

AOI221xp5_ASAP7_75t_L g698 ( 
.A1(n_659),
.A2(n_258),
.B1(n_205),
.B2(n_204),
.C(n_217),
.Y(n_698)
);

A2O1A1Ixp33_ASAP7_75t_L g699 ( 
.A1(n_624),
.A2(n_491),
.B(n_469),
.C(n_473),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_624),
.B(n_475),
.Y(n_700)
);

INVxp67_ASAP7_75t_L g701 ( 
.A(n_520),
.Y(n_701)
);

INVxp67_ASAP7_75t_L g702 ( 
.A(n_520),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_635),
.B(n_475),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_583),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_596),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_635),
.B(n_478),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_580),
.B(n_581),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_583),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_538),
.B(n_493),
.Y(n_709)
);

NOR2xp67_ASAP7_75t_L g710 ( 
.A(n_642),
.B(n_479),
.Y(n_710)
);

NOR2xp67_ASAP7_75t_L g711 ( 
.A(n_622),
.B(n_479),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_621),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_536),
.B(n_566),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_635),
.B(n_636),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_SL g715 ( 
.A(n_613),
.B(n_371),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_635),
.B(n_482),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_536),
.B(n_490),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_621),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_573),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_591),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_552),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_536),
.B(n_490),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_522),
.B(n_492),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_591),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_588),
.B(n_492),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_536),
.B(n_602),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_566),
.B(n_494),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_614),
.Y(n_728)
);

NAND2xp33_ASAP7_75t_L g729 ( 
.A(n_636),
.B(n_494),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_566),
.B(n_500),
.Y(n_730)
);

INVx1_ASAP7_75t_SL g731 ( 
.A(n_573),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_582),
.B(n_500),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_615),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_566),
.B(n_505),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_636),
.B(n_505),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_636),
.B(n_507),
.Y(n_736)
);

INVx4_ASAP7_75t_L g737 ( 
.A(n_616),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_615),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_623),
.B(n_507),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_623),
.Y(n_740)
);

INVxp67_ASAP7_75t_SL g741 ( 
.A(n_633),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_645),
.B(n_488),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_616),
.B(n_488),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_615),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_616),
.B(n_488),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_645),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_616),
.B(n_485),
.Y(n_747)
);

A2O1A1Ixp33_ASAP7_75t_L g748 ( 
.A1(n_647),
.A2(n_515),
.B(n_495),
.C(n_496),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_575),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_617),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_616),
.B(n_487),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_553),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_617),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_617),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_618),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_647),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_648),
.B(n_489),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_522),
.B(n_549),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_648),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_669),
.B(n_489),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_654),
.B(n_489),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_549),
.B(n_489),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_569),
.B(n_493),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_601),
.A2(n_477),
.B1(n_502),
.B2(n_512),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_618),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_SL g766 ( 
.A1(n_553),
.A2(n_393),
.B1(n_406),
.B2(n_379),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_R g767 ( 
.A(n_655),
.B(n_487),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_633),
.B(n_495),
.Y(n_768)
);

NAND2xp33_ASAP7_75t_L g769 ( 
.A(n_643),
.B(n_495),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_660),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_585),
.B(n_512),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_601),
.A2(n_502),
.B1(n_477),
.B2(n_512),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_629),
.B(n_495),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_585),
.B(n_477),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_567),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_567),
.B(n_477),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_601),
.A2(n_502),
.B1(n_511),
.B2(n_499),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_568),
.B(n_502),
.Y(n_778)
);

O2A1O1Ixp5_ASAP7_75t_L g779 ( 
.A1(n_548),
.A2(n_515),
.B(n_496),
.C(n_497),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_660),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_646),
.B(n_656),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_601),
.A2(n_502),
.B1(n_501),
.B2(n_499),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_618),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_568),
.B(n_496),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_569),
.B(n_496),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_633),
.B(n_497),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_569),
.B(n_497),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_661),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_548),
.B(n_497),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_569),
.B(n_515),
.Y(n_790)
);

NAND2xp33_ASAP7_75t_L g791 ( 
.A(n_577),
.B(n_515),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_619),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_601),
.A2(n_501),
.B1(n_285),
.B2(n_287),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_661),
.Y(n_794)
);

INVxp67_ASAP7_75t_L g795 ( 
.A(n_662),
.Y(n_795)
);

NAND2xp33_ASAP7_75t_L g796 ( 
.A(n_577),
.B(n_514),
.Y(n_796)
);

NOR2xp67_ASAP7_75t_L g797 ( 
.A(n_632),
.B(n_271),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_658),
.B(n_278),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_670),
.B(n_320),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_548),
.A2(n_470),
.B(n_271),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_554),
.A2(n_320),
.B1(n_321),
.B2(n_251),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_554),
.A2(n_321),
.B1(n_243),
.B2(n_242),
.Y(n_802)
);

INVx8_ASAP7_75t_L g803 ( 
.A(n_554),
.Y(n_803)
);

NAND2xp33_ASAP7_75t_L g804 ( 
.A(n_519),
.B(n_514),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_665),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_655),
.Y(n_806)
);

AO22x2_ASAP7_75t_L g807 ( 
.A1(n_611),
.A2(n_186),
.B1(n_187),
.B2(n_349),
.Y(n_807)
);

NAND2x1p5_ASAP7_75t_L g808 ( 
.A(n_519),
.B(n_223),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_665),
.B(n_196),
.Y(n_809)
);

AND2x6_ASAP7_75t_SL g810 ( 
.A(n_554),
.B(n_196),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_554),
.B(n_204),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_600),
.B(n_209),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_625),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_630),
.Y(n_814)
);

BUFx6f_ASAP7_75t_SL g815 ( 
.A(n_607),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_600),
.B(n_625),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_619),
.Y(n_817)
);

BUFx5_ASAP7_75t_L g818 ( 
.A(n_521),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_524),
.B(n_194),
.Y(n_819)
);

NOR2x1p5_ASAP7_75t_L g820 ( 
.A(n_560),
.B(n_280),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_667),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_600),
.B(n_224),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_640),
.B(n_641),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_524),
.B(n_211),
.Y(n_824)
);

BUFx5_ASAP7_75t_L g825 ( 
.A(n_521),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_561),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_524),
.B(n_252),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_603),
.B(n_252),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_640),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_603),
.B(n_179),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_641),
.B(n_224),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_649),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_564),
.B(n_297),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_649),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_603),
.B(n_179),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_604),
.A2(n_227),
.B1(n_237),
.B2(n_232),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_652),
.B(n_229),
.Y(n_837)
);

OAI22xp33_ASAP7_75t_L g838 ( 
.A1(n_604),
.A2(n_244),
.B1(n_238),
.B2(n_235),
.Y(n_838)
);

INVx1_ASAP7_75t_SL g839 ( 
.A(n_731),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_779),
.A2(n_529),
.B(n_528),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_701),
.B(n_533),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_673),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_688),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_758),
.B(n_674),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_758),
.B(n_631),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_769),
.A2(n_529),
.B(n_528),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_691),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_713),
.A2(n_542),
.B1(n_559),
.B2(n_606),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_712),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_714),
.A2(n_534),
.B(n_531),
.Y(n_850)
);

OAI21xp5_ASAP7_75t_L g851 ( 
.A1(n_714),
.A2(n_534),
.B(n_531),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_789),
.A2(n_544),
.B(n_540),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_675),
.B(n_668),
.Y(n_853)
);

CKINVDCx20_ASAP7_75t_R g854 ( 
.A(n_721),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_718),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_747),
.A2(n_544),
.B(n_540),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_747),
.A2(n_546),
.B(n_545),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_702),
.B(n_610),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_675),
.B(n_532),
.Y(n_859)
);

NAND2x1p5_ASAP7_75t_L g860 ( 
.A(n_737),
.B(n_532),
.Y(n_860)
);

AO21x1_ASAP7_75t_L g861 ( 
.A1(n_684),
.A2(n_546),
.B(n_545),
.Y(n_861)
);

AO21x1_ASAP7_75t_L g862 ( 
.A1(n_684),
.A2(n_551),
.B(n_550),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_719),
.B(n_605),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_L g864 ( 
.A1(n_678),
.A2(n_551),
.B(n_550),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_688),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_688),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_707),
.B(n_557),
.Y(n_867)
);

NOR3xp33_ASAP7_75t_L g868 ( 
.A(n_693),
.B(n_235),
.C(n_229),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_740),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_707),
.B(n_557),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_715),
.B(n_795),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_751),
.A2(n_579),
.B(n_556),
.Y(n_872)
);

O2A1O1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_751),
.A2(n_666),
.B(n_664),
.C(n_663),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_676),
.B(n_576),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_789),
.A2(n_579),
.B(n_556),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_681),
.A2(n_587),
.B(n_586),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_SL g877 ( 
.A1(n_815),
.A2(n_576),
.B(n_541),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_688),
.B(n_639),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_737),
.B(n_639),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_727),
.A2(n_667),
.B1(n_570),
.B2(n_526),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_681),
.A2(n_587),
.B(n_586),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_692),
.A2(n_590),
.B(n_589),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_692),
.A2(n_590),
.B(n_589),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_677),
.B(n_710),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_749),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_773),
.A2(n_593),
.B(n_592),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_699),
.A2(n_593),
.B(n_592),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_746),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_682),
.B(n_667),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_767),
.B(n_650),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_729),
.A2(n_598),
.B(n_570),
.Y(n_891)
);

AO21x1_ASAP7_75t_L g892 ( 
.A1(n_799),
.A2(n_598),
.B(n_584),
.Y(n_892)
);

O2A1O1Ixp33_ASAP7_75t_SL g893 ( 
.A1(n_748),
.A2(n_572),
.B(n_570),
.C(n_526),
.Y(n_893)
);

BUFx5_ASAP7_75t_L g894 ( 
.A(n_756),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_803),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_767),
.B(n_639),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_742),
.A2(n_570),
.B(n_526),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_705),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_742),
.A2(n_572),
.B(n_526),
.Y(n_899)
);

O2A1O1Ixp33_ASAP7_75t_SL g900 ( 
.A1(n_757),
.A2(n_572),
.B(n_664),
.C(n_663),
.Y(n_900)
);

INVxp67_ASAP7_75t_SL g901 ( 
.A(n_741),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_763),
.B(n_530),
.Y(n_902)
);

NOR3xp33_ASAP7_75t_L g903 ( 
.A(n_833),
.B(n_698),
.C(n_806),
.Y(n_903)
);

AOI21xp33_ASAP7_75t_L g904 ( 
.A1(n_833),
.A2(n_612),
.B(n_652),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_711),
.B(n_639),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_763),
.B(n_521),
.Y(n_906)
);

NAND2x1p5_ASAP7_75t_L g907 ( 
.A(n_726),
.B(n_686),
.Y(n_907)
);

O2A1O1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_775),
.A2(n_666),
.B(n_653),
.C(n_619),
.Y(n_908)
);

A2O1A1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_732),
.A2(n_653),
.B(n_620),
.C(n_518),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_757),
.A2(n_572),
.B(n_657),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_803),
.Y(n_911)
);

NOR2xp67_ASAP7_75t_L g912 ( 
.A(n_728),
.B(n_826),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_814),
.B(n_518),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_723),
.B(n_626),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_771),
.B(n_525),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_761),
.A2(n_657),
.B(n_620),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_761),
.A2(n_786),
.B(n_768),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_768),
.A2(n_657),
.B(n_620),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_776),
.B(n_525),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_778),
.B(n_774),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_709),
.B(n_190),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_781),
.B(n_535),
.Y(n_922)
);

AO21x1_ASAP7_75t_L g923 ( 
.A1(n_828),
.A2(n_584),
.B(n_537),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_725),
.B(n_535),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_803),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_743),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_717),
.B(n_537),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_679),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_671),
.A2(n_563),
.B(n_562),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_722),
.B(n_562),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_732),
.B(n_563),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_725),
.A2(n_607),
.B1(n_574),
.B2(n_609),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_671),
.A2(n_541),
.B(n_530),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_683),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_689),
.A2(n_541),
.B(n_530),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_820),
.Y(n_936)
);

AOI21x1_ASAP7_75t_L g937 ( 
.A1(n_739),
.A2(n_574),
.B(n_565),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_759),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_L g939 ( 
.A1(n_723),
.A2(n_607),
.B1(n_609),
.B2(n_608),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_689),
.A2(n_547),
.B(n_603),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_786),
.A2(n_595),
.B(n_565),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_798),
.B(n_595),
.Y(n_942)
);

OAI21xp33_ASAP7_75t_L g943 ( 
.A1(n_784),
.A2(n_316),
.B(n_312),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_764),
.B(n_626),
.Y(n_944)
);

AOI21x1_ASAP7_75t_L g945 ( 
.A1(n_739),
.A2(n_608),
.B(n_244),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_770),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_685),
.B(n_607),
.Y(n_947)
);

OAI22xp5_ASAP7_75t_L g948 ( 
.A1(n_730),
.A2(n_547),
.B1(n_324),
.B2(n_328),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_687),
.B(n_607),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_690),
.B(n_607),
.Y(n_950)
);

O2A1O1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_785),
.A2(n_238),
.B(n_258),
.C(n_349),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_745),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_780),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_700),
.A2(n_607),
.B(n_547),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_762),
.B(n_603),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_694),
.B(n_603),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_787),
.B(n_628),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_788),
.Y(n_958)
);

AO21x1_ASAP7_75t_L g959 ( 
.A1(n_828),
.A2(n_348),
.B(n_317),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_772),
.B(n_626),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_790),
.B(n_777),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_734),
.A2(n_339),
.B1(n_333),
.B2(n_340),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_802),
.B(n_626),
.Y(n_963)
);

BUFx4f_ASAP7_75t_L g964 ( 
.A(n_808),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_782),
.B(n_628),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_700),
.A2(n_651),
.B(n_634),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_703),
.A2(n_651),
.B(n_634),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_811),
.B(n_628),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_797),
.B(n_628),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_703),
.A2(n_514),
.B(n_578),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_798),
.B(n_628),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_706),
.A2(n_514),
.B(n_578),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_794),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_760),
.B(n_628),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_838),
.B(n_634),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_838),
.B(n_634),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_812),
.B(n_634),
.Y(n_977)
);

INVx4_ASAP7_75t_L g978 ( 
.A(n_680),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_706),
.A2(n_514),
.B(n_543),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_821),
.B(n_281),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_836),
.A2(n_352),
.B1(n_351),
.B2(n_343),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_716),
.A2(n_651),
.B(n_634),
.Y(n_982)
);

O2A1O1Ixp33_ASAP7_75t_SL g983 ( 
.A1(n_716),
.A2(n_317),
.B(n_348),
.C(n_342),
.Y(n_983)
);

AND2x6_ASAP7_75t_L g984 ( 
.A(n_816),
.B(n_651),
.Y(n_984)
);

AOI21x1_ASAP7_75t_L g985 ( 
.A1(n_735),
.A2(n_319),
.B(n_281),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_735),
.A2(n_651),
.B(n_578),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_736),
.A2(n_651),
.B(n_441),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_801),
.B(n_341),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_807),
.B(n_190),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_805),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_736),
.A2(n_441),
.B(n_457),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_791),
.A2(n_294),
.B(n_319),
.C(n_306),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_793),
.A2(n_306),
.B(n_342),
.C(n_330),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_809),
.A2(n_822),
.B(n_750),
.C(n_753),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_823),
.A2(n_578),
.B(n_543),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_766),
.B(n_283),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_754),
.A2(n_578),
.B(n_543),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_755),
.A2(n_578),
.B(n_543),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_819),
.A2(n_457),
.B(n_441),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_821),
.A2(n_315),
.B1(n_294),
.B2(n_330),
.Y(n_1000)
);

OAI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_819),
.A2(n_514),
.B(n_543),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_672),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_697),
.B(n_283),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_765),
.A2(n_783),
.B(n_792),
.C(n_817),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_752),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_695),
.A2(n_543),
.B(n_257),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_680),
.B(n_283),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_696),
.A2(n_178),
.B(n_181),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_704),
.A2(n_275),
.B(n_225),
.Y(n_1009)
);

CKINVDCx10_ASAP7_75t_R g1010 ( 
.A(n_815),
.Y(n_1010)
);

AO21x1_ASAP7_75t_L g1011 ( 
.A1(n_824),
.A2(n_295),
.B(n_457),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_807),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_807),
.B(n_283),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_808),
.B(n_325),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_813),
.B(n_325),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_708),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_824),
.A2(n_457),
.B(n_325),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_829),
.B(n_325),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_832),
.B(n_325),
.Y(n_1019)
);

NOR3xp33_ASAP7_75t_L g1020 ( 
.A(n_796),
.B(n_327),
.C(n_231),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_834),
.B(n_188),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_810),
.B(n_206),
.Y(n_1022)
);

O2A1O1Ixp5_ASAP7_75t_L g1023 ( 
.A1(n_827),
.A2(n_514),
.B(n_338),
.C(n_296),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_827),
.A2(n_269),
.B(n_214),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_720),
.A2(n_277),
.B(n_216),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_724),
.B(n_189),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_733),
.B(n_197),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_844),
.A2(n_818),
.B(n_697),
.Y(n_1028)
);

BUFx2_ASAP7_75t_L g1029 ( 
.A(n_839),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_842),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_934),
.B(n_921),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_863),
.B(n_738),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_871),
.A2(n_804),
.B1(n_831),
.B2(n_837),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_895),
.B(n_744),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_895),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_898),
.Y(n_1036)
);

INVx2_ASAP7_75t_SL g1037 ( 
.A(n_1010),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_847),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_845),
.B(n_800),
.Y(n_1039)
);

CKINVDCx16_ASAP7_75t_R g1040 ( 
.A(n_854),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_849),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_890),
.B(n_206),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_928),
.Y(n_1043)
);

INVxp67_ASAP7_75t_L g1044 ( 
.A(n_885),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_853),
.A2(n_835),
.B(n_830),
.C(n_259),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_859),
.A2(n_825),
.B(n_818),
.Y(n_1046)
);

BUFx5_ASAP7_75t_L g1047 ( 
.A(n_984),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_867),
.B(n_697),
.Y(n_1048)
);

NOR3xp33_ASAP7_75t_SL g1049 ( 
.A(n_962),
.B(n_289),
.C(n_207),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_855),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_920),
.B(n_830),
.Y(n_1051)
);

INVx4_ASAP7_75t_L g1052 ( 
.A(n_895),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_1005),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_869),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_884),
.B(n_835),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_996),
.B(n_296),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_978),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_888),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_993),
.A2(n_259),
.B(n_262),
.C(n_350),
.Y(n_1059)
);

INVx2_ASAP7_75t_SL g1060 ( 
.A(n_978),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_870),
.B(n_697),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_903),
.A2(n_262),
.B(n_350),
.C(n_16),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_889),
.B(n_697),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_961),
.A2(n_825),
.B1(n_818),
.B2(n_697),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_841),
.B(n_818),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_SL g1066 ( 
.A1(n_971),
.A2(n_825),
.B(n_818),
.C(n_17),
.Y(n_1066)
);

AND2x6_ASAP7_75t_SL g1067 ( 
.A(n_1007),
.B(n_12),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_924),
.B(n_818),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_874),
.A2(n_825),
.B1(n_291),
.B2(n_335),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_942),
.A2(n_179),
.B(n_329),
.C(n_250),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_938),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_848),
.B(n_825),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_911),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_901),
.A2(n_825),
.B1(n_286),
.B2(n_334),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_858),
.B(n_296),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_951),
.A2(n_179),
.B(n_250),
.C(n_329),
.Y(n_1076)
);

INVx2_ASAP7_75t_SL g1077 ( 
.A(n_964),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_946),
.B(n_12),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_926),
.B(n_457),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_982),
.A2(n_457),
.B(n_329),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_907),
.B(n_296),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_953),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_1016),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_958),
.A2(n_255),
.B1(n_198),
.B2(n_323),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_973),
.A2(n_990),
.B1(n_956),
.B2(n_976),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_926),
.B(n_457),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_974),
.A2(n_284),
.B(n_218),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1012),
.B(n_14),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_975),
.A2(n_179),
.B(n_329),
.C(n_250),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_919),
.A2(n_208),
.B1(n_219),
.B2(n_230),
.Y(n_1090)
);

O2A1O1Ixp33_ASAP7_75t_SL g1091 ( 
.A1(n_909),
.A2(n_14),
.B(n_17),
.C(n_21),
.Y(n_1091)
);

BUFx12f_ASAP7_75t_L g1092 ( 
.A(n_936),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_980),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_907),
.B(n_338),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_866),
.Y(n_1095)
);

OAI21xp33_ASAP7_75t_L g1096 ( 
.A1(n_981),
.A2(n_239),
.B(n_318),
.Y(n_1096)
);

BUFx3_ASAP7_75t_L g1097 ( 
.A(n_911),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_904),
.A2(n_329),
.B(n_250),
.C(n_314),
.Y(n_1098)
);

AO21x2_ASAP7_75t_L g1099 ( 
.A1(n_861),
.A2(n_338),
.B(n_329),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_955),
.A2(n_308),
.B(n_299),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_902),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_926),
.B(n_250),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_980),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_876),
.A2(n_292),
.B(n_250),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_881),
.A2(n_71),
.B(n_172),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_915),
.Y(n_1106)
);

OAI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_917),
.A2(n_338),
.B(n_23),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_911),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_985),
.Y(n_1109)
);

AOI21x1_ASAP7_75t_L g1110 ( 
.A1(n_862),
.A2(n_171),
.B(n_162),
.Y(n_1110)
);

O2A1O1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_868),
.A2(n_22),
.B(n_23),
.C(n_27),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_989),
.B(n_27),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_866),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_902),
.B(n_922),
.Y(n_1114)
);

NOR3xp33_ASAP7_75t_L g1115 ( 
.A(n_943),
.B(n_988),
.C(n_1000),
.Y(n_1115)
);

OR2x6_ASAP7_75t_L g1116 ( 
.A(n_925),
.B(n_31),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_866),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_925),
.B(n_33),
.Y(n_1118)
);

AOI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1022),
.A2(n_944),
.B1(n_960),
.B2(n_914),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_SL g1120 ( 
.A1(n_1013),
.A2(n_33),
.B1(n_38),
.B2(n_43),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_882),
.A2(n_80),
.B(n_156),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_883),
.A2(n_161),
.B(n_145),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_913),
.B(n_43),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_939),
.B(n_931),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_927),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_964),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_R g1127 ( 
.A(n_925),
.B(n_140),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_937),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_992),
.A2(n_45),
.B(n_46),
.C(n_47),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_930),
.Y(n_1130)
);

INVx4_ASAP7_75t_L g1131 ( 
.A(n_843),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_912),
.B(n_45),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_952),
.B(n_50),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_945),
.Y(n_1134)
);

O2A1O1Ixp33_ASAP7_75t_SL g1135 ( 
.A1(n_1003),
.A2(n_50),
.B(n_51),
.C(n_53),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_894),
.Y(n_1136)
);

AOI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_896),
.A2(n_51),
.B1(n_53),
.B2(n_55),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_965),
.A2(n_56),
.B1(n_58),
.B2(n_62),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_900),
.A2(n_91),
.B(n_137),
.Y(n_1139)
);

AOI21x1_ASAP7_75t_L g1140 ( 
.A1(n_1015),
.A2(n_1019),
.B(n_1018),
.Y(n_1140)
);

O2A1O1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_983),
.A2(n_62),
.B(n_63),
.C(n_64),
.Y(n_1141)
);

AO21x1_ASAP7_75t_L g1142 ( 
.A1(n_994),
.A2(n_93),
.B(n_124),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_957),
.A2(n_89),
.B(n_119),
.Y(n_1143)
);

AOI22xp33_ASAP7_75t_L g1144 ( 
.A1(n_947),
.A2(n_63),
.B1(n_67),
.B2(n_68),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_894),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_886),
.A2(n_82),
.B(n_84),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1021),
.B(n_68),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_856),
.A2(n_95),
.B(n_109),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_843),
.B(n_138),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_865),
.B(n_906),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_952),
.B(n_894),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_857),
.A2(n_872),
.B(n_982),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_952),
.B(n_894),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_917),
.A2(n_977),
.B(n_873),
.Y(n_1154)
);

OR2x2_ASAP7_75t_L g1155 ( 
.A(n_1026),
.B(n_1027),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_949),
.B(n_950),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_SL g1157 ( 
.A(n_860),
.B(n_865),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_846),
.A2(n_967),
.B(n_966),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_846),
.A2(n_910),
.B(n_918),
.Y(n_1159)
);

O2A1O1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_948),
.A2(n_893),
.B(n_908),
.C(n_1025),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_894),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_894),
.B(n_968),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_910),
.A2(n_918),
.B(n_852),
.Y(n_1163)
);

CKINVDCx8_ASAP7_75t_R g1164 ( 
.A(n_984),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_932),
.B(n_984),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_984),
.B(n_1004),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_984),
.B(n_1024),
.Y(n_1167)
);

INVx1_ASAP7_75t_SL g1168 ( 
.A(n_1014),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_851),
.B(n_954),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_929),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1002),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_969),
.B(n_1002),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_860),
.A2(n_963),
.B1(n_879),
.B2(n_905),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_850),
.A2(n_916),
.B(n_899),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_852),
.A2(n_875),
.B(n_916),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_850),
.B(n_941),
.Y(n_1176)
);

OAI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_897),
.A2(n_899),
.B(n_941),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_897),
.B(n_1020),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_877),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_891),
.A2(n_840),
.B(n_940),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_891),
.A2(n_887),
.B1(n_880),
.B2(n_878),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_959),
.Y(n_1182)
);

OA21x2_ASAP7_75t_L g1183 ( 
.A1(n_864),
.A2(n_1017),
.B(n_999),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_987),
.B(n_1009),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1023),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_1011),
.Y(n_1186)
);

AOI21xp33_ASAP7_75t_L g1187 ( 
.A1(n_1075),
.A2(n_1056),
.B(n_1062),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1080),
.A2(n_999),
.B(n_1017),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1159),
.A2(n_1163),
.B(n_1158),
.Y(n_1189)
);

AO32x2_ASAP7_75t_L g1190 ( 
.A1(n_1085),
.A2(n_892),
.A3(n_923),
.B1(n_987),
.B2(n_991),
.Y(n_1190)
);

OAI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1107),
.A2(n_933),
.B(n_935),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1063),
.A2(n_986),
.B(n_991),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1152),
.A2(n_997),
.B(n_998),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1068),
.A2(n_1006),
.B(n_972),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1064),
.A2(n_970),
.B(n_979),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1075),
.B(n_1008),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1028),
.A2(n_1046),
.B(n_1048),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1042),
.B(n_1001),
.Y(n_1198)
);

NOR4xp25_ASAP7_75t_L g1199 ( 
.A(n_1129),
.B(n_995),
.C(n_1111),
.D(n_1141),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_1040),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1032),
.B(n_1031),
.Y(n_1201)
);

O2A1O1Ixp5_ASAP7_75t_L g1202 ( 
.A1(n_1177),
.A2(n_1142),
.B(n_1174),
.C(n_1123),
.Y(n_1202)
);

CKINVDCx9p33_ASAP7_75t_R g1203 ( 
.A(n_1053),
.Y(n_1203)
);

AO32x2_ASAP7_75t_L g1204 ( 
.A1(n_1120),
.A2(n_1138),
.A3(n_1181),
.B1(n_1173),
.B2(n_1131),
.Y(n_1204)
);

INVxp67_ASAP7_75t_L g1205 ( 
.A(n_1029),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1175),
.A2(n_1180),
.B(n_1176),
.Y(n_1206)
);

BUFx12f_ASAP7_75t_L g1207 ( 
.A(n_1037),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1140),
.A2(n_1184),
.B(n_1154),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1048),
.A2(n_1061),
.B(n_1072),
.Y(n_1209)
);

O2A1O1Ixp33_ASAP7_75t_SL g1210 ( 
.A1(n_1065),
.A2(n_1066),
.B(n_1061),
.C(n_1169),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1044),
.B(n_1101),
.Y(n_1211)
);

NOR2xp67_ASAP7_75t_L g1212 ( 
.A(n_1179),
.B(n_1131),
.Y(n_1212)
);

OAI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1112),
.A2(n_1116),
.B1(n_1119),
.B2(n_1103),
.Y(n_1213)
);

NOR2xp67_ASAP7_75t_SL g1214 ( 
.A(n_1092),
.B(n_1164),
.Y(n_1214)
);

CKINVDCx11_ASAP7_75t_R g1215 ( 
.A(n_1067),
.Y(n_1215)
);

OA21x2_ASAP7_75t_L g1216 ( 
.A1(n_1089),
.A2(n_1098),
.B(n_1070),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1030),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1162),
.A2(n_1169),
.B(n_1178),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1160),
.A2(n_1153),
.B(n_1151),
.Y(n_1219)
);

AO32x2_ASAP7_75t_L g1220 ( 
.A1(n_1099),
.A2(n_1090),
.A3(n_1069),
.B1(n_1084),
.B2(n_1091),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1044),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1151),
.A2(n_1153),
.B(n_1039),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1123),
.A2(n_1032),
.B1(n_1155),
.B2(n_1114),
.Y(n_1223)
);

CKINVDCx20_ASAP7_75t_R g1224 ( 
.A(n_1057),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1156),
.A2(n_1066),
.B(n_1165),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1038),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_1036),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1156),
.A2(n_1167),
.B(n_1145),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1128),
.A2(n_1139),
.B(n_1166),
.Y(n_1229)
);

AOI31xp67_ASAP7_75t_L g1230 ( 
.A1(n_1185),
.A2(n_1109),
.A3(n_1134),
.B(n_1172),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1060),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1106),
.B(n_1125),
.Y(n_1232)
);

A2O1A1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1115),
.A2(n_1147),
.B(n_1051),
.C(n_1081),
.Y(n_1233)
);

CKINVDCx11_ASAP7_75t_R g1234 ( 
.A(n_1116),
.Y(n_1234)
);

AOI221x1_ASAP7_75t_L g1235 ( 
.A1(n_1098),
.A2(n_1115),
.B1(n_1129),
.B2(n_1070),
.C(n_1045),
.Y(n_1235)
);

AOI221x1_ASAP7_75t_L g1236 ( 
.A1(n_1045),
.A2(n_1089),
.B1(n_1076),
.B2(n_1182),
.C(n_1088),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1136),
.A2(n_1161),
.B(n_1148),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1041),
.Y(n_1238)
);

BUFx10_ASAP7_75t_L g1239 ( 
.A(n_1118),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1051),
.A2(n_1121),
.B(n_1122),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1105),
.A2(n_1146),
.B(n_1170),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1050),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1054),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1058),
.Y(n_1244)
);

AOI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1110),
.A2(n_1102),
.B(n_1172),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1101),
.B(n_1093),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1144),
.A2(n_1124),
.B1(n_1116),
.B2(n_1049),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_1035),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1071),
.Y(n_1249)
);

AO31x2_ASAP7_75t_L g1250 ( 
.A1(n_1055),
.A2(n_1104),
.A3(n_1130),
.B(n_1083),
.Y(n_1250)
);

INVxp67_ASAP7_75t_L g1251 ( 
.A(n_1082),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1081),
.B(n_1094),
.Y(n_1252)
);

INVx4_ASAP7_75t_L g1253 ( 
.A(n_1035),
.Y(n_1253)
);

NOR4xp25_ASAP7_75t_L g1254 ( 
.A(n_1144),
.B(n_1091),
.C(n_1059),
.D(n_1135),
.Y(n_1254)
);

BUFx4_ASAP7_75t_SL g1255 ( 
.A(n_1126),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1094),
.B(n_1077),
.Y(n_1256)
);

AO32x2_ASAP7_75t_L g1257 ( 
.A1(n_1099),
.A2(n_1052),
.A3(n_1074),
.B1(n_1183),
.B2(n_1135),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1183),
.A2(n_1143),
.B(n_1086),
.Y(n_1258)
);

AOI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1118),
.A2(n_1133),
.B1(n_1096),
.B2(n_1137),
.Y(n_1259)
);

NOR2xp67_ASAP7_75t_L g1260 ( 
.A(n_1095),
.B(n_1113),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1171),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_SL g1262 ( 
.A1(n_1078),
.A2(n_1100),
.B(n_1087),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1097),
.Y(n_1263)
);

O2A1O1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1133),
.A2(n_1049),
.B(n_1132),
.C(n_1150),
.Y(n_1264)
);

NOR2xp67_ASAP7_75t_SL g1265 ( 
.A(n_1035),
.B(n_1073),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_1108),
.Y(n_1266)
);

AO21x2_ASAP7_75t_L g1267 ( 
.A1(n_1079),
.A2(n_1086),
.B(n_1033),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1034),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1052),
.B(n_1035),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1034),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1073),
.B(n_1150),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1079),
.A2(n_1157),
.B(n_1149),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1149),
.A2(n_1168),
.B(n_1117),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1073),
.B(n_1095),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1073),
.B(n_1113),
.Y(n_1275)
);

AO21x1_ASAP7_75t_L g1276 ( 
.A1(n_1047),
.A2(n_1186),
.B(n_1127),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_1117),
.B(n_1127),
.Y(n_1277)
);

AO31x2_ASAP7_75t_L g1278 ( 
.A1(n_1186),
.A2(n_1098),
.A3(n_1089),
.B(n_1128),
.Y(n_1278)
);

NOR2x1_ASAP7_75t_SL g1279 ( 
.A(n_1047),
.B(n_1116),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1047),
.Y(n_1280)
);

OR2x6_ASAP7_75t_L g1281 ( 
.A(n_1047),
.B(n_803),
.Y(n_1281)
);

INVx4_ASAP7_75t_L g1282 ( 
.A(n_1047),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1047),
.A2(n_1063),
.B(n_1068),
.Y(n_1283)
);

O2A1O1Ixp33_ASAP7_75t_SL g1284 ( 
.A1(n_1065),
.A2(n_844),
.B(n_853),
.C(n_1066),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1042),
.B(n_693),
.Y(n_1285)
);

AO21x2_ASAP7_75t_L g1286 ( 
.A1(n_1098),
.A2(n_1140),
.B(n_1045),
.Y(n_1286)
);

INVx2_ASAP7_75t_SL g1287 ( 
.A(n_1036),
.Y(n_1287)
);

OA21x2_ASAP7_75t_L g1288 ( 
.A1(n_1177),
.A2(n_1159),
.B(n_1163),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1080),
.A2(n_1159),
.B(n_1163),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1030),
.Y(n_1290)
);

AOI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1075),
.A2(n_863),
.B1(n_903),
.B2(n_1123),
.Y(n_1291)
);

OAI22x1_ASAP7_75t_L g1292 ( 
.A1(n_1075),
.A2(n_553),
.B1(n_1056),
.B2(n_996),
.Y(n_1292)
);

A2O1A1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1075),
.A2(n_844),
.B(n_1107),
.C(n_707),
.Y(n_1293)
);

INVx5_ASAP7_75t_SL g1294 ( 
.A(n_1116),
.Y(n_1294)
);

AO32x2_ASAP7_75t_L g1295 ( 
.A1(n_1085),
.A2(n_1012),
.A3(n_1120),
.B1(n_1138),
.B2(n_1181),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1080),
.A2(n_1159),
.B(n_1163),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1063),
.A2(n_1068),
.B(n_1064),
.Y(n_1297)
);

INVx5_ASAP7_75t_L g1298 ( 
.A(n_1116),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_SL g1299 ( 
.A(n_1032),
.B(n_867),
.Y(n_1299)
);

OA21x2_ASAP7_75t_L g1300 ( 
.A1(n_1177),
.A2(n_1159),
.B(n_1163),
.Y(n_1300)
);

AO31x2_ASAP7_75t_L g1301 ( 
.A1(n_1098),
.A2(n_1089),
.A3(n_1128),
.B(n_861),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1075),
.A2(n_844),
.B1(n_863),
.B2(n_853),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1040),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1080),
.A2(n_1159),
.B(n_1163),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1101),
.B(n_895),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1075),
.B(n_844),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1080),
.A2(n_1159),
.B(n_1163),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_1040),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1063),
.A2(n_1068),
.B(n_1064),
.Y(n_1309)
);

INVx3_ASAP7_75t_SL g1310 ( 
.A(n_1040),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1043),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1030),
.Y(n_1312)
);

OR2x6_ASAP7_75t_L g1313 ( 
.A(n_1116),
.B(n_803),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1063),
.A2(n_1068),
.B(n_1064),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1043),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1075),
.A2(n_766),
.B1(n_996),
.B2(n_553),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1075),
.B(n_553),
.Y(n_1317)
);

O2A1O1Ixp33_ASAP7_75t_SL g1318 ( 
.A1(n_1065),
.A2(n_844),
.B(n_853),
.C(n_1066),
.Y(n_1318)
);

AO31x2_ASAP7_75t_L g1319 ( 
.A1(n_1098),
.A2(n_1089),
.A3(n_1128),
.B(n_861),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1075),
.A2(n_766),
.B1(n_996),
.B2(n_553),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1063),
.A2(n_1068),
.B(n_1064),
.Y(n_1321)
);

OAI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1107),
.A2(n_844),
.B(n_1156),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1107),
.A2(n_844),
.B(n_1156),
.Y(n_1323)
);

AO31x2_ASAP7_75t_L g1324 ( 
.A1(n_1098),
.A2(n_1089),
.A3(n_1128),
.B(n_861),
.Y(n_1324)
);

OAI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1075),
.A2(n_715),
.B1(n_539),
.B2(n_476),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_SL g1326 ( 
.A1(n_1107),
.A2(n_844),
.B(n_867),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1043),
.Y(n_1327)
);

AO32x2_ASAP7_75t_L g1328 ( 
.A1(n_1085),
.A2(n_1012),
.A3(n_1120),
.B1(n_1138),
.B2(n_1181),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_SL g1329 ( 
.A(n_1032),
.B(n_867),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1063),
.A2(n_1068),
.B(n_1064),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1063),
.A2(n_1068),
.B(n_1064),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1063),
.A2(n_1068),
.B(n_1064),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1063),
.A2(n_1068),
.B(n_1064),
.Y(n_1333)
);

A2O1A1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1075),
.A2(n_844),
.B(n_1107),
.C(n_707),
.Y(n_1334)
);

A2O1A1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1075),
.A2(n_844),
.B(n_1107),
.C(n_707),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1075),
.A2(n_766),
.B1(n_996),
.B2(n_553),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1063),
.A2(n_1068),
.B(n_1064),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1042),
.B(n_693),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1030),
.Y(n_1339)
);

AO31x2_ASAP7_75t_L g1340 ( 
.A1(n_1098),
.A2(n_1089),
.A3(n_1128),
.B(n_861),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1075),
.B(n_553),
.Y(n_1341)
);

O2A1O1Ixp33_ASAP7_75t_SL g1342 ( 
.A1(n_1065),
.A2(n_844),
.B(n_853),
.C(n_1066),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1063),
.A2(n_1068),
.B(n_1064),
.Y(n_1343)
);

OAI21xp33_ASAP7_75t_L g1344 ( 
.A1(n_1075),
.A2(n_853),
.B(n_844),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1075),
.B(n_844),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1063),
.A2(n_1068),
.B(n_1064),
.Y(n_1346)
);

A2O1A1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1075),
.A2(n_844),
.B(n_1107),
.C(n_707),
.Y(n_1347)
);

AOI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1317),
.A2(n_1341),
.B1(n_1291),
.B2(n_1325),
.Y(n_1348)
);

CKINVDCx20_ASAP7_75t_R g1349 ( 
.A(n_1224),
.Y(n_1349)
);

CKINVDCx6p67_ASAP7_75t_R g1350 ( 
.A(n_1310),
.Y(n_1350)
);

AOI21xp33_ASAP7_75t_L g1351 ( 
.A1(n_1291),
.A2(n_1302),
.B(n_1292),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1227),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1217),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1288),
.Y(n_1354)
);

CKINVDCx20_ASAP7_75t_R g1355 ( 
.A(n_1203),
.Y(n_1355)
);

CKINVDCx20_ASAP7_75t_R g1356 ( 
.A(n_1200),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1316),
.A2(n_1320),
.B1(n_1336),
.B2(n_1344),
.Y(n_1357)
);

CKINVDCx11_ASAP7_75t_R g1358 ( 
.A(n_1207),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1226),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1306),
.B(n_1345),
.Y(n_1360)
);

INVx4_ASAP7_75t_L g1361 ( 
.A(n_1266),
.Y(n_1361)
);

INVx6_ASAP7_75t_L g1362 ( 
.A(n_1239),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_SL g1363 ( 
.A1(n_1298),
.A2(n_1247),
.B1(n_1294),
.B2(n_1252),
.Y(n_1363)
);

AOI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1344),
.A2(n_1213),
.B1(n_1223),
.B2(n_1338),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1293),
.A2(n_1347),
.B1(n_1335),
.B2(n_1334),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1285),
.B(n_1201),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1187),
.A2(n_1234),
.B1(n_1323),
.B2(n_1322),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1238),
.Y(n_1368)
);

BUFx10_ASAP7_75t_L g1369 ( 
.A(n_1303),
.Y(n_1369)
);

OAI21xp33_ASAP7_75t_SL g1370 ( 
.A1(n_1322),
.A2(n_1323),
.B(n_1326),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1298),
.A2(n_1259),
.B1(n_1329),
.B2(n_1299),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1298),
.A2(n_1259),
.B1(n_1294),
.B2(n_1313),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1313),
.A2(n_1198),
.B1(n_1232),
.B2(n_1215),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1313),
.A2(n_1196),
.B1(n_1251),
.B2(n_1246),
.Y(n_1374)
);

CKINVDCx11_ASAP7_75t_R g1375 ( 
.A(n_1239),
.Y(n_1375)
);

NAND2x1p5_ASAP7_75t_L g1376 ( 
.A(n_1265),
.B(n_1214),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1221),
.B(n_1211),
.Y(n_1377)
);

INVx6_ASAP7_75t_L g1378 ( 
.A(n_1305),
.Y(n_1378)
);

BUFx2_ASAP7_75t_L g1379 ( 
.A(n_1269),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1242),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1243),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1244),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_1255),
.Y(n_1383)
);

INVx4_ASAP7_75t_L g1384 ( 
.A(n_1231),
.Y(n_1384)
);

INVx3_ASAP7_75t_L g1385 ( 
.A(n_1248),
.Y(n_1385)
);

BUFx2_ASAP7_75t_L g1386 ( 
.A(n_1205),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1249),
.Y(n_1387)
);

INVx4_ASAP7_75t_L g1388 ( 
.A(n_1308),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1233),
.A2(n_1256),
.B1(n_1240),
.B2(n_1225),
.Y(n_1389)
);

NAND2x1p5_ASAP7_75t_L g1390 ( 
.A(n_1277),
.B(n_1305),
.Y(n_1390)
);

AOI21xp33_ASAP7_75t_L g1391 ( 
.A1(n_1264),
.A2(n_1202),
.B(n_1262),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1290),
.Y(n_1392)
);

CKINVDCx20_ASAP7_75t_R g1393 ( 
.A(n_1263),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1312),
.Y(n_1394)
);

NAND2x1p5_ASAP7_75t_L g1395 ( 
.A(n_1212),
.B(n_1253),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_SL g1396 ( 
.A1(n_1279),
.A2(n_1295),
.B1(n_1328),
.B2(n_1216),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1219),
.A2(n_1212),
.B1(n_1272),
.B2(n_1218),
.Y(n_1397)
);

OAI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1235),
.A2(n_1339),
.B1(n_1328),
.B2(n_1295),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1271),
.B(n_1268),
.Y(n_1399)
);

OAI21xp5_ASAP7_75t_SL g1400 ( 
.A1(n_1204),
.A2(n_1328),
.B(n_1295),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1216),
.A2(n_1261),
.B1(n_1327),
.B2(n_1315),
.Y(n_1401)
);

INVx3_ASAP7_75t_L g1402 ( 
.A(n_1253),
.Y(n_1402)
);

BUFx12f_ASAP7_75t_L g1403 ( 
.A(n_1287),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1276),
.A2(n_1270),
.B1(n_1286),
.B2(n_1273),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1286),
.A2(n_1204),
.B1(n_1267),
.B2(n_1191),
.Y(n_1405)
);

BUFx12f_ASAP7_75t_L g1406 ( 
.A(n_1281),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1204),
.A2(n_1267),
.B1(n_1191),
.B2(n_1228),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1288),
.Y(n_1408)
);

CKINVDCx11_ASAP7_75t_R g1409 ( 
.A(n_1281),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1250),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1230),
.Y(n_1411)
);

BUFx2_ASAP7_75t_SL g1412 ( 
.A(n_1260),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1281),
.A2(n_1222),
.B1(n_1260),
.B2(n_1195),
.Y(n_1413)
);

INVx4_ASAP7_75t_L g1414 ( 
.A(n_1282),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1300),
.A2(n_1241),
.B1(n_1254),
.B2(n_1194),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1274),
.Y(n_1416)
);

INVx3_ASAP7_75t_L g1417 ( 
.A(n_1250),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_SL g1418 ( 
.A1(n_1236),
.A2(n_1258),
.B(n_1209),
.Y(n_1418)
);

BUFx2_ASAP7_75t_SL g1419 ( 
.A(n_1282),
.Y(n_1419)
);

BUFx10_ASAP7_75t_L g1420 ( 
.A(n_1280),
.Y(n_1420)
);

BUFx10_ASAP7_75t_L g1421 ( 
.A(n_1275),
.Y(n_1421)
);

BUFx4f_ASAP7_75t_SL g1422 ( 
.A(n_1257),
.Y(n_1422)
);

OAI21xp33_ASAP7_75t_L g1423 ( 
.A1(n_1254),
.A2(n_1199),
.B(n_1206),
.Y(n_1423)
);

BUFx2_ASAP7_75t_SL g1424 ( 
.A(n_1300),
.Y(n_1424)
);

BUFx2_ASAP7_75t_SL g1425 ( 
.A(n_1237),
.Y(n_1425)
);

INVx6_ASAP7_75t_L g1426 ( 
.A(n_1284),
.Y(n_1426)
);

OAI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1297),
.A2(n_1331),
.B1(n_1343),
.B2(n_1314),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1199),
.A2(n_1220),
.B1(n_1208),
.B2(n_1229),
.Y(n_1428)
);

INVx6_ASAP7_75t_L g1429 ( 
.A(n_1318),
.Y(n_1429)
);

INVx1_ASAP7_75t_SL g1430 ( 
.A(n_1283),
.Y(n_1430)
);

BUFx10_ASAP7_75t_L g1431 ( 
.A(n_1342),
.Y(n_1431)
);

CKINVDCx11_ASAP7_75t_R g1432 ( 
.A(n_1257),
.Y(n_1432)
);

BUFx10_ASAP7_75t_L g1433 ( 
.A(n_1257),
.Y(n_1433)
);

INVx4_ASAP7_75t_L g1434 ( 
.A(n_1210),
.Y(n_1434)
);

INVx4_ASAP7_75t_L g1435 ( 
.A(n_1245),
.Y(n_1435)
);

OAI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1309),
.A2(n_1346),
.B1(n_1330),
.B2(n_1332),
.Y(n_1436)
);

OAI21xp5_ASAP7_75t_SL g1437 ( 
.A1(n_1321),
.A2(n_1333),
.B(n_1337),
.Y(n_1437)
);

BUFx3_ASAP7_75t_L g1438 ( 
.A(n_1189),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1301),
.Y(n_1439)
);

INVx5_ASAP7_75t_L g1440 ( 
.A(n_1190),
.Y(n_1440)
);

CKINVDCx11_ASAP7_75t_R g1441 ( 
.A(n_1220),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1319),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1319),
.Y(n_1443)
);

BUFx8_ASAP7_75t_L g1444 ( 
.A(n_1220),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1319),
.Y(n_1445)
);

BUFx10_ASAP7_75t_L g1446 ( 
.A(n_1324),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1278),
.Y(n_1447)
);

OAI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1192),
.A2(n_1197),
.B1(n_1324),
.B2(n_1340),
.Y(n_1448)
);

CKINVDCx20_ASAP7_75t_R g1449 ( 
.A(n_1278),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1324),
.A2(n_1340),
.B1(n_1289),
.B2(n_1296),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1188),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1307),
.Y(n_1452)
);

INVx6_ASAP7_75t_L g1453 ( 
.A(n_1193),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_SL g1454 ( 
.A1(n_1304),
.A2(n_1341),
.B1(n_1317),
.B2(n_989),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1302),
.A2(n_1341),
.B1(n_1317),
.B2(n_1320),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1317),
.A2(n_1341),
.B1(n_1291),
.B2(n_1325),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1227),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1291),
.A2(n_1302),
.B1(n_1345),
.B2(n_1306),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1217),
.Y(n_1459)
);

OAI21xp33_ASAP7_75t_L g1460 ( 
.A1(n_1291),
.A2(n_1344),
.B(n_1302),
.Y(n_1460)
);

INVx4_ASAP7_75t_L g1461 ( 
.A(n_1266),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1302),
.A2(n_1341),
.B1(n_1317),
.B2(n_1320),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_SL g1463 ( 
.A1(n_1317),
.A2(n_1341),
.B1(n_989),
.B2(n_807),
.Y(n_1463)
);

CKINVDCx11_ASAP7_75t_R g1464 ( 
.A(n_1207),
.Y(n_1464)
);

CKINVDCx20_ASAP7_75t_R g1465 ( 
.A(n_1224),
.Y(n_1465)
);

INVx1_ASAP7_75t_SL g1466 ( 
.A(n_1203),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1217),
.Y(n_1467)
);

OAI21xp5_ASAP7_75t_SL g1468 ( 
.A1(n_1291),
.A2(n_1302),
.B(n_1317),
.Y(n_1468)
);

CKINVDCx20_ASAP7_75t_R g1469 ( 
.A(n_1224),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1302),
.A2(n_1341),
.B1(n_1317),
.B2(n_1320),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1302),
.A2(n_1341),
.B1(n_1317),
.B2(n_1320),
.Y(n_1471)
);

NAND2x1p5_ASAP7_75t_L g1472 ( 
.A(n_1298),
.B(n_1265),
.Y(n_1472)
);

AND2x4_ASAP7_75t_SL g1473 ( 
.A(n_1224),
.B(n_854),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1302),
.A2(n_1341),
.B1(n_1317),
.B2(n_1320),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_SL g1475 ( 
.A1(n_1317),
.A2(n_1341),
.B1(n_989),
.B2(n_807),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1217),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1311),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1317),
.A2(n_1341),
.B1(n_989),
.B2(n_807),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1227),
.Y(n_1479)
);

BUFx2_ASAP7_75t_L g1480 ( 
.A(n_1203),
.Y(n_1480)
);

OR2x6_ASAP7_75t_L g1481 ( 
.A(n_1400),
.B(n_1447),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1450),
.A2(n_1415),
.B(n_1397),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1410),
.Y(n_1483)
);

INVx3_ASAP7_75t_L g1484 ( 
.A(n_1438),
.Y(n_1484)
);

AOI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1389),
.A2(n_1452),
.B(n_1365),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1468),
.B(n_1360),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1415),
.A2(n_1451),
.B(n_1411),
.Y(n_1487)
);

BUFx3_ASAP7_75t_L g1488 ( 
.A(n_1409),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1348),
.A2(n_1456),
.B1(n_1470),
.B2(n_1471),
.Y(n_1489)
);

BUFx3_ASAP7_75t_L g1490 ( 
.A(n_1406),
.Y(n_1490)
);

AO21x2_ASAP7_75t_L g1491 ( 
.A1(n_1448),
.A2(n_1398),
.B(n_1439),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1379),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1442),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1440),
.B(n_1405),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1443),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1445),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1463),
.A2(n_1478),
.B1(n_1475),
.B2(n_1441),
.Y(n_1497)
);

OAI211xp5_ASAP7_75t_L g1498 ( 
.A1(n_1460),
.A2(n_1351),
.B(n_1474),
.C(n_1462),
.Y(n_1498)
);

AOI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1427),
.A2(n_1436),
.B(n_1437),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1463),
.A2(n_1475),
.B1(n_1478),
.B2(n_1357),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1353),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1440),
.B(n_1405),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1359),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1377),
.Y(n_1504)
);

INVx1_ASAP7_75t_SL g1505 ( 
.A(n_1393),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1413),
.A2(n_1418),
.B(n_1417),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1416),
.Y(n_1507)
);

BUFx2_ASAP7_75t_SL g1508 ( 
.A(n_1355),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1354),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1368),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1380),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1417),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1381),
.Y(n_1513)
);

BUFx2_ASAP7_75t_L g1514 ( 
.A(n_1422),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1455),
.A2(n_1474),
.B1(n_1462),
.B2(n_1471),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_SL g1516 ( 
.A(n_1349),
.B(n_1465),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1440),
.B(n_1382),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1387),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1354),
.Y(n_1519)
);

BUFx4f_ASAP7_75t_SL g1520 ( 
.A(n_1469),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1408),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_SL g1522 ( 
.A1(n_1444),
.A2(n_1422),
.B1(n_1458),
.B2(n_1449),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_1408),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1455),
.A2(n_1470),
.B1(n_1357),
.B2(n_1367),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1392),
.Y(n_1525)
);

OAI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1370),
.A2(n_1367),
.B(n_1364),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1394),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1459),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1467),
.Y(n_1529)
);

INVx2_ASAP7_75t_SL g1530 ( 
.A(n_1420),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1476),
.Y(n_1531)
);

OA21x2_ASAP7_75t_L g1532 ( 
.A1(n_1423),
.A2(n_1407),
.B(n_1391),
.Y(n_1532)
);

OAI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1454),
.A2(n_1427),
.B(n_1436),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1446),
.Y(n_1534)
);

OAI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1413),
.A2(n_1407),
.B(n_1404),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1424),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1433),
.B(n_1396),
.Y(n_1537)
);

CKINVDCx8_ASAP7_75t_R g1538 ( 
.A(n_1412),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1433),
.B(n_1396),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1430),
.Y(n_1540)
);

NOR2x1_ASAP7_75t_L g1541 ( 
.A(n_1434),
.B(n_1435),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1398),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_SL g1543 ( 
.A1(n_1444),
.A2(n_1432),
.B1(n_1426),
.B2(n_1429),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1453),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1401),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1401),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_1358),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1366),
.B(n_1454),
.Y(n_1548)
);

AO21x2_ASAP7_75t_L g1549 ( 
.A1(n_1448),
.A2(n_1399),
.B(n_1477),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1428),
.B(n_1374),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1428),
.B(n_1374),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1420),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1373),
.B(n_1434),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1435),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1453),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1425),
.Y(n_1556)
);

AOI21xp33_ASAP7_75t_L g1557 ( 
.A1(n_1404),
.A2(n_1372),
.B(n_1371),
.Y(n_1557)
);

OAI221xp5_ASAP7_75t_L g1558 ( 
.A1(n_1373),
.A2(n_1371),
.B1(n_1363),
.B2(n_1372),
.C(n_1429),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1426),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1464),
.Y(n_1560)
);

BUFx4_ASAP7_75t_R g1561 ( 
.A(n_1369),
.Y(n_1561)
);

BUFx4f_ASAP7_75t_SL g1562 ( 
.A(n_1356),
.Y(n_1562)
);

INVx3_ASAP7_75t_SL g1563 ( 
.A(n_1426),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1429),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1386),
.B(n_1480),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1431),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1385),
.B(n_1479),
.Y(n_1567)
);

CKINVDCx10_ASAP7_75t_R g1568 ( 
.A(n_1350),
.Y(n_1568)
);

OAI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1376),
.A2(n_1363),
.B(n_1466),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1431),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1421),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1352),
.B(n_1457),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1421),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1390),
.B(n_1385),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1419),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1414),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1402),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1402),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1395),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1486),
.B(n_1361),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1504),
.B(n_1361),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_1568),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1492),
.B(n_1461),
.Y(n_1583)
);

AOI21x1_ASAP7_75t_L g1584 ( 
.A1(n_1566),
.A2(n_1570),
.B(n_1540),
.Y(n_1584)
);

OAI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1489),
.A2(n_1376),
.B(n_1472),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1507),
.B(n_1461),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1513),
.Y(n_1587)
);

O2A1O1Ixp33_ASAP7_75t_L g1588 ( 
.A1(n_1515),
.A2(n_1383),
.B(n_1472),
.C(n_1390),
.Y(n_1588)
);

AOI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1524),
.A2(n_1362),
.B1(n_1378),
.B2(n_1375),
.Y(n_1589)
);

BUFx2_ASAP7_75t_L g1590 ( 
.A(n_1492),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1498),
.A2(n_1384),
.B1(n_1388),
.B2(n_1362),
.Y(n_1591)
);

O2A1O1Ixp33_ASAP7_75t_L g1592 ( 
.A1(n_1526),
.A2(n_1395),
.B(n_1403),
.C(n_1362),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1537),
.B(n_1384),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1537),
.B(n_1369),
.Y(n_1594)
);

BUFx6f_ASAP7_75t_L g1595 ( 
.A(n_1563),
.Y(n_1595)
);

O2A1O1Ixp5_ASAP7_75t_L g1596 ( 
.A1(n_1533),
.A2(n_1378),
.B(n_1473),
.C(n_1499),
.Y(n_1596)
);

AOI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1500),
.A2(n_1497),
.B1(n_1522),
.B2(n_1558),
.Y(n_1597)
);

INVx4_ASAP7_75t_L g1598 ( 
.A(n_1563),
.Y(n_1598)
);

OAI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1543),
.A2(n_1563),
.B1(n_1566),
.B2(n_1570),
.Y(n_1599)
);

BUFx6f_ASAP7_75t_SL g1600 ( 
.A(n_1488),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1539),
.B(n_1517),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1568),
.Y(n_1602)
);

O2A1O1Ixp33_ASAP7_75t_L g1603 ( 
.A1(n_1569),
.A2(n_1542),
.B(n_1550),
.C(n_1551),
.Y(n_1603)
);

AOI22xp5_ASAP7_75t_SL g1604 ( 
.A1(n_1488),
.A2(n_1560),
.B1(n_1547),
.B2(n_1548),
.Y(n_1604)
);

OAI22xp5_ASAP7_75t_SL g1605 ( 
.A1(n_1488),
.A2(n_1508),
.B1(n_1520),
.B2(n_1562),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1538),
.A2(n_1564),
.B1(n_1565),
.B2(n_1550),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1567),
.B(n_1514),
.Y(n_1607)
);

NAND4xp25_ASAP7_75t_L g1608 ( 
.A(n_1565),
.B(n_1552),
.C(n_1575),
.D(n_1572),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1567),
.B(n_1514),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1538),
.A2(n_1564),
.B1(n_1551),
.B2(n_1553),
.Y(n_1610)
);

OAI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1485),
.A2(n_1540),
.B(n_1482),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1548),
.B(n_1501),
.Y(n_1612)
);

AOI221xp5_ASAP7_75t_L g1613 ( 
.A1(n_1542),
.A2(n_1491),
.B1(n_1557),
.B2(n_1531),
.C(n_1529),
.Y(n_1613)
);

AOI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1491),
.A2(n_1528),
.B1(n_1531),
.B2(n_1510),
.C(n_1529),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1553),
.A2(n_1559),
.B1(n_1481),
.B2(n_1505),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1494),
.B(n_1502),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1503),
.B(n_1510),
.Y(n_1617)
);

INVx3_ASAP7_75t_L g1618 ( 
.A(n_1484),
.Y(n_1618)
);

OA21x2_ASAP7_75t_L g1619 ( 
.A1(n_1482),
.A2(n_1506),
.B(n_1535),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1511),
.B(n_1518),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1511),
.B(n_1518),
.Y(n_1621)
);

INVx3_ASAP7_75t_L g1622 ( 
.A(n_1484),
.Y(n_1622)
);

OAI21x1_ASAP7_75t_SL g1623 ( 
.A1(n_1530),
.A2(n_1559),
.B(n_1575),
.Y(n_1623)
);

OA21x2_ASAP7_75t_L g1624 ( 
.A1(n_1506),
.A2(n_1535),
.B(n_1487),
.Y(n_1624)
);

BUFx6f_ASAP7_75t_SL g1625 ( 
.A(n_1490),
.Y(n_1625)
);

OAI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1485),
.A2(n_1556),
.B(n_1541),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1525),
.B(n_1527),
.Y(n_1627)
);

AOI221xp5_ASAP7_75t_L g1628 ( 
.A1(n_1491),
.A2(n_1528),
.B1(n_1527),
.B2(n_1545),
.C(n_1546),
.Y(n_1628)
);

AO32x2_ASAP7_75t_L g1629 ( 
.A1(n_1530),
.A2(n_1549),
.A3(n_1523),
.B1(n_1481),
.B2(n_1532),
.Y(n_1629)
);

AOI221x1_ASAP7_75t_SL g1630 ( 
.A1(n_1552),
.A2(n_1571),
.B1(n_1573),
.B2(n_1577),
.C(n_1578),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1571),
.B(n_1573),
.Y(n_1631)
);

OA21x2_ASAP7_75t_L g1632 ( 
.A1(n_1487),
.A2(n_1536),
.B(n_1545),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1577),
.B(n_1578),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1574),
.B(n_1523),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1579),
.B(n_1519),
.Y(n_1635)
);

AO32x2_ASAP7_75t_L g1636 ( 
.A1(n_1549),
.A2(n_1532),
.A3(n_1519),
.B1(n_1521),
.B2(n_1509),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1509),
.B(n_1521),
.Y(n_1637)
);

NAND4xp25_ASAP7_75t_L g1638 ( 
.A(n_1516),
.B(n_1541),
.C(n_1554),
.D(n_1536),
.Y(n_1638)
);

AO32x1_ASAP7_75t_L g1639 ( 
.A1(n_1509),
.A2(n_1521),
.A3(n_1519),
.B1(n_1554),
.B2(n_1512),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1532),
.B(n_1544),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1614),
.B(n_1532),
.Y(n_1641)
);

NAND4xp25_ASAP7_75t_L g1642 ( 
.A(n_1630),
.B(n_1561),
.C(n_1579),
.D(n_1490),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_SL g1643 ( 
.A(n_1595),
.B(n_1576),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1597),
.A2(n_1613),
.B1(n_1628),
.B2(n_1585),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1610),
.A2(n_1549),
.B1(n_1594),
.B2(n_1606),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1619),
.B(n_1555),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1621),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1621),
.Y(n_1648)
);

INVx3_ASAP7_75t_L g1649 ( 
.A(n_1618),
.Y(n_1649)
);

INVxp67_ASAP7_75t_L g1650 ( 
.A(n_1590),
.Y(n_1650)
);

INVx3_ASAP7_75t_L g1651 ( 
.A(n_1618),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1637),
.B(n_1483),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1619),
.B(n_1512),
.Y(n_1653)
);

NOR2x1p5_ASAP7_75t_L g1654 ( 
.A(n_1638),
.B(n_1490),
.Y(n_1654)
);

BUFx3_ASAP7_75t_L g1655 ( 
.A(n_1595),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1616),
.B(n_1496),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1627),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1627),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1617),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1616),
.B(n_1640),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1632),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1620),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1632),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1587),
.B(n_1495),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1612),
.B(n_1634),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1636),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1632),
.Y(n_1667)
);

NOR2xp67_ASAP7_75t_L g1668 ( 
.A(n_1640),
.B(n_1534),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1635),
.B(n_1496),
.Y(n_1669)
);

INVx3_ASAP7_75t_L g1670 ( 
.A(n_1622),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1636),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1633),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1601),
.B(n_1493),
.Y(n_1673)
);

INVx4_ASAP7_75t_L g1674 ( 
.A(n_1598),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_1582),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1660),
.B(n_1629),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1660),
.B(n_1629),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1660),
.B(n_1593),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1653),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1661),
.Y(n_1680)
);

OR2x2_ASAP7_75t_SL g1681 ( 
.A(n_1641),
.B(n_1581),
.Y(n_1681)
);

NAND2x1_ASAP7_75t_L g1682 ( 
.A(n_1649),
.B(n_1623),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1647),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1653),
.Y(n_1684)
);

OAI221xp5_ASAP7_75t_L g1685 ( 
.A1(n_1644),
.A2(n_1603),
.B1(n_1596),
.B2(n_1589),
.C(n_1588),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1656),
.B(n_1673),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1641),
.A2(n_1639),
.B(n_1611),
.Y(n_1687)
);

OAI33xp33_ASAP7_75t_L g1688 ( 
.A1(n_1664),
.A2(n_1631),
.A3(n_1608),
.B1(n_1599),
.B2(n_1591),
.B3(n_1615),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1647),
.Y(n_1689)
);

INVxp67_ASAP7_75t_SL g1690 ( 
.A(n_1661),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1647),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1663),
.Y(n_1692)
);

INVx3_ASAP7_75t_L g1693 ( 
.A(n_1649),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1669),
.B(n_1584),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1673),
.B(n_1593),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1656),
.B(n_1629),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1673),
.B(n_1607),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_SL g1698 ( 
.A1(n_1644),
.A2(n_1605),
.B1(n_1580),
.B2(n_1602),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1656),
.B(n_1609),
.Y(n_1699)
);

NAND2x1p5_ASAP7_75t_L g1700 ( 
.A(n_1674),
.B(n_1598),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1669),
.B(n_1626),
.Y(n_1701)
);

BUFx3_ASAP7_75t_L g1702 ( 
.A(n_1655),
.Y(n_1702)
);

NAND2x1_ASAP7_75t_L g1703 ( 
.A(n_1651),
.B(n_1594),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1648),
.B(n_1629),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1664),
.B(n_1601),
.Y(n_1705)
);

OR2x2_ASAP7_75t_SL g1706 ( 
.A(n_1666),
.B(n_1586),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1653),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1701),
.B(n_1665),
.Y(n_1708)
);

AOI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1685),
.A2(n_1645),
.B1(n_1580),
.B2(n_1654),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1701),
.B(n_1659),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_1693),
.B(n_1668),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1676),
.B(n_1648),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1683),
.Y(n_1713)
);

INVx1_ASAP7_75t_SL g1714 ( 
.A(n_1694),
.Y(n_1714)
);

INVx3_ASAP7_75t_L g1715 ( 
.A(n_1682),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1683),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1681),
.B(n_1665),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1693),
.B(n_1651),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1693),
.B(n_1651),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1680),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1693),
.B(n_1651),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1679),
.B(n_1651),
.Y(n_1722)
);

NOR2x1_ASAP7_75t_L g1723 ( 
.A(n_1682),
.B(n_1642),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1679),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1676),
.B(n_1657),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1689),
.Y(n_1726)
);

INVx2_ASAP7_75t_SL g1727 ( 
.A(n_1703),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1676),
.B(n_1657),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1677),
.B(n_1658),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1677),
.B(n_1696),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1681),
.B(n_1652),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1689),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1694),
.B(n_1659),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1677),
.B(n_1658),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1696),
.B(n_1686),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1679),
.B(n_1670),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1684),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1687),
.B(n_1662),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1696),
.B(n_1650),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1686),
.B(n_1650),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1686),
.B(n_1672),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1684),
.Y(n_1742)
);

HB1xp67_ASAP7_75t_L g1743 ( 
.A(n_1680),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1678),
.B(n_1672),
.Y(n_1744)
);

BUFx2_ASAP7_75t_L g1745 ( 
.A(n_1723),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1708),
.B(n_1687),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1708),
.B(n_1705),
.Y(n_1747)
);

INVx3_ASAP7_75t_L g1748 ( 
.A(n_1715),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1713),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1713),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1708),
.B(n_1705),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1713),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1723),
.B(n_1654),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1717),
.B(n_1738),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1723),
.B(n_1678),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1716),
.Y(n_1756)
);

INVxp33_ASAP7_75t_L g1757 ( 
.A(n_1717),
.Y(n_1757)
);

OAI22x1_ASAP7_75t_L g1758 ( 
.A1(n_1709),
.A2(n_1690),
.B1(n_1692),
.B2(n_1688),
.Y(n_1758)
);

OAI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1709),
.A2(n_1698),
.B1(n_1645),
.B2(n_1685),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1717),
.B(n_1704),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1716),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1738),
.B(n_1706),
.Y(n_1762)
);

AND2x4_ASAP7_75t_L g1763 ( 
.A(n_1735),
.B(n_1702),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1716),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1710),
.B(n_1706),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1730),
.B(n_1695),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1730),
.B(n_1695),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1714),
.B(n_1704),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1730),
.B(n_1702),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1735),
.B(n_1702),
.Y(n_1770)
);

NOR2x1_ASAP7_75t_L g1771 ( 
.A(n_1715),
.B(n_1642),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1724),
.Y(n_1772)
);

INVx2_ASAP7_75t_SL g1773 ( 
.A(n_1715),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1724),
.Y(n_1774)
);

NOR2x1p5_ASAP7_75t_SL g1775 ( 
.A(n_1724),
.B(n_1667),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1726),
.Y(n_1776)
);

AOI211xp5_ASAP7_75t_SL g1777 ( 
.A1(n_1715),
.A2(n_1698),
.B(n_1690),
.C(n_1692),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1724),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1710),
.B(n_1691),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1731),
.B(n_1691),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1731),
.B(n_1733),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1714),
.B(n_1704),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1735),
.B(n_1697),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1740),
.B(n_1697),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1740),
.B(n_1699),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1726),
.Y(n_1786)
);

INVx2_ASAP7_75t_SL g1787 ( 
.A(n_1715),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1753),
.B(n_1739),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1749),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1754),
.B(n_1731),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1754),
.B(n_1733),
.Y(n_1791)
);

AO211x2_ASAP7_75t_L g1792 ( 
.A1(n_1758),
.A2(n_1688),
.B(n_1667),
.C(n_1604),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1747),
.B(n_1739),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1747),
.B(n_1739),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1769),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1769),
.Y(n_1796)
);

AND2x4_ASAP7_75t_L g1797 ( 
.A(n_1753),
.B(n_1727),
.Y(n_1797)
);

CKINVDCx5p33_ASAP7_75t_R g1798 ( 
.A(n_1745),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1746),
.B(n_1720),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1749),
.Y(n_1800)
);

INVx2_ASAP7_75t_SL g1801 ( 
.A(n_1753),
.Y(n_1801)
);

INVx3_ASAP7_75t_SL g1802 ( 
.A(n_1763),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1771),
.B(n_1740),
.Y(n_1803)
);

NOR2x1_ASAP7_75t_L g1804 ( 
.A(n_1745),
.B(n_1711),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1758),
.B(n_1744),
.Y(n_1805)
);

AOI211x1_ASAP7_75t_SL g1806 ( 
.A1(n_1759),
.A2(n_1737),
.B(n_1742),
.C(n_1707),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1757),
.B(n_1744),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1784),
.B(n_1785),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1784),
.B(n_1785),
.Y(n_1809)
);

AND2x4_ASAP7_75t_L g1810 ( 
.A(n_1766),
.B(n_1727),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1771),
.B(n_1727),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1770),
.Y(n_1812)
);

OR2x2_ASAP7_75t_L g1813 ( 
.A(n_1751),
.B(n_1720),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1760),
.B(n_1781),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1781),
.B(n_1743),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1766),
.B(n_1744),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1767),
.B(n_1712),
.Y(n_1817)
);

INVx1_ASAP7_75t_SL g1818 ( 
.A(n_1755),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1750),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1767),
.B(n_1712),
.Y(n_1820)
);

INVx1_ASAP7_75t_SL g1821 ( 
.A(n_1755),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1780),
.B(n_1743),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1762),
.B(n_1741),
.Y(n_1823)
);

OR2x2_ASAP7_75t_L g1824 ( 
.A(n_1780),
.B(n_1726),
.Y(n_1824)
);

OAI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1803),
.A2(n_1777),
.B(n_1762),
.Y(n_1825)
);

AOI221xp5_ASAP7_75t_L g1826 ( 
.A1(n_1805),
.A2(n_1765),
.B1(n_1782),
.B2(n_1768),
.C(n_1671),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1789),
.Y(n_1827)
);

OAI221xp5_ASAP7_75t_L g1828 ( 
.A1(n_1806),
.A2(n_1765),
.B1(n_1666),
.B2(n_1671),
.C(n_1663),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1798),
.B(n_1783),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1800),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1798),
.B(n_1783),
.Y(n_1831)
);

AOI211xp5_ASAP7_75t_L g1832 ( 
.A1(n_1803),
.A2(n_1770),
.B(n_1763),
.C(n_1750),
.Y(n_1832)
);

AOI31xp33_ASAP7_75t_L g1833 ( 
.A1(n_1801),
.A2(n_1582),
.A3(n_1602),
.B(n_1675),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1819),
.Y(n_1834)
);

AOI21xp5_ASAP7_75t_L g1835 ( 
.A1(n_1792),
.A2(n_1787),
.B(n_1773),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1822),
.Y(n_1836)
);

AOI21xp33_ASAP7_75t_L g1837 ( 
.A1(n_1792),
.A2(n_1756),
.B(n_1752),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1802),
.B(n_1763),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1818),
.B(n_1779),
.Y(n_1839)
);

OAI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1811),
.A2(n_1773),
.B(n_1787),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1808),
.B(n_1809),
.Y(n_1841)
);

AOI221xp5_ASAP7_75t_L g1842 ( 
.A1(n_1790),
.A2(n_1821),
.B1(n_1823),
.B2(n_1799),
.C(n_1791),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1795),
.B(n_1779),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1822),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1793),
.B(n_1752),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1802),
.B(n_1748),
.Y(n_1846)
);

OAI21xp33_ASAP7_75t_L g1847 ( 
.A1(n_1788),
.A2(n_1775),
.B(n_1756),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_SL g1848 ( 
.A(n_1811),
.B(n_1748),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1795),
.B(n_1712),
.Y(n_1849)
);

OAI32xp33_ASAP7_75t_L g1850 ( 
.A1(n_1799),
.A2(n_1748),
.A3(n_1761),
.B1(n_1776),
.B2(n_1786),
.Y(n_1850)
);

AOI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1826),
.A2(n_1801),
.B1(n_1788),
.B2(n_1807),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1838),
.B(n_1796),
.Y(n_1852)
);

INVx1_ASAP7_75t_SL g1853 ( 
.A(n_1838),
.Y(n_1853)
);

AOI21xp33_ASAP7_75t_L g1854 ( 
.A1(n_1837),
.A2(n_1814),
.B(n_1815),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1845),
.Y(n_1855)
);

AOI22xp5_ASAP7_75t_L g1856 ( 
.A1(n_1825),
.A2(n_1796),
.B1(n_1812),
.B2(n_1666),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1845),
.Y(n_1857)
);

AOI21xp33_ASAP7_75t_L g1858 ( 
.A1(n_1836),
.A2(n_1815),
.B(n_1824),
.Y(n_1858)
);

AOI221xp5_ASAP7_75t_L g1859 ( 
.A1(n_1828),
.A2(n_1671),
.B1(n_1666),
.B2(n_1813),
.C(n_1772),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1844),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1835),
.A2(n_1804),
.B(n_1812),
.Y(n_1861)
);

NAND2x1_ASAP7_75t_SL g1862 ( 
.A(n_1846),
.B(n_1797),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1842),
.B(n_1816),
.Y(n_1863)
);

AOI22xp33_ASAP7_75t_SL g1864 ( 
.A1(n_1850),
.A2(n_1797),
.B1(n_1794),
.B2(n_1813),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_SL g1865 ( 
.A(n_1833),
.B(n_1797),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1841),
.B(n_1816),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1843),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1827),
.Y(n_1868)
);

AOI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1847),
.A2(n_1671),
.B1(n_1810),
.B2(n_1778),
.Y(n_1869)
);

INVxp33_ASAP7_75t_L g1870 ( 
.A(n_1829),
.Y(n_1870)
);

OAI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1864),
.A2(n_1848),
.B(n_1832),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1866),
.Y(n_1872)
);

OAI22xp33_ASAP7_75t_L g1873 ( 
.A1(n_1856),
.A2(n_1849),
.B1(n_1839),
.B2(n_1831),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1863),
.B(n_1817),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1853),
.B(n_1820),
.Y(n_1875)
);

OAI22xp33_ASAP7_75t_L g1876 ( 
.A1(n_1869),
.A2(n_1824),
.B1(n_1840),
.B2(n_1772),
.Y(n_1876)
);

XOR2x2_ASAP7_75t_L g1877 ( 
.A(n_1862),
.B(n_1848),
.Y(n_1877)
);

XNOR2x2_ASAP7_75t_L g1878 ( 
.A(n_1861),
.B(n_1846),
.Y(n_1878)
);

NAND2xp33_ASAP7_75t_L g1879 ( 
.A(n_1870),
.B(n_1675),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1855),
.Y(n_1880)
);

OAI21xp33_ASAP7_75t_L g1881 ( 
.A1(n_1864),
.A2(n_1834),
.B(n_1830),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1857),
.Y(n_1882)
);

AOI211xp5_ASAP7_75t_SL g1883 ( 
.A1(n_1881),
.A2(n_1854),
.B(n_1879),
.C(n_1858),
.Y(n_1883)
);

AND4x1_ASAP7_75t_L g1884 ( 
.A(n_1871),
.B(n_1852),
.C(n_1867),
.D(n_1860),
.Y(n_1884)
);

A2O1A1Ixp33_ASAP7_75t_L g1885 ( 
.A1(n_1871),
.A2(n_1859),
.B(n_1851),
.C(n_1775),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1875),
.B(n_1820),
.Y(n_1886)
);

NAND4xp25_ASAP7_75t_L g1887 ( 
.A(n_1874),
.B(n_1865),
.C(n_1868),
.D(n_1810),
.Y(n_1887)
);

OAI21xp33_ASAP7_75t_SL g1888 ( 
.A1(n_1878),
.A2(n_1865),
.B(n_1761),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1872),
.B(n_1810),
.Y(n_1889)
);

AND2x2_ASAP7_75t_SL g1890 ( 
.A(n_1882),
.B(n_1711),
.Y(n_1890)
);

NAND3xp33_ASAP7_75t_L g1891 ( 
.A(n_1880),
.B(n_1778),
.C(n_1774),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1877),
.Y(n_1892)
);

AOI211xp5_ASAP7_75t_L g1893 ( 
.A1(n_1873),
.A2(n_1786),
.B(n_1776),
.C(n_1764),
.Y(n_1893)
);

AOI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1892),
.A2(n_1876),
.B1(n_1600),
.B2(n_1774),
.Y(n_1894)
);

O2A1O1Ixp33_ASAP7_75t_L g1895 ( 
.A1(n_1888),
.A2(n_1764),
.B(n_1742),
.C(n_1737),
.Y(n_1895)
);

AOI21xp33_ASAP7_75t_SL g1896 ( 
.A1(n_1889),
.A2(n_1711),
.B(n_1736),
.Y(n_1896)
);

AOI321xp33_ASAP7_75t_L g1897 ( 
.A1(n_1883),
.A2(n_1592),
.A3(n_1667),
.B1(n_1737),
.B2(n_1742),
.C(n_1646),
.Y(n_1897)
);

AOI22xp33_ASAP7_75t_L g1898 ( 
.A1(n_1891),
.A2(n_1742),
.B1(n_1737),
.B2(n_1624),
.Y(n_1898)
);

OAI21xp5_ASAP7_75t_SL g1899 ( 
.A1(n_1884),
.A2(n_1700),
.B(n_1711),
.Y(n_1899)
);

OAI211xp5_ASAP7_75t_L g1900 ( 
.A1(n_1899),
.A2(n_1893),
.B(n_1887),
.C(n_1885),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1895),
.Y(n_1901)
);

OAI211xp5_ASAP7_75t_L g1902 ( 
.A1(n_1897),
.A2(n_1894),
.B(n_1896),
.C(n_1886),
.Y(n_1902)
);

AOI222xp33_ASAP7_75t_L g1903 ( 
.A1(n_1898),
.A2(n_1890),
.B1(n_1600),
.B2(n_1625),
.C1(n_1734),
.C2(n_1725),
.Y(n_1903)
);

NOR2xp33_ASAP7_75t_L g1904 ( 
.A(n_1899),
.B(n_1600),
.Y(n_1904)
);

XOR2x2_ASAP7_75t_L g1905 ( 
.A(n_1894),
.B(n_1625),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1901),
.Y(n_1906)
);

HB1xp67_ASAP7_75t_L g1907 ( 
.A(n_1900),
.Y(n_1907)
);

NOR2xp33_ASAP7_75t_L g1908 ( 
.A(n_1902),
.B(n_1625),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1905),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1904),
.Y(n_1910)
);

AOI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1907),
.A2(n_1903),
.B(n_1732),
.Y(n_1911)
);

OAI31xp33_ASAP7_75t_L g1912 ( 
.A1(n_1907),
.A2(n_1711),
.A3(n_1729),
.B(n_1728),
.Y(n_1912)
);

NAND3xp33_ASAP7_75t_L g1913 ( 
.A(n_1906),
.B(n_1711),
.C(n_1732),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1913),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1914),
.Y(n_1915)
);

CKINVDCx20_ASAP7_75t_R g1916 ( 
.A(n_1915),
.Y(n_1916)
);

INVx3_ASAP7_75t_L g1917 ( 
.A(n_1915),
.Y(n_1917)
);

AOI22xp5_ASAP7_75t_L g1918 ( 
.A1(n_1916),
.A2(n_1908),
.B1(n_1910),
.B2(n_1909),
.Y(n_1918)
);

HB1xp67_ASAP7_75t_L g1919 ( 
.A(n_1917),
.Y(n_1919)
);

HB1xp67_ASAP7_75t_L g1920 ( 
.A(n_1919),
.Y(n_1920)
);

OAI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1918),
.A2(n_1911),
.B(n_1912),
.Y(n_1921)
);

AOI221xp5_ASAP7_75t_L g1922 ( 
.A1(n_1920),
.A2(n_1732),
.B1(n_1707),
.B2(n_1725),
.C(n_1734),
.Y(n_1922)
);

OAI21x1_ASAP7_75t_L g1923 ( 
.A1(n_1922),
.A2(n_1921),
.B(n_1725),
.Y(n_1923)
);

AOI21xp5_ASAP7_75t_L g1924 ( 
.A1(n_1923),
.A2(n_1729),
.B(n_1728),
.Y(n_1924)
);

OAI221xp5_ASAP7_75t_R g1925 ( 
.A1(n_1924),
.A2(n_1718),
.B1(n_1719),
.B2(n_1721),
.C(n_1722),
.Y(n_1925)
);

AOI211xp5_ASAP7_75t_L g1926 ( 
.A1(n_1925),
.A2(n_1583),
.B(n_1595),
.C(n_1643),
.Y(n_1926)
);


endmodule