module fake_jpeg_7739_n_115 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_115);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_115;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx10_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_30),
.Y(n_44)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_17),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_31),
.B(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_24),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_15),
.B1(n_24),
.B2(n_23),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_14),
.B1(n_20),
.B2(n_21),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_34),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_19),
.B(n_16),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_25),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_28),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_60),
.C(n_61),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_15),
.B1(n_29),
.B2(n_24),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_51),
.B1(n_53),
.B2(n_57),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_47),
.B(n_48),
.Y(n_66)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_39),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_50),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_15),
.B1(n_27),
.B2(n_21),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_54),
.B1(n_58),
.B2(n_1),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_32),
.B1(n_20),
.B2(n_14),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_16),
.B1(n_19),
.B2(n_22),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_25),
.B1(n_12),
.B2(n_13),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_12),
.B1(n_22),
.B2(n_13),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_13),
.B(n_26),
.Y(n_60)
);

AND2x6_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_0),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_1),
.Y(n_62)
);

AO21x1_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_2),
.B(n_3),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_1),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_62),
.C(n_46),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_67),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_34),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_34),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_72),
.A2(n_10),
.B1(n_11),
.B2(n_26),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_71),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_76),
.B(n_79),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_47),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_80),
.C(n_81),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_61),
.B1(n_53),
.B2(n_57),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_84),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_59),
.B1(n_55),
.B2(n_49),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_83),
.A2(n_75),
.B1(n_64),
.B2(n_74),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_9),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_85),
.B(n_86),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_66),
.B(n_75),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_81),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_83),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_91),
.B(n_64),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_80),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_94),
.A2(n_74),
.B1(n_78),
.B2(n_65),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_SL g101 ( 
.A1(n_95),
.A2(n_92),
.B(n_88),
.C(n_90),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_87),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_100),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_98),
.B1(n_94),
.B2(n_89),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_65),
.C(n_63),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_101),
.A2(n_103),
.B(n_100),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_95),
.Y(n_108)
);

NOR2xp67_ASAP7_75t_SL g103 ( 
.A(n_99),
.B(n_93),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_107),
.Y(n_110)
);

OAI21x1_ASAP7_75t_SL g109 ( 
.A1(n_106),
.A2(n_86),
.B(n_72),
.Y(n_109)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_108),
.B(n_63),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_109),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_110),
.B(n_111),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_11),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_33),
.Y(n_115)
);


endmodule