module fake_jpeg_25925_n_46 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_46);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_46;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_17;
wire n_29;
wire n_37;
wire n_43;
wire n_32;
wire n_15;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

HB1xp67_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_21),
.Y(n_27)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_30),
.Y(n_35)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_25),
.B(n_9),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_21),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_31),
.B1(n_23),
.B2(n_19),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_31),
.B(n_34),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_33),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_SL g38 ( 
.A(n_37),
.B(n_33),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_39),
.C(n_32),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_26),
.B1(n_18),
.B2(n_17),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_40),
.B(n_41),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_17),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_0),
.B(n_12),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_43),
.C(n_20),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_22),
.Y(n_46)
);


endmodule