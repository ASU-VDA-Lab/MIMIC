module real_jpeg_14344_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_38;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_0),
.B(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_0),
.B(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_1),
.B(n_13),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_1),
.B(n_15),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_1),
.B(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_1),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_1),
.B(n_3),
.Y(n_42)
);

OR2x2_ASAP7_75t_SL g8 ( 
.A(n_2),
.B(n_9),
.Y(n_8)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_2),
.B(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_3),
.B(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_3),
.B(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_4),
.Y(n_9)
);

AO21x1_ASAP7_75t_L g15 ( 
.A1(n_5),
.A2(n_16),
.B(n_18),
.Y(n_15)
);

AO21x1_ASAP7_75t_SL g32 ( 
.A1(n_5),
.A2(n_33),
.B(n_35),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g6 ( 
.A(n_7),
.B(n_27),
.Y(n_6)
);

OAI22xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_10),
.B1(n_19),
.B2(n_21),
.Y(n_7)
);

AND2x2_ASAP7_75t_SL g37 ( 
.A(n_9),
.B(n_38),
.Y(n_37)
);

OR2x2_ASAP7_75t_SL g43 ( 
.A(n_9),
.B(n_38),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_14),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_12),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_13),
.B(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_17),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

INVxp33_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_36),
.B1(n_39),
.B2(n_43),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_42),
.Y(n_39)
);


endmodule