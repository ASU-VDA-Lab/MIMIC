module fake_jpeg_962_n_358 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_358);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_358;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_0),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_2),
.B(n_4),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_46),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_10),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_47),
.B(n_68),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_18),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_48),
.B(n_52),
.Y(n_102)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_49),
.Y(n_143)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_31),
.Y(n_55)
);

NAND2xp33_ASAP7_75t_SL g140 ( 
.A(n_55),
.B(n_75),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_57),
.Y(n_126)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_31),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_58),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

AND2x4_ASAP7_75t_SL g66 ( 
.A(n_44),
.B(n_32),
.Y(n_66)
);

AND2x4_ASAP7_75t_SL g142 ( 
.A(n_66),
.B(n_41),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_67),
.B(n_81),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_18),
.B(n_11),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_16),
.B(n_11),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_71),
.B(n_89),
.Y(n_98)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

INVxp67_ASAP7_75t_SL g75 ( 
.A(n_26),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_84),
.Y(n_104)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_80),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_35),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_42),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_87),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_24),
.B(n_8),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_42),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_91),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_90),
.A2(n_27),
.B1(n_29),
.B2(n_33),
.Y(n_101)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_93),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_16),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_94),
.B(n_95),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_24),
.B(n_12),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_51),
.A2(n_43),
.B1(n_17),
.B2(n_29),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_110),
.A2(n_115),
.B1(n_116),
.B2(n_124),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_48),
.A2(n_25),
.B1(n_33),
.B2(n_30),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_57),
.A2(n_25),
.B1(n_43),
.B2(n_30),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_82),
.A2(n_17),
.B1(n_39),
.B2(n_22),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_66),
.A2(n_41),
.B1(n_22),
.B2(n_21),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_127),
.A2(n_131),
.B1(n_21),
.B2(n_2),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_83),
.A2(n_41),
.B1(n_22),
.B2(n_13),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_84),
.A2(n_41),
.B1(n_13),
.B2(n_14),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_56),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_75),
.A2(n_73),
.B1(n_85),
.B2(n_63),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_136),
.A2(n_0),
.B1(n_2),
.B2(n_5),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_91),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_55),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_145),
.B(n_147),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_111),
.A2(n_89),
.B1(n_62),
.B2(n_74),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_146),
.A2(n_180),
.B1(n_107),
.B2(n_104),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_98),
.B(n_59),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_102),
.B(n_119),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_148),
.B(n_159),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_140),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_149),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_78),
.C(n_61),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_178),
.Y(n_190)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_153),
.Y(n_192)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

INVx11_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_155),
.Y(n_199)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_156),
.Y(n_197)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_157),
.Y(n_214)
);

O2A1O1Ixp33_ASAP7_75t_SL g158 ( 
.A1(n_142),
.A2(n_127),
.B(n_110),
.C(n_66),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_158),
.A2(n_107),
.B(n_136),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_103),
.B(n_70),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_129),
.B(n_79),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_165),
.Y(n_186)
);

AND2x2_ASAP7_75t_SL g189 ( 
.A(n_161),
.B(n_138),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_130),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_172),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_76),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_163),
.Y(n_202)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_106),
.Y(n_164)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_76),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_166),
.B(n_167),
.Y(n_207)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_126),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_15),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_168),
.B(n_170),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_105),
.B(n_60),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_173),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_96),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_171),
.Y(n_200)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_125),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_141),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_104),
.B(n_14),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_177),
.Y(n_210)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_176),
.Y(n_212)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_41),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_121),
.B(n_13),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_97),
.A2(n_54),
.B1(n_90),
.B2(n_21),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_179),
.A2(n_182),
.B1(n_183),
.B2(n_116),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_109),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_181),
.A2(n_184),
.B1(n_109),
.B2(n_132),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_97),
.A2(n_0),
.B1(n_2),
.B2(n_5),
.Y(n_183)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_132),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_185),
.A2(n_193),
.B1(n_144),
.B2(n_158),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_187),
.A2(n_144),
.B1(n_149),
.B2(n_161),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_188),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_189),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_177),
.A2(n_101),
.B1(n_117),
.B2(n_123),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_151),
.A2(n_114),
.B1(n_123),
.B2(n_112),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_195),
.A2(n_203),
.B1(n_206),
.B2(n_209),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_146),
.A2(n_112),
.B1(n_114),
.B2(n_100),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_180),
.A2(n_100),
.B1(n_118),
.B2(n_139),
.Y(n_206)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_208),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_170),
.A2(n_117),
.B1(n_128),
.B2(n_5),
.Y(n_209)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_214),
.Y(n_216)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_202),
.Y(n_217)
);

INVxp33_ASAP7_75t_L g252 ( 
.A(n_217),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_147),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_221),
.Y(n_245)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_220),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_154),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_145),
.Y(n_221)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_214),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_230),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_192),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_224),
.Y(n_255)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_225),
.B(n_229),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_161),
.C(n_148),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_190),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_227),
.A2(n_228),
.B1(n_189),
.B2(n_185),
.Y(n_253)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_169),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_231),
.B(n_194),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_204),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_234),
.Y(n_238)
);

NOR2x1_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_158),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_232),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_195),
.A2(n_159),
.B1(n_182),
.B2(n_183),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_236),
.A2(n_193),
.B1(n_187),
.B2(n_205),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_205),
.B(n_172),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_237),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_222),
.A2(n_188),
.B(n_213),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_240),
.A2(n_242),
.B(n_251),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_226),
.C(n_231),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_189),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_248),
.A2(n_249),
.B1(n_227),
.B2(n_221),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_229),
.A2(n_211),
.B1(n_213),
.B2(n_200),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_234),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_250),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_222),
.A2(n_200),
.B(n_204),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_253),
.A2(n_254),
.B1(n_236),
.B2(n_232),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_228),
.A2(n_189),
.B1(n_203),
.B2(n_206),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_218),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_263),
.Y(n_284)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_256),
.Y(n_259)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_259),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_260),
.A2(n_262),
.B1(n_270),
.B2(n_248),
.Y(n_280)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_256),
.Y(n_261)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_261),
.Y(n_290)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_269),
.C(n_241),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_239),
.B(n_186),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_265),
.B(n_266),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_186),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_247),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_267),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_230),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_235),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_253),
.A2(n_248),
.B1(n_254),
.B2(n_251),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_246),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_272),
.Y(n_285)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_246),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_244),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_288),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_243),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_275),
.B(n_282),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_243),
.C(n_238),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_283),
.C(n_287),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_257),
.A2(n_249),
.B(n_240),
.Y(n_277)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_277),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_280),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_238),
.C(n_242),
.Y(n_283)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_263),
.B(n_242),
.C(n_245),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_210),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_259),
.A2(n_250),
.B1(n_239),
.B2(n_251),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_289),
.A2(n_273),
.B(n_204),
.Y(n_299)
);

BUFx5_ASAP7_75t_L g291 ( 
.A(n_285),
.Y(n_291)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_291),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_261),
.Y(n_292)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_292),
.Y(n_314)
);

NAND3xp33_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_210),
.C(n_245),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_298),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_270),
.C(n_257),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_297),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_260),
.C(n_271),
.Y(n_298)
);

AO21x1_ASAP7_75t_L g307 ( 
.A1(n_299),
.A2(n_301),
.B(n_289),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_272),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_300),
.B(n_290),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_278),
.A2(n_219),
.B(n_225),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_305),
.A2(n_310),
.B1(n_311),
.B2(n_313),
.Y(n_322)
);

AOI21x1_ASAP7_75t_L g320 ( 
.A1(n_307),
.A2(n_314),
.B(n_298),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_276),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_309),
.B(n_316),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_302),
.A2(n_287),
.B1(n_279),
.B2(n_283),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_296),
.A2(n_233),
.B1(n_282),
.B2(n_255),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_296),
.A2(n_255),
.B1(n_209),
.B2(n_215),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_294),
.A2(n_215),
.B1(n_233),
.B2(n_223),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_315),
.A2(n_301),
.B1(n_291),
.B2(n_224),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_216),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_308),
.A2(n_299),
.B(n_300),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_318),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_297),
.C(n_295),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_320),
.B(n_198),
.Y(n_335)
);

XOR2x2_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_295),
.Y(n_321)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_321),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_304),
.C(n_292),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_323),
.B(n_324),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_312),
.B(n_304),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_325),
.A2(n_307),
.B1(n_305),
.B2(n_224),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_196),
.C(n_150),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_157),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_311),
.B(n_196),
.C(n_207),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_327),
.B(n_199),
.C(n_207),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_329),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_330),
.B(n_333),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_322),
.A2(n_171),
.B1(n_181),
.B2(n_192),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_332),
.B(n_334),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_318),
.B(n_198),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_335),
.A2(n_327),
.B(n_321),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_339),
.B(n_340),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_328),
.B(n_319),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_156),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_341),
.B(n_343),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_331),
.B(n_164),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_342),
.B(n_336),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_345),
.A2(n_346),
.B1(n_184),
.B2(n_162),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_337),
.A2(n_338),
.B1(n_332),
.B2(n_341),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_337),
.A2(n_329),
.B(n_330),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_348),
.A2(n_166),
.B(n_155),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_347),
.A2(n_176),
.B1(n_175),
.B2(n_152),
.Y(n_349)
);

OR2x2_ASAP7_75t_L g353 ( 
.A(n_349),
.B(n_350),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_344),
.B(n_153),
.C(n_167),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_351),
.B(n_352),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_353),
.A2(n_350),
.B(n_128),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_355),
.A2(n_354),
.B(n_12),
.Y(n_356)
);

AOI21x1_ASAP7_75t_L g357 ( 
.A1(n_356),
.A2(n_15),
.B(n_6),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_357),
.B(n_6),
.Y(n_358)
);


endmodule