module fake_jpeg_31404_n_550 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_550);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_550;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_49),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_59),
.B(n_63),
.Y(n_129)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_60),
.Y(n_122)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_61),
.Y(n_153)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx11_ASAP7_75t_L g138 ( 
.A(n_62),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_21),
.B(n_36),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_66),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_21),
.A2(n_17),
.B1(n_9),
.B2(n_4),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_67),
.A2(n_36),
.B1(n_33),
.B2(n_51),
.Y(n_151)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_69),
.Y(n_161)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_70),
.B(n_73),
.Y(n_149)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_71),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_72),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_75),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_78),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_82),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_30),
.B(n_11),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_83),
.B(n_89),
.Y(n_154)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_84),
.Y(n_170)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_49),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_18),
.B(n_11),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_90),
.B(n_95),
.Y(n_176)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_30),
.B(n_11),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_94),
.B(n_55),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_21),
.B(n_9),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_101),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_104),
.Y(n_159)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_25),
.Y(n_105)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_25),
.Y(n_106)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_106),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

BUFx8_ASAP7_75t_L g160 ( 
.A(n_107),
.Y(n_160)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_108),
.Y(n_162)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_39),
.Y(n_109)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_109),
.Y(n_174)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_38),
.Y(n_110)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

INVx4_ASAP7_75t_SL g111 ( 
.A(n_39),
.Y(n_111)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_38),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

INVx4_ASAP7_75t_SL g115 ( 
.A(n_111),
.Y(n_115)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_115),
.Y(n_186)
);

HAxp5_ASAP7_75t_SL g141 ( 
.A(n_63),
.B(n_39),
.CON(n_141),
.SN(n_141)
);

HAxp5_ASAP7_75t_SL g214 ( 
.A(n_141),
.B(n_39),
.CON(n_214),
.SN(n_214)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_143),
.B(n_45),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_151),
.A2(n_23),
.B1(n_28),
.B2(n_50),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_83),
.A2(n_55),
.B1(n_54),
.B2(n_37),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_155),
.A2(n_164),
.B1(n_175),
.B2(n_26),
.Y(n_201)
);

AND2x2_ASAP7_75t_SL g157 ( 
.A(n_70),
.B(n_14),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_32),
.C(n_46),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_158),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_61),
.A2(n_51),
.B1(n_28),
.B2(n_33),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_65),
.A2(n_36),
.B1(n_52),
.B2(n_41),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_165),
.A2(n_52),
.B1(n_41),
.B2(n_0),
.Y(n_221)
);

INVx4_ASAP7_75t_SL g167 ( 
.A(n_107),
.Y(n_167)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_167),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_102),
.Y(n_171)
);

BUFx8_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_90),
.A2(n_54),
.B1(n_50),
.B2(n_37),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_97),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_178),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g179 ( 
.A(n_107),
.Y(n_179)
);

INVx11_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_123),
.Y(n_180)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_180),
.Y(n_241)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_181),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_115),
.A2(n_93),
.B1(n_112),
.B2(n_32),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_182),
.A2(n_202),
.B1(n_212),
.B2(n_124),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_120),
.B(n_95),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_183),
.B(n_193),
.Y(n_242)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_136),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_184),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_185),
.A2(n_210),
.B1(n_233),
.B2(n_178),
.Y(n_263)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_136),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_187),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_129),
.B(n_38),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_188),
.B(n_190),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_176),
.A2(n_80),
.B1(n_99),
.B2(n_91),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_189),
.A2(n_198),
.B1(n_207),
.B2(n_222),
.Y(n_277)
);

OA22x2_ASAP7_75t_L g190 ( 
.A1(n_141),
.A2(n_67),
.B1(n_62),
.B2(n_64),
.Y(n_190)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_191),
.Y(n_282)
);

BUFx16f_ASAP7_75t_L g192 ( 
.A(n_167),
.Y(n_192)
);

CKINVDCx6p67_ASAP7_75t_R g280 ( 
.A(n_192),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_130),
.B(n_45),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_195),
.B(n_217),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_196),
.B(n_201),
.Y(n_247)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_138),
.Y(n_197)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_197),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_148),
.A2(n_101),
.B1(n_79),
.B2(n_78),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_118),
.Y(n_199)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_199),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_149),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_205),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_121),
.A2(n_52),
.B1(n_41),
.B2(n_74),
.Y(n_202)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_162),
.Y(n_203)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_132),
.Y(n_204)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_204),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_149),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_174),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_206),
.B(n_216),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_176),
.A2(n_76),
.B1(n_72),
.B2(n_69),
.Y(n_207)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_208),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_164),
.A2(n_77),
.B1(n_46),
.B2(n_34),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_168),
.A2(n_52),
.B1(n_41),
.B2(n_34),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_122),
.Y(n_213)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_213),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_214),
.B(n_218),
.Y(n_253)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_163),
.Y(n_215)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_215),
.Y(n_281)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_135),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_154),
.B(n_26),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_129),
.B(n_52),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_177),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_219),
.B(n_220),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_140),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_221),
.A2(n_119),
.B1(n_147),
.B2(n_125),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_L g222 ( 
.A1(n_127),
.A2(n_41),
.B1(n_12),
.B2(n_5),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_154),
.B(n_9),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_223),
.B(n_225),
.Y(n_258)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_158),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_224),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_117),
.B(n_12),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_126),
.A2(n_137),
.B1(n_145),
.B2(n_114),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_226),
.A2(n_237),
.B1(n_166),
.B2(n_139),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_116),
.B(n_0),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_218),
.Y(n_260)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_152),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_229),
.B(n_230),
.Y(n_265)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_159),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_172),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_231),
.Y(n_252)
);

OA22x2_ASAP7_75t_L g233 ( 
.A1(n_165),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_160),
.B(n_12),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_234),
.B(n_160),
.Y(n_249)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_131),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_235),
.Y(n_268)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_153),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_236),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_134),
.A2(n_17),
.B1(n_5),
.B2(n_6),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_157),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_240),
.B(n_246),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_153),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_249),
.B(n_256),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_250),
.A2(n_270),
.B1(n_273),
.B2(n_279),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_205),
.B(n_173),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_251),
.B(n_254),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_201),
.B(n_188),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_255),
.A2(n_233),
.B1(n_232),
.B2(n_204),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_196),
.B(n_133),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_260),
.B(n_263),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_266),
.A2(n_199),
.B1(n_211),
.B2(n_192),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_190),
.A2(n_156),
.B1(n_144),
.B2(n_146),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_269),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_185),
.A2(n_173),
.B1(n_170),
.B2(n_169),
.Y(n_270)
);

NAND3xp33_ASAP7_75t_SL g271 ( 
.A(n_214),
.B(n_142),
.C(n_179),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_271),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_190),
.A2(n_150),
.B1(n_171),
.B2(n_179),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_190),
.A2(n_142),
.B1(n_6),
.B2(n_7),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_278),
.A2(n_277),
.B1(n_266),
.B2(n_254),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_237),
.A2(n_226),
.B1(n_207),
.B2(n_189),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_283),
.Y(n_337)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_284),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_279),
.A2(n_236),
.B1(n_208),
.B2(n_191),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_285),
.A2(n_268),
.B1(n_274),
.B2(n_252),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_286),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_238),
.B(n_218),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_288),
.A2(n_292),
.B(n_264),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_262),
.A2(n_197),
.B1(n_216),
.B2(n_219),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_290),
.A2(n_295),
.B1(n_244),
.B2(n_276),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_238),
.A2(n_233),
.B(n_188),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_265),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_294),
.B(n_301),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_262),
.A2(n_233),
.B1(n_186),
.B2(n_232),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_277),
.A2(n_181),
.B1(n_180),
.B2(n_235),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_238),
.A2(n_231),
.B1(n_222),
.B2(n_199),
.Y(n_298)
);

AND2x2_ASAP7_75t_SL g300 ( 
.A(n_246),
.B(n_184),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_300),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_280),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_267),
.Y(n_302)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_302),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_273),
.A2(n_253),
.B(n_263),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_303),
.A2(n_292),
.B(n_312),
.Y(n_326)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_281),
.Y(n_304)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_304),
.Y(n_331)
);

OAI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_270),
.A2(n_203),
.B1(n_224),
.B2(n_187),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_306),
.A2(n_272),
.B1(n_268),
.B2(n_252),
.Y(n_339)
);

BUFx5_ASAP7_75t_L g307 ( 
.A(n_280),
.Y(n_307)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_307),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_280),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_308),
.Y(n_323)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_259),
.Y(n_309)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_309),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_251),
.B(n_209),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_314),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_280),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_311),
.Y(n_348)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_281),
.Y(n_313)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_313),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_247),
.B(n_192),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_247),
.B(n_1),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_317),
.Y(n_320)
);

OAI32xp33_ASAP7_75t_L g316 ( 
.A1(n_250),
.A2(n_6),
.A3(n_7),
.B1(n_12),
.B2(n_14),
.Y(n_316)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_316),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_247),
.B(n_6),
.Y(n_317)
);

OAI32xp33_ASAP7_75t_L g318 ( 
.A1(n_305),
.A2(n_243),
.A3(n_256),
.B1(n_240),
.B2(n_242),
.Y(n_318)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_318),
.Y(n_353)
);

INVxp33_ASAP7_75t_L g322 ( 
.A(n_301),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g378 ( 
.A(n_322),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_326),
.A2(n_292),
.B(n_303),
.Y(n_352)
);

INVx13_ASAP7_75t_L g327 ( 
.A(n_307),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_327),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_329),
.A2(n_333),
.B1(n_346),
.B2(n_306),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_293),
.B(n_260),
.C(n_253),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_330),
.B(n_293),
.C(n_288),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_305),
.B(n_249),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_332),
.B(n_289),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_296),
.A2(n_253),
.B1(n_258),
.B2(n_257),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_287),
.B(n_248),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_334),
.B(n_294),
.Y(n_351)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_307),
.Y(n_335)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_335),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_336),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_339),
.A2(n_343),
.B1(n_295),
.B2(n_283),
.Y(n_350)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_304),
.Y(n_342)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_342),
.Y(n_358)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_313),
.Y(n_344)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_344),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_296),
.A2(n_274),
.B1(n_276),
.B2(n_282),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_330),
.B(n_293),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_349),
.B(n_320),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_350),
.A2(n_346),
.B1(n_343),
.B2(n_291),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_351),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_352),
.A2(n_354),
.B(n_337),
.Y(n_379)
);

AND2x6_ASAP7_75t_L g354 ( 
.A(n_326),
.B(n_293),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_332),
.B(n_310),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_355),
.B(n_361),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_356),
.B(n_357),
.C(n_364),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_330),
.B(n_314),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_338),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_359),
.B(n_308),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_360),
.A2(n_367),
.B1(n_370),
.B2(n_315),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_336),
.B(n_288),
.C(n_289),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_319),
.B(n_287),
.Y(n_365)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_365),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_319),
.B(n_300),
.Y(n_366)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_366),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_341),
.A2(n_286),
.B1(n_297),
.B2(n_298),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_331),
.Y(n_368)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_368),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_338),
.B(n_300),
.Y(n_369)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_369),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_341),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_370)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_331),
.Y(n_372)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_372),
.Y(n_408)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_340),
.Y(n_374)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_374),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_323),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_375),
.B(n_348),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_323),
.B(n_300),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_376),
.B(n_377),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_348),
.B(n_300),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_379),
.A2(n_388),
.B(n_390),
.Y(n_417)
);

OA22x2_ASAP7_75t_L g381 ( 
.A1(n_360),
.A2(n_324),
.B1(n_339),
.B2(n_296),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_381),
.B(n_396),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_371),
.Y(n_382)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_382),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_357),
.B(n_336),
.C(n_345),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_384),
.B(n_363),
.C(n_358),
.Y(n_428)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_385),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_387),
.A2(n_394),
.B1(n_366),
.B2(n_291),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_352),
.A2(n_288),
.B(n_334),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_373),
.A2(n_290),
.B(n_317),
.Y(n_390)
);

XOR2x1_ASAP7_75t_L g392 ( 
.A(n_354),
.B(n_345),
.Y(n_392)
);

OAI21xp33_ASAP7_75t_L g435 ( 
.A1(n_392),
.A2(n_342),
.B(n_335),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_349),
.B(n_333),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_393),
.B(n_395),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_350),
.A2(n_329),
.B1(n_324),
.B2(n_285),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_376),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_354),
.A2(n_339),
.B(n_324),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_397),
.A2(n_370),
.B(n_369),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_365),
.B(n_321),
.Y(n_398)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_398),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_399),
.A2(n_353),
.B1(n_359),
.B2(n_367),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_356),
.B(n_318),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_400),
.B(n_364),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_355),
.B(n_325),
.Y(n_403)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_403),
.Y(n_427)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_404),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_377),
.Y(n_405)
);

O2A1O1Ixp33_ASAP7_75t_L g421 ( 
.A1(n_405),
.A2(n_363),
.B(n_358),
.C(n_321),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_351),
.B(n_353),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_406),
.B(n_372),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_411),
.A2(n_416),
.B1(n_430),
.B2(n_409),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_413),
.A2(n_418),
.B(n_437),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_414),
.B(n_388),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_415),
.A2(n_429),
.B1(n_402),
.B2(n_381),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_407),
.A2(n_375),
.B1(n_378),
.B2(n_374),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_397),
.A2(n_361),
.B(n_368),
.Y(n_418)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_419),
.Y(n_448)
);

AOI32xp33_ASAP7_75t_L g420 ( 
.A1(n_407),
.A2(n_392),
.A3(n_389),
.B1(n_379),
.B2(n_405),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_420),
.B(n_422),
.Y(n_460)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_421),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_389),
.B(n_311),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_383),
.B(n_320),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_423),
.B(n_431),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_398),
.B(n_347),
.Y(n_424)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_424),
.Y(n_450)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_386),
.Y(n_426)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_426),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_428),
.B(n_435),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_387),
.A2(n_316),
.B1(n_325),
.B2(n_371),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_396),
.A2(n_362),
.B1(n_340),
.B2(n_344),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_383),
.B(n_393),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_403),
.Y(n_433)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_433),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_395),
.B(n_302),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_436),
.B(n_400),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_386),
.A2(n_347),
.B(n_284),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_421),
.B(n_391),
.Y(n_440)
);

CKINVDCx14_ASAP7_75t_R g481 ( 
.A(n_440),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_423),
.B(n_431),
.C(n_428),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_441),
.B(n_447),
.C(n_436),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_432),
.B(n_384),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_442),
.B(n_446),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_410),
.B(n_391),
.Y(n_444)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_444),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_445),
.A2(n_459),
.B1(n_413),
.B2(n_418),
.Y(n_466)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_416),
.Y(n_454)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_454),
.Y(n_465)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_434),
.Y(n_455)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_455),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_411),
.A2(n_394),
.B1(n_380),
.B2(n_402),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_456),
.B(n_461),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_457),
.A2(n_429),
.B1(n_381),
.B2(n_409),
.Y(n_473)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_426),
.Y(n_458)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_458),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_415),
.A2(n_381),
.B1(n_390),
.B2(n_401),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_430),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_432),
.B(n_414),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_462),
.B(n_347),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_466),
.A2(n_467),
.B1(n_446),
.B2(n_327),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_445),
.A2(n_425),
.B1(n_412),
.B2(n_427),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_451),
.A2(n_417),
.B(n_425),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_469),
.B(n_244),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_444),
.B(n_401),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_470),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_SL g491 ( 
.A(n_471),
.B(n_462),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_441),
.B(n_417),
.C(n_437),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_472),
.B(n_474),
.C(n_439),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_473),
.A2(n_475),
.B1(n_459),
.B2(n_450),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_443),
.B(n_380),
.C(n_438),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_461),
.A2(n_408),
.B1(n_362),
.B2(n_316),
.Y(n_475)
);

FAx1_ASAP7_75t_L g476 ( 
.A(n_447),
.B(n_408),
.CI(n_362),
.CON(n_476),
.SN(n_476)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_476),
.B(n_479),
.Y(n_482)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_440),
.Y(n_480)
);

AOI22xp33_ASAP7_75t_SL g492 ( 
.A1(n_480),
.A2(n_453),
.B1(n_457),
.B2(n_328),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_474),
.B(n_448),
.Y(n_483)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_483),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_477),
.B(n_442),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_484),
.B(n_485),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_468),
.B(n_460),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_486),
.B(n_494),
.Y(n_502)
);

XNOR2x1_ASAP7_75t_L g507 ( 
.A(n_487),
.B(n_498),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_480),
.A2(n_449),
.B1(n_452),
.B2(n_451),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_489),
.A2(n_469),
.B1(n_467),
.B2(n_476),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_472),
.B(n_439),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_490),
.B(n_491),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_492),
.A2(n_493),
.B1(n_475),
.B2(n_470),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_SL g493 ( 
.A1(n_481),
.A2(n_328),
.B1(n_309),
.B2(n_327),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_468),
.B(n_443),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_495),
.B(n_499),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_477),
.B(n_471),
.C(n_464),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_496),
.B(n_497),
.C(n_282),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_464),
.B(n_245),
.C(n_261),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_466),
.B(n_272),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_490),
.A2(n_487),
.B(n_496),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_505),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_506),
.A2(n_241),
.B1(n_228),
.B2(n_194),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_495),
.B(n_499),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_508),
.B(n_514),
.C(n_484),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_485),
.A2(n_465),
.B1(n_463),
.B2(n_476),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_509),
.B(n_261),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_488),
.A2(n_473),
.B1(n_465),
.B2(n_463),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_510),
.B(n_511),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_482),
.A2(n_478),
.B1(n_245),
.B2(n_282),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_512),
.B(n_515),
.Y(n_521)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_489),
.B(n_478),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g525 ( 
.A1(n_513),
.A2(n_275),
.B(n_241),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_497),
.A2(n_261),
.B1(n_259),
.B2(n_239),
.Y(n_515)
);

INVx5_ASAP7_75t_L g516 ( 
.A(n_507),
.Y(n_516)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_516),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_518),
.B(n_520),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_502),
.B(n_491),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g528 ( 
.A(n_522),
.B(n_524),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_501),
.B(n_259),
.C(n_239),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_523),
.B(n_520),
.C(n_508),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_504),
.B(n_275),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_525),
.B(n_526),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_501),
.B(n_228),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_527),
.B(n_507),
.C(n_500),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_519),
.A2(n_514),
.B(n_513),
.Y(n_530)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_530),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_533),
.B(n_535),
.C(n_523),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_SL g534 ( 
.A(n_517),
.B(n_500),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_SL g538 ( 
.A1(n_534),
.A2(n_518),
.B(n_516),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_536),
.B(n_539),
.C(n_540),
.Y(n_542)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_538),
.Y(n_541)
);

NOR2xp67_ASAP7_75t_L g539 ( 
.A(n_528),
.B(n_531),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_SL g540 ( 
.A1(n_532),
.A2(n_521),
.B(n_509),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_537),
.B(n_535),
.C(n_529),
.Y(n_543)
);

AO221x1_ASAP7_75t_L g544 ( 
.A1(n_543),
.A2(n_541),
.B1(n_542),
.B2(n_526),
.C(n_511),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_SL g546 ( 
.A1(n_544),
.A2(n_545),
.B(n_7),
.Y(n_546)
);

A2O1A1O1Ixp25_ASAP7_75t_L g545 ( 
.A1(n_541),
.A2(n_503),
.B(n_194),
.C(n_15),
.D(n_16),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_546),
.B(n_14),
.Y(n_547)
);

AO21x1_ASAP7_75t_L g548 ( 
.A1(n_547),
.A2(n_15),
.B(n_17),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_548),
.A2(n_15),
.B(n_17),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_549),
.B(n_503),
.Y(n_550)
);


endmodule