module real_jpeg_23931_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_0),
.B(n_49),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_0),
.B(n_40),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_0),
.B(n_52),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_0),
.B(n_84),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_0),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_0),
.B(n_29),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_0),
.B(n_25),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_0),
.B(n_34),
.Y(n_282)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_2),
.B(n_40),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_2),
.B(n_29),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_2),
.B(n_49),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_2),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_2),
.B(n_84),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_2),
.B(n_25),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_4),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_4),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_4),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_4),
.B(n_84),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_4),
.B(n_52),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_4),
.B(n_49),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_4),
.B(n_40),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_4),
.B(n_29),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_5),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_6),
.B(n_84),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_6),
.B(n_52),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_6),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_6),
.B(n_49),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_6),
.B(n_40),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_6),
.B(n_29),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_6),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_6),
.B(n_107),
.Y(n_336)
);

INVx8_ASAP7_75t_SL g27 ( 
.A(n_7),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_8),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_8),
.B(n_25),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_8),
.B(n_29),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_8),
.B(n_17),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_8),
.B(n_84),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_8),
.B(n_52),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_8),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_10),
.B(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_10),
.B(n_29),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_10),
.B(n_40),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_10),
.B(n_17),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_10),
.B(n_84),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_10),
.B(n_52),
.Y(n_264)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_12),
.B(n_52),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_12),
.B(n_49),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_12),
.B(n_84),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_12),
.B(n_17),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_12),
.B(n_40),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_12),
.B(n_29),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_12),
.B(n_25),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_12),
.B(n_300),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_14),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_14),
.B(n_25),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_14),
.B(n_52),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_14),
.B(n_49),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_14),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_14),
.B(n_84),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_29),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_15),
.B(n_34),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_15),
.B(n_49),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_15),
.B(n_40),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_15),
.B(n_236),
.Y(n_235)
);

INVxp33_ASAP7_75t_L g276 ( 
.A(n_15),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_15),
.B(n_52),
.Y(n_312)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_16),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_16),
.B(n_40),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_16),
.B(n_29),
.Y(n_71)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_17),
.Y(n_102)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_17),
.Y(n_145)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_17),
.Y(n_190)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_17),
.Y(n_281)
);

HAxp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_117),
.CON(n_18),
.SN(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_74),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_62),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_43),
.C(n_54),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_22),
.B(n_116),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_23),
.B(n_63),
.Y(n_62)
);

FAx1_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_28),
.CI(n_32),
.CON(n_23),
.SN(n_23)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_26),
.B(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_26),
.B(n_295),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_38),
.C(n_41),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_33),
.B(n_96),
.Y(n_95)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_37),
.Y(n_107)
);

INVx8_ASAP7_75t_L g300 ( 
.A(n_37),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_38),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_40),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_43),
.B(n_54),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_46),
.C(n_51),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_44),
.B(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_45),
.B(n_48),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_46),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_58),
.C(n_60),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_46),
.A2(n_51),
.B1(n_59),
.B2(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_47),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_48),
.B(n_255),
.Y(n_254)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_81),
.B1(n_82),
.B2(n_86),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_51),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_SL g114 ( 
.A(n_51),
.B(n_79),
.C(n_82),
.Y(n_114)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_52),
.Y(n_185)
);

BUFx24_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_60),
.B2(n_61),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_55),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_58),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_72),
.B2(n_73),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_72),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_109),
.C(n_115),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_75),
.A2(n_76),
.B1(n_367),
.B2(n_368),
.Y(n_366)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_95),
.C(n_97),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_77),
.B(n_363),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_87),
.C(n_91),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_78),
.B(n_345),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_82),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_100),
.C(n_103),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_82),
.A2(n_86),
.B1(n_100),
.B2(n_101),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_83),
.B(n_276),
.Y(n_275)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_87),
.B(n_91),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.C(n_90),
.Y(n_87)
);

FAx1_ASAP7_75t_SL g327 ( 
.A(n_88),
.B(n_89),
.CI(n_90),
.CON(n_327),
.SN(n_327)
);

BUFx24_ASAP7_75t_SL g372 ( 
.A(n_91),
.Y(n_372)
);

FAx1_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_93),
.CI(n_94),
.CON(n_91),
.SN(n_91)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_93),
.C(n_94),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_95),
.A2(n_97),
.B1(n_98),
.B2(n_364),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_95),
.Y(n_364)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_105),
.C(n_108),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_99),
.B(n_351),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_100),
.A2(n_101),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_100),
.B(n_304),
.C(n_305),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_103),
.B(n_324),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_105),
.A2(n_106),
.B1(n_108),
.B2(n_337),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_107),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_108),
.A2(n_336),
.B1(n_337),
.B2(n_338),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_108),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_108),
.B(n_333),
.C(n_336),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_109),
.B(n_115),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.C(n_114),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_110),
.A2(n_111),
.B1(n_359),
.B2(n_360),
.Y(n_358)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_113),
.B(n_114),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_365),
.C(n_366),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_353),
.C(n_354),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_341),
.C(n_342),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_317),
.C(n_318),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_284),
.C(n_285),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_247),
.C(n_248),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_215),
.C(n_216),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_195),
.C(n_196),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_155),
.C(n_167),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_140),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_135),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_128),
.B(n_135),
.C(n_140),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.C(n_133),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_130),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_136),
.B(n_138),
.C(n_139),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_148),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_141),
.B(n_149),
.C(n_150),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_142),
.A2(n_143),
.B1(n_146),
.B2(n_147),
.Y(n_166)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_150)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_151),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_152),
.B(n_154),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.C(n_166),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_159),
.A2(n_160),
.B1(n_166),
.B2(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_171)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_166),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_191),
.C(n_192),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_176),
.C(n_181),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_174),
.C(n_175),
.Y(n_191)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.C(n_186),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_184),
.B(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx8_ASAP7_75t_L g236 ( 
.A(n_190),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_209),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_210),
.C(n_214),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_205),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_204),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_204),
.C(n_205),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_200),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_203),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx24_ASAP7_75t_SL g373 ( 
.A(n_205),
.Y(n_373)
);

FAx1_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_207),
.CI(n_208),
.CON(n_205),
.SN(n_205)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_207),
.C(n_208),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_214),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_210),
.Y(n_232)
);

FAx1_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_212),
.CI(n_213),
.CON(n_210),
.SN(n_210)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_231),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_220),
.C(n_231),
.Y(n_247)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_226),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_227),
.C(n_230),
.Y(n_251)
);

BUFx24_ASAP7_75t_SL g369 ( 
.A(n_222),
.Y(n_369)
);

FAx1_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_224),
.CI(n_225),
.CON(n_222),
.SN(n_222)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_223),
.B(n_224),
.C(n_225),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_232),
.B(n_239),
.C(n_245),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_239),
.B1(n_245),
.B2(n_246),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_234),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_237),
.B(n_238),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_237),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_238),
.B(n_272),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_238),
.B(n_272),
.C(n_273),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_239),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_243),
.C(n_244),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_268),
.B2(n_283),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_269),
.C(n_270),
.Y(n_284)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_251),
.B(n_253),
.C(n_261),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_261),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_254),
.B(n_257),
.C(n_260),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_255),
.B(n_293),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_259),
.B2(n_260),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_259),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_267),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_263),
.B(n_266),
.C(n_267),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_265),
.Y(n_266)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_273),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_282),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_275),
.B(n_277),
.C(n_282),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_315),
.B2(n_316),
.Y(n_285)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_286),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_287),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_306),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_288),
.B(n_306),
.C(n_315),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_296),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_289),
.B(n_297),
.C(n_298),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_290),
.B(n_292),
.C(n_294),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_294),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_301),
.B1(n_302),
.B2(n_305),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_299),
.Y(n_305)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_309),
.C(n_310),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_314),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_312),
.B(n_313),
.C(n_314),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_319),
.B(n_321),
.C(n_340),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_328),
.B2(n_340),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_325),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_323),
.B(n_326),
.C(n_327),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

BUFx24_ASAP7_75t_SL g371 ( 
.A(n_327),
.Y(n_371)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_328),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_329),
.B(n_331),
.C(n_332),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_333),
.A2(n_334),
.B1(n_335),
.B2(n_339),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_335),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_336),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_352),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_346),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_344),
.B(n_346),
.C(n_352),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_347),
.B(n_349),
.C(n_350),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_355),
.B(n_357),
.C(n_362),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_358),
.B1(n_361),
.B2(n_362),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_367),
.Y(n_368)
);


endmodule