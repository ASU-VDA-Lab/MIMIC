module fake_jpeg_14159_n_367 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_367);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_367;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_19),
.B(n_6),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_45),
.B(n_56),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_46),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_23),
.B(n_19),
.C(n_31),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_47),
.A2(n_30),
.B(n_40),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_48),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_50),
.Y(n_117)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_52),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_17),
.B(n_6),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_64),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_23),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_69),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_17),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_73),
.Y(n_111)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_71),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_25),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_75),
.Y(n_99)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_42),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_25),
.B(n_5),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_77),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_21),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_100),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_54),
.A2(n_18),
.B1(n_41),
.B2(n_37),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_79),
.A2(n_88),
.B1(n_94),
.B2(n_101),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_26),
.B(n_40),
.C(n_30),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_80),
.A2(n_3),
.B(n_4),
.C(n_11),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_27),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_83),
.B(n_84),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_27),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_55),
.A2(n_18),
.B1(n_41),
.B2(n_37),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_48),
.A2(n_24),
.B1(n_29),
.B2(n_39),
.Y(n_90)
);

OA22x2_ASAP7_75t_L g162 ( 
.A1(n_90),
.A2(n_113),
.B1(n_53),
.B2(n_2),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_93),
.B(n_104),
.C(n_109),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_58),
.A2(n_41),
.B1(n_24),
.B2(n_29),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_42),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_96),
.B(n_97),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_52),
.B(n_24),
.Y(n_97)
);

AOI21xp33_ASAP7_75t_L g98 ( 
.A1(n_59),
.A2(n_28),
.B(n_38),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_98),
.B(n_116),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_51),
.A2(n_29),
.B1(n_32),
.B2(n_36),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_63),
.A2(n_36),
.B1(n_32),
.B2(n_39),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_66),
.A2(n_39),
.B1(n_32),
.B2(n_36),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_107),
.A2(n_112),
.B1(n_53),
.B2(n_1),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_68),
.A2(n_39),
.B1(n_36),
.B2(n_38),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_L g112 ( 
.A1(n_57),
.A2(n_33),
.B1(n_28),
.B2(n_35),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_62),
.A2(n_35),
.B1(n_33),
.B2(n_21),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_15),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_115),
.B(n_118),
.Y(n_149)
);

AOI21xp33_ASAP7_75t_L g116 ( 
.A1(n_59),
.A2(n_5),
.B(n_11),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_50),
.B(n_0),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_71),
.B(n_9),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_120),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_65),
.B(n_12),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_73),
.B(n_12),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_5),
.Y(n_146)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_121),
.Y(n_127)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_128),
.Y(n_177)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_129),
.Y(n_183)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_131),
.B(n_159),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_132),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_133),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_83),
.B(n_75),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_134),
.B(n_155),
.C(n_160),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_102),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_135),
.B(n_165),
.Y(n_176)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_137),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_92),
.A2(n_70),
.B1(n_1),
.B2(n_2),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_138),
.A2(n_140),
.B1(n_156),
.B2(n_136),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_111),
.B1(n_110),
.B2(n_91),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

INVx4_ASAP7_75t_SL g171 ( 
.A(n_142),
.Y(n_171)
);

BUFx6f_ASAP7_75t_SL g143 ( 
.A(n_117),
.Y(n_143)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_144),
.A2(n_162),
.B1(n_166),
.B2(n_107),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_145),
.B(n_146),
.C(n_161),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_85),
.B(n_8),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_147),
.B(n_154),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_153),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_105),
.B(n_8),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_0),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_111),
.A2(n_110),
.B1(n_91),
.B2(n_114),
.Y(n_156)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_114),
.Y(n_158)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_158),
.Y(n_206)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_78),
.B(n_84),
.Y(n_160)
);

AND2x2_ASAP7_75t_SL g163 ( 
.A(n_97),
.B(n_80),
.Y(n_163)
);

AND2x4_ASAP7_75t_SL g200 ( 
.A(n_163),
.B(n_160),
.Y(n_200)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_124),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_93),
.B(n_99),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_109),
.A2(n_4),
.B1(n_12),
.B2(n_0),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_111),
.A2(n_4),
.B(n_87),
.C(n_103),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_81),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_117),
.B(n_123),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_168),
.B(n_87),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_143),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_169),
.B(n_194),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_159),
.A2(n_104),
.B1(n_86),
.B2(n_126),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_174),
.A2(n_190),
.B1(n_201),
.B2(n_205),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_178),
.B(n_185),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_193),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_181),
.A2(n_192),
.B(n_131),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_139),
.B(n_103),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_189),
.Y(n_210)
);

INVx13_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_184),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_149),
.B(n_89),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_141),
.B(n_89),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_187),
.B(n_148),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_139),
.B(n_86),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_157),
.A2(n_126),
.B1(n_106),
.B2(n_123),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_160),
.A2(n_106),
.B(n_81),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_135),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_163),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_195),
.B(n_158),
.Y(n_236)
);

AND2x6_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_152),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_153),
.Y(n_235)
);

XNOR2x1_ASAP7_75t_SL g207 ( 
.A(n_200),
.B(n_199),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_L g201 ( 
.A1(n_151),
.A2(n_162),
.B1(n_167),
.B2(n_129),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_151),
.A2(n_152),
.B1(n_134),
.B2(n_162),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_233),
.Y(n_242)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_180),
.A2(n_162),
.B1(n_134),
.B2(n_145),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_211),
.A2(n_218),
.B1(n_226),
.B2(n_128),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_175),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_225),
.Y(n_241)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_173),
.Y(n_213)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_214),
.Y(n_250)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_215),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_161),
.B1(n_127),
.B2(n_164),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_219),
.Y(n_257)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_220),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_175),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_222),
.B(n_224),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_184),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_194),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_195),
.A2(n_142),
.B1(n_132),
.B2(n_131),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_228),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_229),
.B(n_230),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_176),
.B(n_155),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_231),
.B(n_235),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_182),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_236),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_188),
.B(n_155),
.Y(n_233)
);

O2A1O1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_181),
.A2(n_137),
.B(n_133),
.C(n_130),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_234),
.A2(n_203),
.B(n_206),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_203),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_237),
.A2(n_202),
.B1(n_171),
.B2(n_172),
.Y(n_267)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_239),
.Y(n_254)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_206),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_225),
.A2(n_201),
.B(n_192),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_245),
.A2(n_246),
.B(n_256),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_209),
.A2(n_197),
.B(n_200),
.Y(n_246)
);

AOI322xp5_ASAP7_75t_L g247 ( 
.A1(n_232),
.A2(n_205),
.A3(n_200),
.B1(n_198),
.B2(n_170),
.C1(n_188),
.C2(n_174),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_248),
.Y(n_270)
);

AND2x6_ASAP7_75t_L g248 ( 
.A(n_207),
.B(n_188),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_210),
.B(n_199),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_259),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_209),
.A2(n_179),
.B(n_191),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_263),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_210),
.B(n_190),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_179),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_264),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_216),
.A2(n_191),
.B(n_169),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_211),
.A2(n_177),
.B1(n_191),
.B2(n_202),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_218),
.B(n_177),
.Y(n_265)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_265),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_266),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_267),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_233),
.C(n_229),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_271),
.Y(n_302)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_240),
.Y(n_269)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_269),
.Y(n_296)
);

XOR2x2_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_227),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_226),
.C(n_216),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_280),
.Y(n_295)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_241),
.Y(n_279)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_279),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_216),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_241),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_281),
.B(n_282),
.Y(n_308)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_254),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_254),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_284),
.Y(n_294)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_240),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_252),
.B(n_231),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_287),
.Y(n_299)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_243),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_262),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_288),
.B(n_246),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_261),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_289),
.Y(n_305)
);

AOI21xp33_ASAP7_75t_L g290 ( 
.A1(n_270),
.A2(n_251),
.B(n_252),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_290),
.B(n_273),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_277),
.A2(n_245),
.B(n_264),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_298),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_292),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_275),
.A2(n_266),
.B1(n_265),
.B2(n_244),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_293),
.B(n_307),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_268),
.B(n_248),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_297),
.B(n_304),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_277),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_275),
.A2(n_259),
.B1(n_244),
.B2(n_221),
.Y(n_300)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_300),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_274),
.A2(n_221),
.B1(n_249),
.B2(n_260),
.Y(n_301)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_301),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_258),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_276),
.B(n_253),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_271),
.C(n_283),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_279),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_276),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_311),
.B(n_319),
.Y(n_331)
);

A2O1A1O1Ixp25_ASAP7_75t_L g314 ( 
.A1(n_308),
.A2(n_273),
.B(n_297),
.C(n_281),
.D(n_278),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_314),
.A2(n_308),
.B(n_305),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_315),
.B(n_212),
.Y(n_336)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_294),
.Y(n_316)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_316),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_320),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_302),
.C(n_304),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_318),
.B(n_320),
.C(n_323),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_291),
.B(n_272),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_295),
.B(n_272),
.C(n_282),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_302),
.B(n_274),
.C(n_289),
.Y(n_323)
);

AO221x1_ASAP7_75t_L g324 ( 
.A1(n_303),
.A2(n_217),
.B1(n_287),
.B2(n_243),
.C(n_257),
.Y(n_324)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_324),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_325),
.B(n_330),
.C(n_336),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_326),
.B(n_327),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_312),
.A2(n_293),
.B1(n_305),
.B2(n_307),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_313),
.A2(n_303),
.B1(n_286),
.B2(n_306),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_328),
.A2(n_322),
.B1(n_310),
.B2(n_317),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_296),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_296),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_332),
.B(n_322),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_309),
.A2(n_263),
.B(n_256),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_334),
.A2(n_314),
.B(n_321),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_330),
.B(n_321),
.C(n_319),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_337),
.B(n_339),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_338),
.B(n_343),
.Y(n_353)
);

NAND3xp33_ASAP7_75t_SL g352 ( 
.A(n_341),
.B(n_234),
.C(n_223),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_327),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_342),
.B(n_345),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_329),
.A2(n_269),
.B1(n_284),
.B2(n_260),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_335),
.A2(n_328),
.B1(n_331),
.B2(n_250),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_332),
.B(n_249),
.C(n_253),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_333),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_347),
.B(n_351),
.Y(n_355)
);

OAI21x1_ASAP7_75t_SL g350 ( 
.A1(n_340),
.A2(n_334),
.B(n_333),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_350),
.A2(n_352),
.B(n_354),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_344),
.B(n_325),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_346),
.A2(n_257),
.B(n_250),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_349),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_356),
.B(n_357),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_353),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_348),
.B(n_337),
.C(n_341),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_358),
.A2(n_228),
.B(n_238),
.Y(n_362)
);

AOI322xp5_ASAP7_75t_L g360 ( 
.A1(n_357),
.A2(n_353),
.A3(n_215),
.B1(n_208),
.B2(n_213),
.C1(n_214),
.C2(n_220),
.Y(n_360)
);

AOI322xp5_ASAP7_75t_L g364 ( 
.A1(n_360),
.A2(n_219),
.A3(n_239),
.B1(n_223),
.B2(n_361),
.C1(n_237),
.C2(n_172),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_362),
.A2(n_359),
.B(n_355),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_363),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_365),
.A2(n_364),
.B(n_237),
.Y(n_366)
);

FAx1_ASAP7_75t_SL g367 ( 
.A(n_366),
.B(n_171),
.CI(n_361),
.CON(n_367),
.SN(n_367)
);


endmodule