module real_aes_13745_n_16 (n_13, n_4, n_0, n_3, n_5, n_2, n_15, n_7, n_8, n_6, n_9, n_12, n_1, n_14, n_10, n_11, n_16);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_15;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_14;
input n_10;
input n_11;
output n_16;
wire n_17;
wire n_28;
wire n_22;
wire n_24;
wire n_41;
wire n_34;
wire n_19;
wire n_40;
wire n_49;
wire n_46;
wire n_53;
wire n_25;
wire n_47;
wire n_48;
wire n_43;
wire n_32;
wire n_30;
wire n_51;
wire n_37;
wire n_54;
wire n_35;
wire n_42;
wire n_39;
wire n_45;
wire n_27;
wire n_50;
wire n_38;
wire n_23;
wire n_29;
wire n_20;
wire n_52;
wire n_44;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
NOR3xp33_ASAP7_75t_SL g23 ( .A(n_0), .B(n_9), .C(n_24), .Y(n_23) );
INVx1_ASAP7_75t_L g29 ( .A(n_1), .Y(n_29) );
NOR2xp33_ASAP7_75t_R g18 ( .A(n_2), .B(n_19), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g38 ( .A(n_2), .Y(n_38) );
NOR2xp33_ASAP7_75t_R g26 ( .A(n_3), .B(n_14), .Y(n_26) );
CKINVDCx5p33_ASAP7_75t_R g35 ( .A(n_3), .Y(n_35) );
NAND2xp33_ASAP7_75t_R g47 ( .A(n_3), .B(n_14), .Y(n_47) );
NOR2xp33_ASAP7_75t_R g50 ( .A(n_3), .B(n_51), .Y(n_50) );
CKINVDCx5p33_ASAP7_75t_R g40 ( .A(n_4), .Y(n_40) );
CKINVDCx5p33_ASAP7_75t_R g20 ( .A(n_5), .Y(n_20) );
NAND5xp2_ASAP7_75t_SL g36 ( .A(n_5), .B(n_8), .C(n_37), .D(n_38), .E(n_39), .Y(n_36) );
CKINVDCx20_ASAP7_75t_R g52 ( .A(n_6), .Y(n_52) );
CKINVDCx20_ASAP7_75t_R g54 ( .A(n_7), .Y(n_54) );
NOR2xp33_ASAP7_75t_R g21 ( .A(n_8), .B(n_22), .Y(n_21) );
CKINVDCx5p33_ASAP7_75t_R g25 ( .A(n_10), .Y(n_25) );
AOI221xp5_ASAP7_75t_R g41 ( .A1(n_11), .A2(n_13), .B1(n_42), .B2(n_45), .C(n_48), .Y(n_41) );
NAND3xp33_ASAP7_75t_SL g19 ( .A(n_12), .B(n_20), .C(n_21), .Y(n_19) );
CKINVDCx5p33_ASAP7_75t_R g39 ( .A(n_12), .Y(n_39) );
NOR2xp33_ASAP7_75t_R g34 ( .A(n_14), .B(n_35), .Y(n_34) );
CKINVDCx5p33_ASAP7_75t_R g51 ( .A(n_14), .Y(n_51) );
CKINVDCx5p33_ASAP7_75t_R g24 ( .A(n_15), .Y(n_24) );
OAI221xp5_ASAP7_75t_L g16 ( .A1(n_17), .A2(n_27), .B1(n_30), .B2(n_40), .C(n_41), .Y(n_16) );
NAND2xp33_ASAP7_75t_R g17 ( .A(n_18), .B(n_26), .Y(n_17) );
NAND2xp33_ASAP7_75t_R g53 ( .A(n_18), .B(n_50), .Y(n_53) );
CKINVDCx5p33_ASAP7_75t_R g37 ( .A(n_22), .Y(n_37) );
NAND2xp33_ASAP7_75t_R g22 ( .A(n_23), .B(n_25), .Y(n_22) );
NAND2xp33_ASAP7_75t_R g43 ( .A(n_26), .B(n_44), .Y(n_43) );
CKINVDCx5p33_ASAP7_75t_R g27 ( .A(n_28), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_29), .Y(n_28) );
CKINVDCx20_ASAP7_75t_R g30 ( .A(n_31), .Y(n_30) );
HB1xp67_ASAP7_75t_L g31 ( .A(n_32), .Y(n_31) );
NOR2xp33_ASAP7_75t_R g32 ( .A(n_33), .B(n_36), .Y(n_32) );
CKINVDCx5p33_ASAP7_75t_R g33 ( .A(n_34), .Y(n_33) );
CKINVDCx5p33_ASAP7_75t_R g44 ( .A(n_36), .Y(n_44) );
NOR2xp33_ASAP7_75t_R g46 ( .A(n_36), .B(n_47), .Y(n_46) );
CKINVDCx5p33_ASAP7_75t_R g42 ( .A(n_43), .Y(n_42) );
NAND2xp33_ASAP7_75t_R g49 ( .A(n_44), .B(n_50), .Y(n_49) );
HB1xp67_ASAP7_75t_L g45 ( .A(n_46), .Y(n_45) );
OAI22xp33_ASAP7_75t_R g48 ( .A1(n_49), .A2(n_52), .B1(n_53), .B2(n_54), .Y(n_48) );
endmodule