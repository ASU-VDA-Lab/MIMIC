module fake_jpeg_7107_n_73 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_73);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_73;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_9),
.B(n_7),
.Y(n_10)
);

INVx2_ASAP7_75t_SL g11 ( 
.A(n_5),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx12f_ASAP7_75t_SL g14 ( 
.A(n_9),
.Y(n_14)
);

INVx6_ASAP7_75t_SL g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_0),
.B(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_21),
.B(n_23),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_24),
.Y(n_31)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx9p33_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_11),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_27),
.A2(n_10),
.B1(n_19),
.B2(n_12),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_16),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_33),
.Y(n_48)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_34),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_18),
.C(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_SL g40 ( 
.A(n_36),
.B(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_28),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_32),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_26),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_46),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_24),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_42),
.C(n_39),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_31),
.B(n_10),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_29),
.B1(n_37),
.B2(n_12),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_36),
.B1(n_29),
.B2(n_24),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_51),
.B(n_48),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_53),
.C(n_54),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_34),
.C(n_30),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_12),
.B1(n_20),
.B2(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_50),
.B1(n_20),
.B2(n_17),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_45),
.C(n_28),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_62),
.C(n_54),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_45),
.C(n_28),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_64),
.C(n_17),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_59),
.C(n_60),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_58),
.B(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_66),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_69),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_64),
.A2(n_3),
.B(n_4),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_1),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_2),
.C(n_3),
.Y(n_72)
);

OR3x1_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_8),
.C(n_70),
.Y(n_73)
);


endmodule