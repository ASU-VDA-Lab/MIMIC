module fake_jpeg_19131_n_81 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_81);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_81;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_24),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_18),
.Y(n_44)
);

CKINVDCx9p33_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_26),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_51),
.Y(n_57)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_49),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_59),
.A2(n_36),
.B1(n_52),
.B2(n_43),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_50),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_30),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_62),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_42),
.B(n_41),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_37),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_34),
.B1(n_54),
.B2(n_29),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_70),
.Y(n_72)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_71),
.A2(n_39),
.B(n_28),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_9),
.B(n_12),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_8),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_74),
.B(n_13),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_76),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_14),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_17),
.B(n_19),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_77),
.C(n_38),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_20),
.Y(n_81)
);


endmodule