module fake_ibex_232_n_16 (n_3, n_1, n_4, n_2, n_0, n_16);

input n_3;
input n_1;
input n_4;
input n_2;
input n_0;

output n_16;



endmodule