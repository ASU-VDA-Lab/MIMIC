module fake_jpeg_13746_n_150 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_150);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_15),
.B(n_28),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_19),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_30),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_27),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_25),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_33),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_7),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_17),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_44),
.Y(n_62)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_64),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

CKINVDCx6p67_ASAP7_75t_R g84 ( 
.A(n_66),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_69),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_1),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_2),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_51),
.B1(n_58),
.B2(n_46),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_76),
.A2(n_22),
.B1(n_42),
.B2(n_41),
.Y(n_98)
);

BUFx10_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

BUFx24_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_80),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_56),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_48),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_82),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_45),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_62),
.A2(n_59),
.B(n_57),
.Y(n_83)
);

OAI32xp33_ASAP7_75t_L g89 ( 
.A1(n_83),
.A2(n_51),
.A3(n_58),
.B1(n_49),
.B2(n_55),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_77),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_90),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_84),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_89),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_79),
.C(n_80),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_84),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_94),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_53),
.C(n_61),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_93),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_54),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_66),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_23),
.Y(n_116)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_6),
.Y(n_117)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

NAND2x1_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_3),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_3),
.B(n_4),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_85),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_103),
.B(n_115),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_108),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_110),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_101),
.B(n_4),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_97),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_116),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_101),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_21),
.B1(n_24),
.B2(n_26),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_5),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_31),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_105),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_13),
.C(n_14),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_123),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_16),
.C(n_20),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_125),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_106),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_127),
.A2(n_128),
.B(n_130),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_34),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_102),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_36),
.B(n_37),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_120),
.A2(n_114),
.B1(n_118),
.B2(n_43),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_128),
.C(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_138),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_119),
.Y(n_140)
);

NOR3xp33_ASAP7_75t_SL g143 ( 
.A(n_140),
.B(n_141),
.C(n_131),
.Y(n_143)
);

AND2x4_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_119),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_136),
.B(n_134),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_139),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_142),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_135),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_147),
.B(n_38),
.Y(n_148)
);

FAx1_ASAP7_75t_SL g149 ( 
.A(n_148),
.B(n_39),
.CI(n_114),
.CON(n_149),
.SN(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_118),
.Y(n_150)
);


endmodule