module fake_jpeg_31823_n_63 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_63);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_63;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_43;
wire n_50;
wire n_37;
wire n_32;

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_30),
.Y(n_37)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_32),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_35),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_32),
.B(n_2),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_6),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_27),
.B1(n_13),
.B2(n_14),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_43),
.B1(n_6),
.B2(n_7),
.Y(n_49)
);

A2O1A1O1Ixp25_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_12),
.B(n_22),
.C(n_21),
.D(n_20),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_10),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_31),
.A2(n_27),
.B1(n_3),
.B2(n_4),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_35),
.B1(n_4),
.B2(n_5),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_49),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_2),
.B(n_5),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_46),
.Y(n_56)
);

OA21x2_ASAP7_75t_SL g52 ( 
.A1(n_47),
.A2(n_50),
.B(n_38),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_16),
.B1(n_18),
.B2(n_17),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_48),
.A2(n_41),
.B1(n_42),
.B2(n_36),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_7),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_53),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_40),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_54),
.A2(n_55),
.B(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_58),
.Y(n_61)
);

HAxp5_ASAP7_75t_SL g58 ( 
.A(n_56),
.B(n_8),
.CON(n_58),
.SN(n_58)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_55),
.Y(n_60)
);

A2O1A1O1Ixp25_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_51),
.B(n_53),
.C(n_54),
.D(n_8),
.Y(n_62)
);

A2O1A1O1Ixp25_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_61),
.B(n_19),
.C(n_11),
.D(n_60),
.Y(n_63)
);


endmodule