module fake_jpeg_20966_n_204 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_204);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_31),
.Y(n_39)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_20),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_32),
.A2(n_21),
.B1(n_16),
.B2(n_15),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_30),
.B1(n_24),
.B2(n_26),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_21),
.B1(n_25),
.B2(n_24),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_41),
.B1(n_42),
.B2(n_23),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_34),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_27),
.A2(n_21),
.B1(n_14),
.B2(n_19),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_29),
.A2(n_21),
.B1(n_25),
.B2(n_24),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_19),
.C(n_14),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_47),
.C(n_42),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_35),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_62),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_52),
.B(n_54),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_53),
.A2(n_58),
.B1(n_66),
.B2(n_70),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_55),
.A2(n_43),
.B1(n_44),
.B2(n_20),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_16),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_56),
.B(n_57),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_16),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_38),
.B1(n_40),
.B2(n_49),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_68),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_15),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_61),
.B(n_0),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_47),
.B(n_15),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_63),
.B(n_51),
.Y(n_82)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_64),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_26),
.B1(n_25),
.B2(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_69),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_26),
.B1(n_23),
.B2(n_17),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_17),
.B1(n_35),
.B2(n_19),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_53),
.B1(n_58),
.B2(n_43),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_90),
.Y(n_99)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_84),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_46),
.C(n_37),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_67),
.C(n_65),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_17),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_78),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_44),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_79),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_82),
.B(n_85),
.Y(n_109)
);

NAND3xp33_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_8),
.C(n_12),
.Y(n_85)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_20),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_86),
.A2(n_92),
.B(n_1),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_54),
.A2(n_20),
.B1(n_19),
.B2(n_14),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_89),
.Y(n_96)
);

AOI22x1_ASAP7_75t_L g89 ( 
.A1(n_51),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_0),
.Y(n_92)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_101),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_60),
.C(n_2),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_1),
.B(n_3),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_89),
.B(n_82),
.Y(n_124)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_83),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_107),
.B(n_111),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_110),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_6),
.C(n_3),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_83),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_113),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_107),
.Y(n_121)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_115),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_77),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_116),
.B(n_117),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_80),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_1),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_118),
.B(n_92),
.Y(n_136)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_93),
.B1(n_73),
.B2(n_86),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_123),
.A2(n_131),
.B1(n_137),
.B2(n_96),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_136),
.Y(n_140)
);

NOR3xp33_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_89),
.C(n_95),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_99),
.A2(n_93),
.B1(n_95),
.B2(n_92),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_74),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_132),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_72),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_133),
.B(n_134),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_109),
.B(n_97),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_99),
.A2(n_88),
.B1(n_5),
.B2(n_7),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_96),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_137),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_141),
.B(n_147),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_98),
.C(n_118),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_144),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_103),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_145),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_101),
.C(n_108),
.Y(n_147)
);

FAx1_ASAP7_75t_SL g148 ( 
.A(n_130),
.B(n_110),
.CI(n_100),
.CON(n_148),
.SN(n_148)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_154),
.Y(n_163)
);

BUFx12_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

INVx13_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_152),
.A2(n_105),
.B1(n_135),
.B2(n_119),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_153),
.Y(n_162)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_106),
.C(n_104),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_155),
.B(n_143),
.Y(n_167)
);

AOI322xp5_ASAP7_75t_L g156 ( 
.A1(n_151),
.A2(n_124),
.A3(n_126),
.B1(n_135),
.B2(n_102),
.C1(n_128),
.C2(n_129),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_156),
.A2(n_151),
.B(n_140),
.Y(n_170)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_126),
.B1(n_120),
.B2(n_128),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_160),
.A2(n_153),
.B1(n_146),
.B2(n_141),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_155),
.A2(n_129),
.B1(n_139),
.B2(n_113),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_164),
.A2(n_146),
.B(n_142),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_144),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_171),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_157),
.C(n_148),
.Y(n_184)
);

NOR2xp67_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_148),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_173),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_147),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_166),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_162),
.Y(n_175)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_177),
.A2(n_162),
.B(n_163),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_166),
.C(n_161),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_181),
.C(n_182),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_168),
.Y(n_179)
);

INVxp67_ASAP7_75t_SL g186 ( 
.A(n_179),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_171),
.C(n_169),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_191),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_160),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_190),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_176),
.C(n_164),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_185),
.A2(n_173),
.B(n_140),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_182),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_180),
.Y(n_198)
);

OAI321xp33_ASAP7_75t_L g194 ( 
.A1(n_186),
.A2(n_154),
.A3(n_150),
.B1(n_158),
.B2(n_180),
.C(n_112),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_158),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_196),
.B(n_197),
.Y(n_199)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_195),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_198),
.B(n_192),
.C(n_150),
.Y(n_200)
);

AOI321xp33_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_197),
.A3(n_150),
.B1(n_115),
.B2(n_114),
.C(n_11),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_201),
.A2(n_199),
.B(n_9),
.Y(n_202)
);

AOI321xp33_ASAP7_75t_L g203 ( 
.A1(n_202),
.A2(n_4),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C(n_114),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_4),
.Y(n_204)
);


endmodule