module real_jpeg_9737_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_0),
.A2(n_1),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_0),
.A2(n_27),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g21 ( 
.A1(n_1),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_1),
.B(n_22),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_2),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_2),
.B(n_61),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_4),
.A2(n_43),
.B1(n_46),
.B2(n_52),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_L g121 ( 
.A1(n_4),
.A2(n_9),
.B(n_43),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_5),
.A2(n_6),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_5),
.A2(n_25),
.B(n_31),
.C(n_35),
.Y(n_34)
);

NAND2xp33_ASAP7_75t_SL g35 ( 
.A(n_5),
.B(n_25),
.Y(n_35)
);

OAI32xp33_ASAP7_75t_L g142 ( 
.A1(n_5),
.A2(n_6),
.A3(n_25),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_6),
.A2(n_52),
.B(n_53),
.C(n_54),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_6),
.B(n_52),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_6),
.A2(n_9),
.B1(n_28),
.B2(n_33),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_6),
.A2(n_10),
.B1(n_33),
.B2(n_47),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_6),
.A2(n_28),
.B(n_52),
.C(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_7),
.Y(n_22)
);

HAxp5_ASAP7_75t_SL g27 ( 
.A(n_7),
.B(n_28),
.CON(n_27),
.SN(n_27)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_8),
.A2(n_43),
.B1(n_46),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_9),
.A2(n_25),
.B(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_9),
.B(n_25),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_9),
.A2(n_28),
.B1(n_43),
.B2(n_46),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_9),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_9),
.B(n_31),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_10),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_89),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_87),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_73),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_14),
.B(n_73),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_65),
.Y(n_14)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_57),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_40),
.B2(n_56),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_17),
.A2(n_18),
.B1(n_66),
.B2(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_17),
.A2(n_18),
.B1(n_81),
.B2(n_82),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_29),
.B1(n_38),
.B2(n_39),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_19),
.B(n_39),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_19),
.B(n_39),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_19),
.A2(n_38),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_27),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_24),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_24),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_25),
.B(n_26),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_28),
.B(n_54),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_28),
.B(n_44),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_29),
.A2(n_39),
.B1(n_50),
.B2(n_79),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_29),
.B(n_86),
.C(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_29),
.A2(n_39),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_36),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_32),
.B(n_33),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_37),
.Y(n_143)
);

AOI211xp5_ASAP7_75t_SL g94 ( 
.A1(n_38),
.A2(n_50),
.B(n_72),
.C(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_39),
.B(n_79),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_39),
.A2(n_79),
.B(n_146),
.C(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_50),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_41),
.A2(n_50),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_41),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_45),
.B2(n_48),
.Y(n_41)
);

INVxp33_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_44),
.B1(n_45),
.B2(n_68),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_42),
.A2(n_44),
.B(n_68),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_46),
.B(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_48),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_67),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_50),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_50),
.A2(n_67),
.B1(n_79),
.B2(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_50),
.A2(n_79),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_50),
.A2(n_79),
.B1(n_120),
.B2(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_50),
.B(n_86),
.C(n_124),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_50),
.A2(n_79),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_50),
.B(n_152),
.C(n_158),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_54),
.B(n_55),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_51),
.A2(n_54),
.B1(n_55),
.B2(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_62),
.B2(n_64),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_62),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_69),
.B(n_71),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_66),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_67),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_72),
.B(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.C(n_80),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_74),
.A2(n_75),
.B1(n_77),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_77),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_120),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_80),
.B(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_86),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_83),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_86),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_86),
.A2(n_107),
.B1(n_123),
.B2(n_126),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_86),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_86),
.B(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_86),
.A2(n_107),
.B1(n_142),
.B2(n_145),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_86),
.A2(n_107),
.B1(n_110),
.B2(n_111),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_86),
.B(n_142),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_113),
.B(n_169),
.C(n_174),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_100),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_91),
.B(n_100),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_99),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_93),
.B(n_97),
.C(n_99),
.Y(n_170)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_95),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.C(n_109),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_101),
.A2(n_102),
.B1(n_164),
.B2(n_166),
.Y(n_163)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_103),
.A2(n_104),
.B1(n_141),
.B2(n_146),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_105),
.A2(n_106),
.B1(n_109),
.B2(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_107),
.B(n_135),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_109),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_168),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_161),
.B(n_167),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_148),
.B(n_160),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_138),
.B(n_147),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_127),
.B(n_137),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_122),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_120),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_123),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_134),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_140),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_141),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_142),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_149),
.B(n_151),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_156),
.B2(n_157),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_162),
.B(n_163),
.Y(n_167)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_164),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_170),
.B(n_171),
.Y(n_174)
);


endmodule