module fake_jpeg_17659_n_314 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_314);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_31),
.B(n_8),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_44),
.Y(n_69)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_29),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_34),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_32),
.Y(n_55)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_18),
.B1(n_25),
.B2(n_27),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_52),
.B1(n_53),
.B2(n_60),
.Y(n_72)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_31),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_55),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_27),
.B(n_24),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_L g75 ( 
.A1(n_51),
.A2(n_45),
.B(n_23),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_25),
.B1(n_31),
.B2(n_32),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_25),
.B1(n_33),
.B2(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_59),
.B(n_66),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_32),
.B1(n_33),
.B2(n_17),
.Y(n_60)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_38),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_67),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_23),
.B1(n_30),
.B2(n_21),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_65),
.A2(n_20),
.B1(n_30),
.B2(n_17),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_38),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_74),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_58),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_84),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_44),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_76),
.B(n_82),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_78),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_46),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_79),
.A2(n_56),
.B1(n_48),
.B2(n_67),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_88),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_62),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_59),
.A2(n_21),
.B1(n_20),
.B2(n_19),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_83),
.A2(n_49),
.B1(n_1),
.B2(n_2),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_40),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_28),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_26),
.Y(n_89)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_60),
.B(n_28),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_99),
.Y(n_122)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_101),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_57),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_28),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_102),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_85),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_103),
.B(n_118),
.Y(n_153)
);

INVx5_ASAP7_75t_SL g107 ( 
.A(n_90),
.Y(n_107)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_81),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_110),
.B(n_116),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_95),
.A2(n_56),
.B1(n_63),
.B2(n_41),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_119),
.B1(n_124),
.B2(n_121),
.Y(n_137)
);

BUFx24_ASAP7_75t_SL g118 ( 
.A(n_87),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_72),
.A2(n_56),
.B1(n_49),
.B2(n_64),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_120),
.A2(n_16),
.B(n_4),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_82),
.A2(n_47),
.B1(n_43),
.B2(n_68),
.Y(n_124)
);

AND2x6_ASAP7_75t_L g125 ( 
.A(n_73),
.B(n_12),
.Y(n_125)
);

A2O1A1O1Ixp25_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_87),
.B(n_1),
.C(n_2),
.D(n_3),
.Y(n_139)
);

NAND3xp33_ASAP7_75t_L g126 ( 
.A(n_84),
.B(n_26),
.C(n_1),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_126),
.B(n_130),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_76),
.A2(n_43),
.B(n_26),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_124),
.C(n_114),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_86),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_104),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_132),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_104),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_133),
.B(n_136),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_134),
.A2(n_129),
.B(n_113),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_123),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_137),
.A2(n_147),
.B1(n_152),
.B2(n_154),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_89),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_141),
.C(n_35),
.Y(n_181)
);

OAI21xp33_ASAP7_75t_SL g189 ( 
.A1(n_139),
.A2(n_161),
.B(n_4),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_43),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_112),
.A2(n_80),
.B1(n_70),
.B2(n_93),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_142),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_105),
.B(n_86),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_144),
.B(n_160),
.Y(n_175)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_100),
.B1(n_70),
.B2(n_91),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_101),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_155),
.Y(n_166)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_149),
.Y(n_191)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_151),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_122),
.A2(n_117),
.B1(n_111),
.B2(n_105),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_91),
.B1(n_97),
.B2(n_78),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_26),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_103),
.Y(n_156)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_115),
.B(n_26),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_159),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_110),
.B(n_22),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_158),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_115),
.B(n_77),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_130),
.B(n_16),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_22),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_162),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_149),
.A2(n_125),
.B1(n_113),
.B2(n_120),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_164),
.A2(n_174),
.B1(n_194),
.B2(n_154),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_155),
.A2(n_125),
.B(n_108),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_167),
.A2(n_183),
.B(n_6),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_145),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_186),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_170),
.B(n_181),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_150),
.A2(n_107),
.B(n_24),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_171),
.A2(n_176),
.B(n_147),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_134),
.A2(n_113),
.B1(n_99),
.B2(n_107),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_132),
.A2(n_24),
.B(n_28),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_152),
.B(n_22),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_135),
.Y(n_196)
);

OAI32xp33_ASAP7_75t_L g180 ( 
.A1(n_148),
.A2(n_28),
.A3(n_35),
.B1(n_106),
.B2(n_0),
.Y(n_180)
);

AOI221xp5_ASAP7_75t_L g210 ( 
.A1(n_180),
.A2(n_189),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_35),
.Y(n_183)
);

AND2x4_ASAP7_75t_SL g185 ( 
.A(n_142),
.B(n_128),
.Y(n_185)
);

NAND2x1_ASAP7_75t_SL g198 ( 
.A(n_185),
.B(n_156),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_156),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_138),
.B(n_106),
.Y(n_187)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_141),
.B(n_96),
.Y(n_190)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_190),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_159),
.Y(n_192)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_192),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_137),
.A2(n_92),
.B1(n_85),
.B2(n_98),
.Y(n_194)
);

AO21x1_ASAP7_75t_L g237 ( 
.A1(n_196),
.A2(n_198),
.B(n_210),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_188),
.Y(n_197)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_197),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_199),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_201),
.A2(n_206),
.B1(n_208),
.B2(n_215),
.Y(n_225)
);

BUFx12f_ASAP7_75t_SL g202 ( 
.A(n_185),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_202),
.A2(n_207),
.B(n_219),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_183),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_213),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_151),
.Y(n_205)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_205),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_163),
.A2(n_139),
.B1(n_140),
.B2(n_143),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_191),
.A2(n_140),
.B1(n_161),
.B2(n_153),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_195),
.Y(n_209)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_92),
.Y(n_212)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_212),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_165),
.B(n_6),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_96),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_217),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_184),
.A2(n_96),
.B1(n_90),
.B2(n_10),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_90),
.Y(n_217)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_185),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_218),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_167),
.A2(n_7),
.B(n_11),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_220),
.A2(n_221),
.B1(n_175),
.B2(n_169),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_193),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_202),
.A2(n_184),
.B1(n_164),
.B2(n_166),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_224),
.A2(n_234),
.B1(n_243),
.B2(n_244),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_187),
.C(n_181),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_231),
.C(n_211),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_190),
.C(n_170),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_232),
.A2(n_239),
.B1(n_200),
.B2(n_196),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_182),
.Y(n_233)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_233),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_218),
.A2(n_166),
.B1(n_185),
.B2(n_174),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_192),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_242),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_208),
.A2(n_193),
.B1(n_173),
.B2(n_169),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_171),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_204),
.A2(n_182),
.B1(n_194),
.B2(n_180),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_211),
.A2(n_216),
.B1(n_203),
.B2(n_198),
.Y(n_244)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

BUFx24_ASAP7_75t_SL g247 ( 
.A(n_226),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_256),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_244),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_251),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_223),
.A2(n_206),
.B(n_207),
.Y(n_250)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_217),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_245),
.A2(n_220),
.B1(n_219),
.B2(n_215),
.Y(n_253)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_259),
.C(n_224),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_231),
.B(n_198),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_242),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_225),
.A2(n_209),
.B1(n_195),
.B2(n_186),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_245),
.A2(n_179),
.B(n_165),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_258),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_223),
.A2(n_172),
.B1(n_175),
.B2(n_209),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_176),
.C(n_11),
.Y(n_259)
);

BUFx12_ASAP7_75t_L g262 ( 
.A(n_230),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_262),
.B(n_263),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_233),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_272),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_268),
.B(n_263),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_236),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_251),
.B(n_241),
.Y(n_273)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_273),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_234),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_276),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_254),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_237),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_277),
.B(n_237),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_262),
.Y(n_279)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_271),
.A2(n_248),
.B(n_269),
.Y(n_280)
);

AOI21xp33_ASAP7_75t_L g293 ( 
.A1(n_280),
.A2(n_252),
.B(n_256),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_283),
.C(n_238),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_262),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_286),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_227),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_287),
.A2(n_274),
.B1(n_272),
.B2(n_276),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_264),
.A2(n_260),
.B(n_261),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_288),
.A2(n_240),
.B(n_227),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_240),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_7),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_291),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_284),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_265),
.C(n_235),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_297),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_296),
.B(n_298),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_235),
.C(n_238),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_300),
.B(n_302),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_286),
.Y(n_302)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_292),
.Y(n_303)
);

AOI322xp5_ASAP7_75t_L g309 ( 
.A1(n_303),
.A2(n_305),
.A3(n_12),
.B1(n_14),
.B2(n_15),
.C1(n_278),
.C2(n_304),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_280),
.Y(n_305)
);

AOI322xp5_ASAP7_75t_L g307 ( 
.A1(n_303),
.A2(n_287),
.A3(n_294),
.B1(n_278),
.B2(n_14),
.C1(n_7),
.C2(n_13),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_307),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_299),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_309),
.C(n_301),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_311),
.A2(n_306),
.B(n_300),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_312),
.A2(n_310),
.B1(n_14),
.B2(n_15),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_12),
.Y(n_314)
);


endmodule