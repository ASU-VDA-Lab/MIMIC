module real_aes_9371_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
NAND2xp5_ASAP7_75t_L g545 ( .A(n_0), .B(n_58), .Y(n_545) );
INVx1_ASAP7_75t_L g570 ( .A(n_0), .Y(n_570) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_0), .Y(n_591) );
AND2x2_ASAP7_75t_L g602 ( .A(n_0), .B(n_569), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_1), .B(n_145), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_2), .B(n_111), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g678 ( .A(n_3), .Y(n_678) );
INVx2_ASAP7_75t_L g484 ( .A(n_4), .Y(n_484) );
BUFx2_ASAP7_75t_L g532 ( .A(n_5), .Y(n_532) );
BUFx2_ASAP7_75t_L g641 ( .A(n_5), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_6), .A2(n_48), .B1(n_581), .B2(n_582), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_6), .A2(n_48), .B1(n_635), .B2(n_637), .Y(n_634) );
AOI221xp5_ASAP7_75t_L g583 ( .A1(n_7), .A2(n_36), .B1(n_584), .B2(n_588), .C(n_590), .Y(n_583) );
INVx1_ASAP7_75t_L g628 ( .A(n_7), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_8), .B(n_108), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_9), .B(n_90), .Y(n_206) );
NAND2x1p5_ASAP7_75t_L g151 ( .A(n_10), .B(n_90), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_11), .B(n_213), .Y(n_231) );
AND2x2_ASAP7_75t_L g182 ( .A(n_12), .B(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g609 ( .A(n_13), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_13), .A2(n_44), .B1(n_635), .B2(n_648), .Y(n_647) );
CKINVDCx5p33_ASAP7_75t_R g673 ( .A(n_14), .Y(n_673) );
BUFx6f_ASAP7_75t_L g103 ( .A(n_15), .Y(n_103) );
NAND2xp5_ASAP7_75t_SL g118 ( .A(n_16), .B(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_17), .B(n_138), .Y(n_218) );
NAND2xp33_ASAP7_75t_L g146 ( .A(n_18), .B(n_147), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g604 ( .A(n_19), .Y(n_604) );
NAND2xp33_ASAP7_75t_L g204 ( .A(n_20), .B(n_147), .Y(n_204) );
BUFx6f_ASAP7_75t_L g100 ( .A(n_21), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_22), .Y(n_160) );
INVx1_ASAP7_75t_L g530 ( .A(n_23), .Y(n_530) );
INVx1_ASAP7_75t_L g701 ( .A(n_23), .Y(n_701) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_24), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_25), .B(n_110), .Y(n_150) );
OAI21x1_ASAP7_75t_L g92 ( .A1(n_26), .A2(n_52), .B(n_93), .Y(n_92) );
A2O1A1Ixp33_ASAP7_75t_L g187 ( .A1(n_27), .A2(n_131), .B(n_188), .C(n_190), .Y(n_187) );
INVx1_ASAP7_75t_L g510 ( .A(n_28), .Y(n_510) );
OAI221xp5_ASAP7_75t_L g571 ( .A1(n_28), .A2(n_50), .B1(n_572), .B2(n_577), .C(n_579), .Y(n_571) );
CKINVDCx5p33_ASAP7_75t_R g661 ( .A(n_29), .Y(n_661) );
INVx1_ASAP7_75t_L g497 ( .A(n_30), .Y(n_497) );
AOI221xp5_ASAP7_75t_L g546 ( .A1(n_30), .A2(n_46), .B1(n_547), .B2(n_552), .C(n_557), .Y(n_546) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_31), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g101 ( .A(n_32), .B(n_102), .Y(n_101) );
NAND2xp33_ASAP7_75t_L g234 ( .A(n_33), .B(n_167), .Y(n_234) );
AND2x6_ASAP7_75t_L g116 ( .A(n_34), .B(n_117), .Y(n_116) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_34), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_34), .B(n_654), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_35), .B(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g633 ( .A(n_36), .Y(n_633) );
XNOR2xp5_ASAP7_75t_L g474 ( .A(n_37), .B(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_38), .B(n_189), .Y(n_203) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_38), .Y(n_703) );
NAND2xp33_ASAP7_75t_L g217 ( .A(n_39), .B(n_167), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g598 ( .A(n_40), .Y(n_598) );
INVx1_ASAP7_75t_L g117 ( .A(n_41), .Y(n_117) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_41), .Y(n_654) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_42), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_43), .B(n_167), .Y(n_230) );
INVx1_ASAP7_75t_L g607 ( .A(n_44), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_45), .Y(n_96) );
INVx1_ASAP7_75t_L g524 ( .A(n_46), .Y(n_524) );
AND2x2_ASAP7_75t_L g192 ( .A(n_47), .B(n_138), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_49), .B(n_129), .Y(n_128) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_49), .Y(n_672) );
INVx1_ASAP7_75t_L g516 ( .A(n_50), .Y(n_516) );
INVx2_ASAP7_75t_L g540 ( .A(n_51), .Y(n_540) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_53), .Y(n_149) );
NAND2xp33_ASAP7_75t_L g127 ( .A(n_54), .B(n_99), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_55), .B(n_145), .Y(n_233) );
BUFx10_ASAP7_75t_L g695 ( .A(n_56), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_57), .B(n_98), .Y(n_201) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_57), .Y(n_711) );
INVx2_ASAP7_75t_L g569 ( .A(n_58), .Y(n_569) );
NAND2xp33_ASAP7_75t_L g135 ( .A(n_59), .B(n_108), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_60), .B(n_147), .Y(n_200) );
INVx1_ASAP7_75t_L g665 ( .A(n_61), .Y(n_665) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_62), .Y(n_191) );
INVx2_ASAP7_75t_L g93 ( .A(n_63), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_64), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_65), .B(n_119), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g109 ( .A(n_66), .B(n_110), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_67), .Y(n_211) );
INVx1_ASAP7_75t_L g181 ( .A(n_68), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_69), .Y(n_162) );
AND2x2_ASAP7_75t_L g173 ( .A(n_70), .B(n_90), .Y(n_173) );
INVx1_ASAP7_75t_L g520 ( .A(n_71), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_71), .A2(n_561), .B(n_565), .Y(n_560) );
INVx2_ASAP7_75t_L g542 ( .A(n_72), .Y(n_542) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_73), .Y(n_490) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_74), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_75), .B(n_138), .Y(n_137) );
BUFx3_ASAP7_75t_L g487 ( .A(n_76), .Y(n_487) );
INVx1_ASAP7_75t_L g503 ( .A(n_76), .Y(n_503) );
BUFx3_ASAP7_75t_L g488 ( .A(n_77), .Y(n_488) );
INVx1_ASAP7_75t_L g527 ( .A(n_77), .Y(n_527) );
AOI21xp33_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_466), .B(n_473), .Y(n_78) );
INVx3_ASAP7_75t_L g79 ( .A(n_80), .Y(n_79) );
AND2x4_ASAP7_75t_L g80 ( .A(n_81), .B(n_374), .Y(n_80) );
NOR4xp25_ASAP7_75t_L g81 ( .A(n_82), .B(n_271), .C(n_315), .D(n_334), .Y(n_81) );
NAND2xp5_ASAP7_75t_L g82 ( .A(n_83), .B(n_256), .Y(n_82) );
AOI222xp33_ASAP7_75t_L g83 ( .A1(n_84), .A2(n_152), .B1(n_193), .B2(n_222), .C1(n_237), .C2(n_246), .Y(n_83) );
AOI221xp5_ASAP7_75t_L g453 ( .A1(n_84), .A2(n_279), .B1(n_399), .B2(n_454), .C(n_456), .Y(n_453) );
AND2x2_ASAP7_75t_L g84 ( .A(n_85), .B(n_121), .Y(n_84) );
BUFx2_ASAP7_75t_L g390 ( .A(n_85), .Y(n_390) );
INVx2_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
AND2x4_ASAP7_75t_L g290 ( .A(n_86), .B(n_275), .Y(n_290) );
AND2x4_ASAP7_75t_L g368 ( .A(n_86), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g425 ( .A(n_86), .B(n_365), .Y(n_425) );
INVx2_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx2_ASAP7_75t_L g251 ( .A(n_88), .Y(n_251) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_88), .Y(n_371) );
OAI21x1_ASAP7_75t_L g88 ( .A1(n_89), .A2(n_94), .B(n_118), .Y(n_88) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_89), .A2(n_142), .B(n_151), .Y(n_141) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_89), .A2(n_209), .B(n_218), .Y(n_208) );
OAI21x1_ASAP7_75t_L g226 ( .A1(n_89), .A2(n_94), .B(n_118), .Y(n_226) );
OAI21x1_ASAP7_75t_L g255 ( .A1(n_89), .A2(n_142), .B(n_151), .Y(n_255) );
BUFx4f_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
OA21x2_ASAP7_75t_L g124 ( .A1(n_90), .A2(n_125), .B(n_137), .Y(n_124) );
INVx4_ASAP7_75t_L g156 ( .A(n_90), .Y(n_156) );
INVx3_ASAP7_75t_L g197 ( .A(n_90), .Y(n_197) );
OA21x2_ASAP7_75t_L g249 ( .A1(n_90), .A2(n_125), .B(n_137), .Y(n_249) );
OA21x2_ASAP7_75t_L g281 ( .A1(n_90), .A2(n_125), .B(n_137), .Y(n_281) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx2_ASAP7_75t_L g120 ( .A(n_91), .Y(n_120) );
INVx2_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g139 ( .A(n_92), .Y(n_139) );
OAI21x1_ASAP7_75t_L g94 ( .A1(n_95), .A2(n_104), .B(n_114), .Y(n_94) );
O2A1O1Ixp33_ASAP7_75t_L g95 ( .A1(n_96), .A2(n_97), .B(n_101), .C(n_103), .Y(n_95) );
INVx1_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_98), .Y(n_472) );
INVx1_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
INVx2_ASAP7_75t_L g129 ( .A(n_99), .Y(n_129) );
INVx2_ASAP7_75t_L g213 ( .A(n_99), .Y(n_213) );
BUFx6f_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
BUFx6f_ASAP7_75t_L g102 ( .A(n_100), .Y(n_102) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_100), .Y(n_108) );
INVx2_ASAP7_75t_L g111 ( .A(n_100), .Y(n_111) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_100), .Y(n_170) );
INVx1_ASAP7_75t_L g185 ( .A(n_100), .Y(n_185) );
INVx5_ASAP7_75t_L g134 ( .A(n_102), .Y(n_134) );
BUFx12f_ASAP7_75t_L g113 ( .A(n_103), .Y(n_113) );
INVx5_ASAP7_75t_L g131 ( .A(n_103), .Y(n_131) );
INVx5_ASAP7_75t_L g136 ( .A(n_103), .Y(n_136) );
O2A1O1Ixp33_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_106), .B(n_109), .C(n_112), .Y(n_104) );
O2A1O1Ixp5_ASAP7_75t_L g148 ( .A1(n_106), .A2(n_112), .B(n_149), .C(n_150), .Y(n_148) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g145 ( .A(n_108), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_108), .B(n_160), .Y(n_159) );
INVx2_ASAP7_75t_SL g189 ( .A(n_108), .Y(n_189) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g147 ( .A(n_111), .Y(n_147) );
INVx2_ASAP7_75t_L g167 ( .A(n_111), .Y(n_167) );
O2A1O1Ixp5_ASAP7_75t_L g210 ( .A1(n_112), .A2(n_211), .B(n_212), .C(n_214), .Y(n_210) );
INVx3_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_113), .Y(n_172) );
BUFx2_ASAP7_75t_L g186 ( .A(n_113), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_113), .A2(n_233), .B(n_234), .Y(n_232) );
OAI21x1_ASAP7_75t_L g125 ( .A1(n_114), .A2(n_126), .B(n_132), .Y(n_125) );
OAI21x1_ASAP7_75t_L g142 ( .A1(n_114), .A2(n_143), .B(n_148), .Y(n_142) );
OAI21x1_ASAP7_75t_L g198 ( .A1(n_114), .A2(n_199), .B(n_202), .Y(n_198) );
OAI21xp5_ASAP7_75t_L g209 ( .A1(n_114), .A2(n_210), .B(n_215), .Y(n_209) );
INVx8_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_115), .A2(n_158), .B(n_164), .Y(n_157) );
NOR2xp67_ASAP7_75t_L g176 ( .A(n_115), .B(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g469 ( .A(n_115), .Y(n_469) );
INVx8_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g235 ( .A(n_116), .Y(n_235) );
INVx3_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g330 ( .A(n_121), .B(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVxp67_ASAP7_75t_SL g393 ( .A(n_122), .Y(n_393) );
NAND2x1p5_ASAP7_75t_L g122 ( .A(n_123), .B(n_140), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g341 ( .A(n_124), .B(n_253), .Y(n_341) );
AND2x2_ASAP7_75t_L g398 ( .A(n_124), .B(n_253), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_124), .B(n_306), .Y(n_407) );
AOI21xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_128), .B(n_130), .Y(n_126) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_130), .A2(n_144), .B(n_146), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_130), .A2(n_216), .B(n_217), .Y(n_215) );
CKINVDCx6p67_ASAP7_75t_R g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_SL g163 ( .A(n_131), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_135), .B(n_136), .Y(n_132) );
NOR2xp67_ASAP7_75t_L g161 ( .A(n_134), .B(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g205 ( .A(n_136), .Y(n_205) );
AOI21x1_ASAP7_75t_L g229 ( .A1(n_136), .A2(n_230), .B(n_231), .Y(n_229) );
BUFx5_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g223 ( .A(n_140), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_140), .B(n_251), .Y(n_294) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g282 ( .A(n_141), .B(n_259), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_147), .B(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_L g372 ( .A(n_154), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g417 ( .A(n_154), .B(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g154 ( .A(n_155), .B(n_174), .Y(n_154) );
AND2x2_ASAP7_75t_L g263 ( .A(n_155), .B(n_221), .Y(n_263) );
OR2x2_ASAP7_75t_L g270 ( .A(n_155), .B(n_195), .Y(n_270) );
AND2x2_ASAP7_75t_L g423 ( .A(n_155), .B(n_208), .Y(n_423) );
AO21x2_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_173), .Y(n_155) );
INVx3_ASAP7_75t_L g177 ( .A(n_156), .Y(n_177) );
AO21x2_ASAP7_75t_L g244 ( .A1(n_156), .A2(n_157), .B(n_173), .Y(n_244) );
OAI21xp5_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_161), .B(n_163), .Y(n_158) );
OAI21xp33_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_168), .B(n_172), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_166), .A2(n_664), .B1(n_665), .B2(n_666), .Y(n_663) );
INVx1_ASAP7_75t_L g666 ( .A(n_166), .Y(n_666) );
NOR2xp33_ASAP7_75t_SL g168 ( .A(n_169), .B(n_171), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_169), .B(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_172), .A2(n_200), .B(n_201), .Y(n_199) );
INVx1_ASAP7_75t_L g221 ( .A(n_174), .Y(n_221) );
AND2x2_ASAP7_75t_L g323 ( .A(n_174), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g402 ( .A(n_174), .Y(n_402) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g241 ( .A(n_175), .Y(n_241) );
AOI21x1_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_178), .B(n_192), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_179), .B(n_187), .Y(n_178) );
OAI21x1_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_182), .B(n_186), .Y(n_179) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_186), .B(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AOI221xp5_ASAP7_75t_L g335 ( .A1(n_193), .A2(n_336), .B1(n_338), .B2(n_342), .C(n_347), .Y(n_335) );
AND2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_219), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_194), .B(n_353), .Y(n_352) );
NAND2xp67_ASAP7_75t_L g389 ( .A(n_194), .B(n_263), .Y(n_389) );
AND2x4_ASAP7_75t_L g444 ( .A(n_194), .B(n_323), .Y(n_444) );
AND2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_207), .Y(n_194) );
INVx1_ASAP7_75t_L g245 ( .A(n_195), .Y(n_245) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_195), .Y(n_266) );
INVx1_ASAP7_75t_L g311 ( .A(n_195), .Y(n_311) );
INVx1_ASAP7_75t_L g360 ( .A(n_195), .Y(n_360) );
AND2x2_ASAP7_75t_L g401 ( .A(n_195), .B(n_402), .Y(n_401) );
OAI21x1_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_198), .B(n_206), .Y(n_195) );
OAI21xp5_ASAP7_75t_L g227 ( .A1(n_196), .A2(n_228), .B(n_236), .Y(n_227) );
OAI21x1_ASAP7_75t_L g261 ( .A1(n_196), .A2(n_228), .B(n_236), .Y(n_261) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_205), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_207), .B(n_244), .Y(n_301) );
OR2x2_ASAP7_75t_L g359 ( .A(n_207), .B(n_360), .Y(n_359) );
BUFx3_ASAP7_75t_L g448 ( .A(n_207), .Y(n_448) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g242 ( .A(n_208), .Y(n_242) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AOI22xp33_ASAP7_75t_SL g449 ( .A1(n_219), .A2(n_290), .B1(n_450), .B2(n_451), .Y(n_449) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g408 ( .A(n_220), .B(n_344), .Y(n_408) );
OR2x2_ASAP7_75t_L g452 ( .A(n_220), .B(n_270), .Y(n_452) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g256 ( .A1(n_222), .A2(n_257), .B1(n_262), .B2(n_267), .Y(n_256) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
OR2x2_ASAP7_75t_L g434 ( .A(n_223), .B(n_350), .Y(n_434) );
BUFx3_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g328 ( .A(n_225), .Y(n_328) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
INVx1_ASAP7_75t_L g306 ( .A(n_226), .Y(n_306) );
OR2x2_ASAP7_75t_L g319 ( .A(n_226), .B(n_260), .Y(n_319) );
AND2x2_ASAP7_75t_L g416 ( .A(n_226), .B(n_253), .Y(n_416) );
BUFx2_ASAP7_75t_L g351 ( .A(n_227), .Y(n_351) );
OAI21x1_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_232), .B(n_235), .Y(n_228) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_243), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_240), .B(n_242), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_240), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g269 ( .A(n_241), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_241), .B(n_242), .Y(n_297) );
INVxp67_ASAP7_75t_SL g354 ( .A(n_241), .Y(n_354) );
OR2x2_ASAP7_75t_L g265 ( .A(n_242), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g345 ( .A(n_242), .Y(n_345) );
AND2x2_ASAP7_75t_L g395 ( .A(n_242), .B(n_311), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_242), .B(n_346), .Y(n_420) );
OR2x2_ASAP7_75t_L g296 ( .A(n_243), .B(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
INVx1_ASAP7_75t_L g313 ( .A(n_244), .Y(n_313) );
INVx2_ASAP7_75t_SL g324 ( .A(n_244), .Y(n_324) );
INVx1_ASAP7_75t_L g380 ( .A(n_245), .Y(n_380) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_250), .Y(n_247) );
OR2x2_ASAP7_75t_L g432 ( .A(n_248), .B(n_307), .Y(n_432) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx2_ASAP7_75t_SL g278 ( .A(n_249), .Y(n_278) );
INVx1_ASAP7_75t_SL g289 ( .A(n_249), .Y(n_289) );
BUFx2_ASAP7_75t_L g438 ( .A(n_249), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_250), .B(n_443), .Y(n_442) );
NAND2x1_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
AND2x4_ASAP7_75t_SL g274 ( .A(n_251), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g331 ( .A(n_251), .Y(n_331) );
BUFx2_ASAP7_75t_L g339 ( .A(n_251), .Y(n_339) );
INVx1_ASAP7_75t_L g387 ( .A(n_252), .Y(n_387) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_253), .B(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g277 ( .A(n_253), .B(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g369 ( .A(n_254), .B(n_260), .Y(n_369) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g365 ( .A(n_255), .B(n_260), .Y(n_365) );
AND2x2_ASAP7_75t_L g314 ( .A(n_257), .B(n_281), .Y(n_314) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g370 ( .A(n_258), .B(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g275 ( .A(n_259), .Y(n_275) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AOI22xp5_ASAP7_75t_L g376 ( .A1(n_262), .A2(n_280), .B1(n_377), .B2(n_382), .Y(n_376) );
AND2x4_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx1_ASAP7_75t_L g332 ( .A(n_263), .Y(n_332) );
INVx1_ASAP7_75t_L g465 ( .A(n_263), .Y(n_465) );
INVx1_ASAP7_75t_L g411 ( .A(n_264), .Y(n_411) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OAI211xp5_ASAP7_75t_L g271 ( .A1(n_268), .A2(n_272), .B(n_283), .C(n_298), .Y(n_271) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx1_ASAP7_75t_L g429 ( .A(n_269), .Y(n_429) );
INVx2_ASAP7_75t_L g346 ( .A(n_270), .Y(n_346) );
INVxp67_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
AO21x1_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_276), .B(n_279), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_274), .B(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g337 ( .A(n_274), .Y(n_337) );
INVx1_ASAP7_75t_L g415 ( .A(n_275), .Y(n_415) );
BUFx2_ASAP7_75t_L g450 ( .A(n_275), .Y(n_450) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NOR2x1_ASAP7_75t_SL g327 ( .A(n_277), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_278), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g358 ( .A(n_278), .Y(n_358) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
OR2x6_ASAP7_75t_SL g318 ( .A(n_280), .B(n_319), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_280), .B(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g286 ( .A(n_281), .Y(n_286) );
INVx2_ASAP7_75t_L g307 ( .A(n_282), .Y(n_307) );
OAI31xp33_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_287), .A3(n_291), .B(n_295), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g447 ( .A(n_286), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NOR2x1p5_ASAP7_75t_L g412 ( .A(n_289), .B(n_367), .Y(n_412) );
INVx2_ASAP7_75t_L g381 ( .A(n_290), .Y(n_381) );
INVxp67_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g455 ( .A(n_297), .Y(n_455) );
AOI22xp33_ASAP7_75t_SL g298 ( .A1(n_299), .A2(n_302), .B1(n_308), .B2(n_314), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g439 ( .A(n_300), .B(n_310), .Y(n_439) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_303), .A2(n_348), .B(n_352), .Y(n_347) );
OR2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_307), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_304), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_SL g364 ( .A(n_305), .B(n_365), .Y(n_364) );
BUFx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx1_ASAP7_75t_L g333 ( .A(n_310), .Y(n_333) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
BUFx2_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g400 ( .A(n_313), .B(n_401), .Y(n_400) );
O2A1O1Ixp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_320), .B(n_325), .C(n_333), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVxp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_318), .B(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g457 ( .A(n_319), .B(n_358), .Y(n_457) );
OAI21xp5_ASAP7_75t_L g459 ( .A1(n_319), .A2(n_460), .B(n_462), .Y(n_459) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g379 ( .A(n_323), .B(n_380), .Y(n_379) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_324), .Y(n_363) );
AO21x1_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_329), .B(n_332), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_328), .A2(n_332), .B1(n_378), .B2(n_381), .Y(n_377) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OAI21xp5_ASAP7_75t_L g404 ( .A1(n_330), .A2(n_405), .B(n_408), .Y(n_404) );
AND2x2_ASAP7_75t_L g397 ( .A(n_331), .B(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_355), .Y(n_334) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g441 ( .A(n_341), .Y(n_441) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx3_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x4_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
AND2x4_ASAP7_75t_L g399 ( .A(n_345), .B(n_400), .Y(n_399) );
OR2x2_ASAP7_75t_L g464 ( .A(n_345), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g443 ( .A(n_351), .Y(n_443) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AOI32xp33_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_361), .A3(n_364), .B1(n_366), .B2(n_372), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx1_ASAP7_75t_L g384 ( .A(n_358), .Y(n_384) );
INVx1_ASAP7_75t_L g373 ( .A(n_359), .Y(n_373) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_362), .B(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI21xp33_ASAP7_75t_L g462 ( .A1(n_364), .A2(n_417), .B(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g437 ( .A(n_365), .B(n_438), .Y(n_437) );
NAND2xp33_ASAP7_75t_SL g366 ( .A(n_367), .B(n_370), .Y(n_366) );
INVx3_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NOR4xp75_ASAP7_75t_L g374 ( .A(n_375), .B(n_403), .C(n_445), .D(n_459), .Y(n_374) );
NAND3xp33_ASAP7_75t_L g375 ( .A(n_376), .B(n_385), .C(n_396), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g418 ( .A(n_380), .Y(n_418) );
A2O1A1Ixp33_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_388), .B(n_390), .C(n_391), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OAI21xp5_ASAP7_75t_L g391 ( .A1(n_390), .A2(n_392), .B(n_394), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g430 ( .A(n_395), .Y(n_430) );
NAND2x1_ASAP7_75t_L g396 ( .A(n_397), .B(n_399), .Y(n_396) );
AND2x4_ASAP7_75t_L g422 ( .A(n_401), .B(n_423), .Y(n_422) );
NAND4xp75_ASAP7_75t_L g403 ( .A(n_404), .B(n_409), .C(n_426), .D(n_435), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AOI211x1_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_412), .B(n_413), .C(n_419), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_410), .A2(n_427), .B1(n_431), .B2(n_433), .Y(n_426) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
NOR3xp33_ASAP7_75t_L g456 ( .A(n_411), .B(n_457), .C(n_458), .Y(n_456) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_417), .Y(n_413) );
AND2x4_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B(n_424), .Y(n_419) );
NOR2xp67_ASAP7_75t_L g461 ( .A(n_421), .B(n_438), .Y(n_461) );
INVx2_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_L g458 ( .A(n_429), .Y(n_458) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OA21x2_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_439), .B(n_440), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OAI21xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_442), .B(n_444), .Y(n_440) );
OAI21xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_449), .B(n_453), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVxp67_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_470), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVxp67_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
AO21x1_ASAP7_75t_L g713 ( .A1(n_471), .A2(n_714), .B(n_715), .Y(n_713) );
OAI221xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B1(n_652), .B2(n_657), .C(n_707), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_475), .A2(n_708), .B1(n_711), .B2(n_712), .Y(n_707) );
HB1xp67_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
AOI221x1_ASAP7_75t_SL g476 ( .A1(n_477), .A2(n_528), .B1(n_533), .B2(n_613), .C(n_615), .Y(n_476) );
NAND4xp25_ASAP7_75t_L g477 ( .A(n_478), .B(n_489), .C(n_504), .D(n_519), .Y(n_477) );
BUFx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx5_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x4_ASAP7_75t_L g480 ( .A(n_481), .B(n_485), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x6_ASAP7_75t_L g525 ( .A(n_482), .B(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x6_ASAP7_75t_L g517 ( .A(n_483), .B(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_484), .Y(n_493) );
INVx1_ASAP7_75t_L g500 ( .A(n_484), .Y(n_500) );
AND2x2_ASAP7_75t_L g620 ( .A(n_484), .B(n_530), .Y(n_620) );
INVx2_ASAP7_75t_L g643 ( .A(n_484), .Y(n_643) );
INVx2_ASAP7_75t_L g509 ( .A(n_485), .Y(n_509) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
INVx2_ASAP7_75t_L g495 ( .A(n_487), .Y(n_495) );
AND2x4_ASAP7_75t_L g526 ( .A(n_487), .B(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g496 ( .A(n_488), .Y(n_496) );
AND2x4_ASAP7_75t_L g502 ( .A(n_488), .B(n_503), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_491), .B1(n_497), .B2(n_498), .Y(n_489) );
AOI222xp33_ASAP7_75t_L g593 ( .A1(n_490), .A2(n_594), .B1(n_598), .B2(n_599), .C1(n_604), .C2(n_605), .Y(n_593) );
AND2x4_ASAP7_75t_L g491 ( .A(n_492), .B(n_494), .Y(n_491) );
AND2x4_ASAP7_75t_L g512 ( .A(n_492), .B(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx6_ASAP7_75t_L g523 ( .A(n_494), .Y(n_523) );
AND2x4_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
INVx1_ASAP7_75t_L g518 ( .A(n_495), .Y(n_518) );
INVx1_ASAP7_75t_L g515 ( .A(n_496), .Y(n_515) );
AND2x6_ASAP7_75t_L g498 ( .A(n_499), .B(n_501), .Y(n_498) );
AND2x4_ASAP7_75t_L g521 ( .A(n_499), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx6f_ASAP7_75t_L g638 ( .A(n_502), .Y(n_638) );
INVx2_ASAP7_75t_L g651 ( .A(n_502), .Y(n_651) );
INVx1_ASAP7_75t_L g626 ( .A(n_503), .Y(n_626) );
AOI222xp33_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_506), .B1(n_510), .B2(n_511), .C1(n_516), .C2(n_517), .Y(n_504) );
OAI21xp5_ASAP7_75t_SL g557 ( .A1(n_505), .A2(n_558), .B(n_560), .Y(n_557) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx3_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx4f_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g693 ( .A(n_515), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_521), .B1(n_524), .B2(n_525), .Y(n_519) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
BUFx3_ASAP7_75t_L g636 ( .A(n_526), .Y(n_636) );
INVx1_ASAP7_75t_L g627 ( .A(n_527), .Y(n_627) );
AND2x4_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x4_ASAP7_75t_L g642 ( .A(n_530), .B(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g614 ( .A(n_531), .Y(n_614) );
BUFx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g621 ( .A(n_532), .Y(n_621) );
NAND3xp33_ASAP7_75t_L g533 ( .A(n_534), .B(n_593), .C(n_606), .Y(n_533) );
NOR3xp33_ASAP7_75t_SL g534 ( .A(n_535), .B(n_546), .C(n_571), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OR2x6_ASAP7_75t_L g536 ( .A(n_537), .B(n_543), .Y(n_536) );
INVx1_ASAP7_75t_L g559 ( .A(n_537), .Y(n_559) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_541), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g551 ( .A(n_540), .Y(n_551) );
INVx2_ASAP7_75t_L g556 ( .A(n_540), .Y(n_556) );
AND2x2_ASAP7_75t_L g564 ( .A(n_540), .B(n_542), .Y(n_564) );
INVx1_ASAP7_75t_L g575 ( .A(n_540), .Y(n_575) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g549 ( .A(n_542), .Y(n_549) );
AND2x4_ASAP7_75t_L g555 ( .A(n_542), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g587 ( .A(n_542), .Y(n_587) );
INVx1_ASAP7_75t_L g576 ( .A(n_543), .Y(n_576) );
OR2x6_ASAP7_75t_L g577 ( .A(n_543), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g596 ( .A(n_543), .Y(n_596) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_548), .Y(n_581) );
AND2x2_ASAP7_75t_L g608 ( .A(n_548), .B(n_602), .Y(n_608) );
AND2x4_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
INVx1_ASAP7_75t_L g578 ( .A(n_549), .Y(n_578) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx3_ASAP7_75t_L g582 ( .A(n_553), .Y(n_582) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx3_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g612 ( .A(n_555), .Y(n_612) );
AND2x4_ASAP7_75t_L g586 ( .A(n_556), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx3_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x4_ASAP7_75t_L g605 ( .A(n_563), .B(n_602), .Y(n_605) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx3_ASAP7_75t_L g589 ( .A(n_564), .Y(n_589) );
INVx2_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NAND2x1p5_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g592 ( .A(n_569), .Y(n_592) );
NAND2x1p5_ASAP7_75t_L g572 ( .A(n_573), .B(n_576), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_583), .Y(n_579) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
BUFx3_ASAP7_75t_L g603 ( .A(n_586), .Y(n_603) );
INVx2_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_SL g597 ( .A(n_589), .Y(n_597) );
OR2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
OAI221xp5_ASAP7_75t_L g644 ( .A1(n_598), .A2(n_604), .B1(n_629), .B2(n_645), .C(n_647), .Y(n_644) );
AND2x4_ASAP7_75t_L g599 ( .A(n_600), .B(n_603), .Y(n_599) );
AND2x4_ASAP7_75t_L g610 ( .A(n_600), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .B1(n_609), .B2(n_610), .Y(n_606) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
BUFx8_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_622), .B1(n_639), .B2(n_644), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OR2x6_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_SL g689 ( .A(n_620), .Y(n_689) );
OAI221xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_628), .B1(n_629), .B2(n_633), .C(n_634), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_624), .Y(n_646) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
AND2x2_ASAP7_75t_L g632 ( .A(n_626), .B(n_627), .Y(n_632) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
BUFx3_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
BUFx3_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx4_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AND2x4_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
AND2x4_ASAP7_75t_L g699 ( .A(n_643), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
BUFx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_654), .B(n_656), .Y(n_685) );
INVx1_ASAP7_75t_SL g714 ( .A(n_654), .Y(n_714) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_682), .B1(n_703), .B2(n_704), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_658), .A2(n_703), .B1(n_709), .B2(n_710), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B1(n_668), .B2(n_669), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_662), .B1(n_663), .B2(n_667), .Y(n_660) );
INVx1_ASAP7_75t_L g667 ( .A(n_661), .Y(n_667) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
CKINVDCx14_ASAP7_75t_R g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_671), .B1(n_676), .B2(n_677), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .B1(n_674), .B2(n_675), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_672), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_673), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B1(n_680), .B2(n_681), .Y(n_677) );
INVx1_ASAP7_75t_L g681 ( .A(n_678), .Y(n_681) );
INVx1_ASAP7_75t_L g680 ( .A(n_679), .Y(n_680) );
BUFx12f_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g709 ( .A(n_683), .Y(n_709) );
CKINVDCx20_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
OR2x6_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
OR2x4_ASAP7_75t_L g706 ( .A(n_685), .B(n_687), .Y(n_706) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AOI31xp33_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_690), .A3(n_694), .B(n_696), .Y(n_687) );
BUFx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVxp67_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g702 ( .A(n_693), .Y(n_702) );
INVx6_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVxp67_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
INVx2_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
AND2x4_ASAP7_75t_L g698 ( .A(n_699), .B(n_702), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
BUFx6f_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g710 ( .A(n_705), .Y(n_710) );
INVx8_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
BUFx2_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
endmodule