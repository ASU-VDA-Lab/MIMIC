module fake_jpeg_4367_n_79 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_79);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_79;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

CKINVDCx16_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_1),
.B(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_17),
.B(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_21),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_25),
.Y(n_31)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_1),
.Y(n_22)
);

OR2x2_ASAP7_75t_SL g32 ( 
.A(n_22),
.B(n_3),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_24),
.A2(n_10),
.B1(n_13),
.B2(n_11),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_2),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_20),
.A2(n_12),
.B1(n_16),
.B2(n_15),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_26),
.A2(n_29),
.B1(n_19),
.B2(n_20),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_21),
.A2(n_12),
.B1(n_16),
.B2(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_22),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_32),
.B(n_22),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_33),
.A2(n_35),
.B1(n_38),
.B2(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_26),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_37),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_21),
.B1(n_18),
.B2(n_24),
.Y(n_35)
);

OR2x4_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_19),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_41),
.Y(n_47)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_25),
.B1(n_27),
.B2(n_18),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_25),
.C(n_24),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_22),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_45),
.B(n_48),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_23),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_50),
.A2(n_36),
.B1(n_40),
.B2(n_22),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_51),
.B(n_3),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_49),
.A2(n_34),
.B1(n_39),
.B2(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_57),
.Y(n_63)
);

AO21x1_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_58),
.B(n_59),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_24),
.Y(n_55)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_45),
.A2(n_10),
.B1(n_9),
.B2(n_5),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_50),
.C(n_43),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_60),
.B(n_63),
.Y(n_68)
);

NOR3xp33_ASAP7_75t_SL g65 ( 
.A(n_57),
.B(n_51),
.C(n_9),
.Y(n_65)
);

AOI322xp5_ASAP7_75t_SL g67 ( 
.A1(n_65),
.A2(n_9),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_4),
.Y(n_67)
);

FAx1_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_53),
.CI(n_56),
.CON(n_66),
.SN(n_66)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_67),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_69),
.Y(n_71)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_61),
.C(n_65),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_72),
.B(n_62),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_72),
.C(n_62),
.Y(n_76)
);

BUFx24_ASAP7_75t_SL g74 ( 
.A(n_71),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_74),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_70),
.C(n_75),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_5),
.B(n_6),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_7),
.B(n_8),
.Y(n_79)
);


endmodule