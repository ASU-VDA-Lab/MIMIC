module fake_ariane_1713_n_1722 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1722);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1722;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_1067;
wire n_968;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

BUFx3_ASAP7_75t_L g155 ( 
.A(n_153),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_98),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_118),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_57),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_116),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_42),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_68),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_91),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_4),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_79),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_111),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_114),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_41),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_80),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_151),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_11),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_147),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_121),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_136),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_70),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_10),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_75),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_1),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_102),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_144),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_56),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_24),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_41),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_105),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_103),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_52),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_122),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_17),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_89),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_11),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_152),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_109),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_9),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_27),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_17),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_74),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_127),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_2),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_44),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_87),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_4),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_146),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_140),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_131),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_22),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_7),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_86),
.Y(n_207)
);

BUFx8_ASAP7_75t_SL g208 ( 
.A(n_63),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_126),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_16),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_132),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_90),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_29),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_124),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g215 ( 
.A(n_128),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_16),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_123),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_45),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_39),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_88),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_76),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_49),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_48),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_154),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_48),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_5),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_62),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_65),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_141),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_36),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_29),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_50),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g233 ( 
.A(n_34),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_134),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_72),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_19),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_5),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_110),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_32),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_83),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_30),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_143),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_23),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_60),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_137),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_28),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_42),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_82),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_95),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_61),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_54),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_13),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_14),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_139),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_97),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_94),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_37),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_33),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_115),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_13),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_30),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_125),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_66),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_84),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_71),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_39),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_113),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_59),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_28),
.Y(n_269)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_101),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_107),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_120),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_99),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_104),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_0),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_64),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_53),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_25),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_100),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_149),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_138),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_26),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_77),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_27),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_50),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_21),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_22),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_26),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_12),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_23),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_73),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_32),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_43),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_145),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_78),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_150),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_7),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_112),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_24),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_58),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_0),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_33),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_47),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_37),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_1),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_208),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_194),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_159),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_161),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_159),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_175),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_226),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_181),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_216),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_266),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_175),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_177),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_177),
.B(n_2),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_167),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_155),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_216),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_282),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_L g323 ( 
.A(n_236),
.B(n_3),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_204),
.B(n_3),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_237),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_184),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_282),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_184),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_160),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_207),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_207),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_220),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_220),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_288),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_304),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_164),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_164),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_212),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_224),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_266),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_286),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_212),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_163),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_224),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_182),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_229),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_190),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_244),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_244),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_198),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_229),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_234),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_199),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_234),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_195),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_277),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_250),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_250),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_205),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_264),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_233),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_286),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_215),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_167),
.Y(n_364)
);

NAND2xp33_ASAP7_75t_R g365 ( 
.A(n_157),
.B(n_106),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_206),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_264),
.Y(n_367)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_215),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_210),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_213),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_170),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_279),
.B(n_6),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_267),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_267),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_195),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_219),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_271),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_271),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_218),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_222),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_215),
.Y(n_381)
);

OAI21x1_ASAP7_75t_L g382 ( 
.A1(n_355),
.A2(n_172),
.B(n_156),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_355),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_308),
.B(n_291),
.Y(n_384)
);

INVx6_ASAP7_75t_L g385 ( 
.A(n_320),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_375),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_375),
.Y(n_387)
);

INVx2_ASAP7_75t_SL g388 ( 
.A(n_308),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_310),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_310),
.Y(n_390)
);

BUFx8_ASAP7_75t_L g391 ( 
.A(n_379),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_311),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_311),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_316),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_316),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_317),
.B(n_291),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_317),
.B(n_218),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_326),
.B(n_225),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_326),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_328),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_328),
.Y(n_401)
);

NAND3xp33_ASAP7_75t_L g402 ( 
.A(n_318),
.B(n_178),
.C(n_170),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_320),
.B(n_300),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_330),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_330),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_331),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_331),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_332),
.B(n_225),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_332),
.B(n_300),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_333),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_333),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_339),
.B(n_236),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_339),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_344),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_344),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_346),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_346),
.B(n_195),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_351),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_351),
.B(n_268),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_352),
.B(n_178),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_352),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_354),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_354),
.B(n_195),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_357),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_357),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_358),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_358),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_360),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_360),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_319),
.B(n_268),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_367),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_324),
.B(n_372),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_367),
.B(n_296),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_314),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_373),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_373),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_374),
.B(n_296),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_374),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_377),
.Y(n_439)
);

BUFx10_ASAP7_75t_L g440 ( 
.A(n_377),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_378),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_378),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_379),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_364),
.B(n_368),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_338),
.B(n_195),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_329),
.Y(n_446)
);

OAI21x1_ASAP7_75t_L g447 ( 
.A1(n_323),
.A2(n_172),
.B(n_156),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_371),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_343),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_315),
.B(n_155),
.Y(n_450)
);

BUFx4f_ASAP7_75t_L g451 ( 
.A(n_446),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_399),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_446),
.B(n_338),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_399),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_L g455 ( 
.A1(n_402),
.A2(n_340),
.B1(n_341),
.B2(n_362),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_388),
.B(n_348),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_444),
.B(n_348),
.Y(n_457)
);

INVxp33_ASAP7_75t_L g458 ( 
.A(n_434),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_388),
.B(n_349),
.Y(n_459)
);

AO22x2_ASAP7_75t_L g460 ( 
.A1(n_402),
.A2(n_292),
.B1(n_201),
.B2(n_284),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_399),
.Y(n_461)
);

INVxp67_ASAP7_75t_SL g462 ( 
.A(n_391),
.Y(n_462)
);

NAND2xp33_ASAP7_75t_L g463 ( 
.A(n_446),
.B(n_270),
.Y(n_463)
);

NAND3xp33_ASAP7_75t_L g464 ( 
.A(n_446),
.B(n_347),
.C(n_345),
.Y(n_464)
);

NAND3xp33_ASAP7_75t_L g465 ( 
.A(n_446),
.B(n_430),
.C(n_402),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_448),
.B(n_183),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_432),
.A2(n_381),
.B1(n_363),
.B2(n_349),
.Y(n_467)
);

INVx5_ASAP7_75t_L g468 ( 
.A(n_399),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_388),
.B(n_350),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_446),
.B(n_353),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_440),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_399),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_446),
.B(n_449),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_399),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_444),
.B(n_359),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_399),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_399),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_446),
.B(n_366),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_449),
.B(n_369),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_446),
.B(n_449),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_449),
.B(n_370),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_446),
.B(n_376),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_399),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_399),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_445),
.B(n_380),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_445),
.B(n_321),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_400),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_400),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_440),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_440),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_448),
.B(n_361),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_400),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_400),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_388),
.B(n_322),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_440),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_400),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_389),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_440),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_400),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_400),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_448),
.B(n_327),
.Y(n_501)
);

INVx5_ASAP7_75t_L g502 ( 
.A(n_400),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_440),
.Y(n_503)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_391),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_443),
.B(n_448),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_430),
.B(n_356),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_432),
.A2(n_183),
.B1(n_188),
.B2(n_193),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_400),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_400),
.Y(n_509)
);

INVx8_ASAP7_75t_L g510 ( 
.A(n_417),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_421),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_393),
.B(n_259),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_443),
.B(n_306),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_443),
.B(n_309),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_393),
.B(n_273),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_443),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g517 ( 
.A(n_385),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_421),
.Y(n_518)
);

BUFx4f_ASAP7_75t_L g519 ( 
.A(n_421),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_393),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_412),
.B(n_420),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_412),
.B(n_420),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_393),
.B(n_158),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_385),
.Y(n_524)
);

AND2x6_ASAP7_75t_L g525 ( 
.A(n_417),
.B(n_423),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_393),
.B(n_162),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_421),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_434),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_450),
.B(n_313),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_421),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_393),
.B(n_165),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_385),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_391),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_385),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_401),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_421),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_421),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_421),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_421),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_421),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_385),
.B(n_307),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_391),
.A2(n_223),
.B1(n_257),
.B2(n_247),
.Y(n_542)
);

BUFx10_ASAP7_75t_L g543 ( 
.A(n_385),
.Y(n_543)
);

INVxp67_ASAP7_75t_SL g544 ( 
.A(n_391),
.Y(n_544)
);

BUFx10_ASAP7_75t_L g545 ( 
.A(n_385),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_438),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_391),
.A2(n_223),
.B1(n_257),
.B2(n_247),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_450),
.B(n_336),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_385),
.B(n_312),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_438),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_438),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_438),
.Y(n_552)
);

NAND3xp33_ASAP7_75t_L g553 ( 
.A(n_450),
.B(n_365),
.C(n_232),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_438),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_433),
.B(n_337),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_394),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_438),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_447),
.A2(n_258),
.B1(n_305),
.B2(n_302),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_397),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_433),
.B(n_342),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_438),
.Y(n_561)
);

NAND2xp33_ASAP7_75t_SL g562 ( 
.A(n_433),
.B(n_230),
.Y(n_562)
);

BUFx8_ASAP7_75t_SL g563 ( 
.A(n_420),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_412),
.B(n_233),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_438),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_394),
.B(n_166),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_438),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_438),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_401),
.Y(n_569)
);

INVx1_ASAP7_75t_SL g570 ( 
.A(n_397),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_397),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_397),
.B(n_188),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_401),
.B(n_231),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_394),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_394),
.Y(n_575)
);

INVxp67_ASAP7_75t_R g576 ( 
.A(n_447),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_382),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_403),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_437),
.B(n_246),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_390),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_394),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_437),
.B(n_252),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_398),
.B(n_325),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_398),
.B(n_193),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_394),
.B(n_168),
.Y(n_585)
);

AND2x6_ASAP7_75t_L g586 ( 
.A(n_417),
.B(n_200),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_437),
.B(n_253),
.Y(n_587)
);

AND2x6_ASAP7_75t_L g588 ( 
.A(n_417),
.B(n_200),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_428),
.B(n_169),
.Y(n_589)
);

INVx6_ASAP7_75t_L g590 ( 
.A(n_417),
.Y(n_590)
);

OR2x6_ASAP7_75t_L g591 ( 
.A(n_420),
.B(n_239),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_404),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_419),
.B(n_260),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_447),
.A2(n_243),
.B1(n_305),
.B2(n_258),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_428),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_390),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_428),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_479),
.B(n_428),
.Y(n_598)
);

INVxp67_ASAP7_75t_L g599 ( 
.A(n_491),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_460),
.A2(n_447),
.B1(n_416),
.B2(n_441),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_578),
.B(n_428),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_481),
.B(n_428),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_580),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_528),
.B(n_398),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_516),
.B(n_435),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_SL g606 ( 
.A(n_578),
.B(n_404),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_457),
.B(n_435),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_497),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_485),
.B(n_435),
.Y(n_609)
);

AND2x2_ASAP7_75t_SL g610 ( 
.A(n_504),
.B(n_384),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_535),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_556),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_475),
.B(n_435),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_569),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_456),
.B(n_435),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_592),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_521),
.B(n_398),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_573),
.B(n_404),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_459),
.B(n_405),
.Y(n_619)
);

CKINVDCx11_ASAP7_75t_R g620 ( 
.A(n_571),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_596),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_486),
.B(n_405),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_581),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_506),
.B(n_405),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_583),
.B(n_408),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_L g626 ( 
.A1(n_465),
.A2(n_407),
.B1(n_413),
.B2(n_439),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_581),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_490),
.B(n_407),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_595),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_469),
.B(n_407),
.Y(n_630)
);

NOR2xp67_ASAP7_75t_L g631 ( 
.A(n_464),
.B(n_419),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_570),
.B(n_413),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_460),
.A2(n_416),
.B1(n_441),
.B2(n_392),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g634 ( 
.A(n_491),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_595),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_559),
.B(n_413),
.Y(n_636)
);

INVxp67_ASAP7_75t_L g637 ( 
.A(n_501),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_559),
.B(n_418),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_563),
.Y(n_639)
);

BUFx6f_ASAP7_75t_SL g640 ( 
.A(n_572),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_458),
.B(n_408),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_553),
.B(n_418),
.Y(n_642)
);

OR2x2_ASAP7_75t_L g643 ( 
.A(n_583),
.B(n_408),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_505),
.B(n_418),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_556),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_575),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_490),
.B(n_424),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_505),
.B(n_424),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_574),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_525),
.A2(n_564),
.B1(n_453),
.B2(n_501),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_521),
.B(n_424),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_503),
.B(n_425),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_555),
.B(n_408),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_563),
.Y(n_654)
);

BUFx5_ASAP7_75t_L g655 ( 
.A(n_543),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_494),
.B(n_425),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_533),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_574),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_522),
.B(n_564),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_510),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_590),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_575),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_529),
.B(n_427),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_466),
.B(n_427),
.Y(n_664)
);

NOR3xp33_ASAP7_75t_L g665 ( 
.A(n_560),
.B(n_176),
.C(n_384),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_590),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_471),
.B(n_431),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_466),
.B(n_431),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_451),
.A2(n_396),
.B(n_384),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_466),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_590),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_590),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_575),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_597),
.B(n_431),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_597),
.B(n_436),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_597),
.B(n_436),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_572),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_454),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_510),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_454),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_520),
.B(n_436),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_548),
.B(n_412),
.Y(n_682)
);

NOR3xp33_ASAP7_75t_L g683 ( 
.A(n_579),
.B(n_409),
.C(n_396),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_471),
.B(n_439),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_510),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_582),
.B(n_442),
.Y(n_686)
);

BUFx5_ASAP7_75t_L g687 ( 
.A(n_543),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_471),
.B(n_442),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_510),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_489),
.B(n_396),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_461),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_461),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_525),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_572),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_525),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_571),
.B(n_403),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_587),
.B(n_409),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_474),
.Y(n_698)
);

INVxp67_ASAP7_75t_SL g699 ( 
.A(n_489),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_520),
.B(n_390),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_593),
.B(n_409),
.Y(n_701)
);

NAND3xp33_ASAP7_75t_L g702 ( 
.A(n_455),
.B(n_395),
.C(n_392),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_520),
.B(n_392),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_474),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_591),
.B(n_417),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_525),
.Y(n_706)
);

AO221x1_ASAP7_75t_L g707 ( 
.A1(n_460),
.A2(n_230),
.B1(n_301),
.B2(n_261),
.C(n_302),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_591),
.B(n_417),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_525),
.B(n_512),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_525),
.B(n_392),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_584),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_514),
.B(n_395),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_584),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_515),
.B(n_395),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_SL g715 ( 
.A(n_504),
.B(n_395),
.Y(n_715)
);

INVx5_ASAP7_75t_L g716 ( 
.A(n_543),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_584),
.Y(n_717)
);

O2A1O1Ixp5_ASAP7_75t_L g718 ( 
.A1(n_473),
.A2(n_441),
.B(n_429),
.C(n_426),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_591),
.B(n_462),
.Y(n_719)
);

OR2x6_ASAP7_75t_L g720 ( 
.A(n_591),
.B(n_423),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_483),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_541),
.B(n_406),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_549),
.B(n_406),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_451),
.B(n_406),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_489),
.B(n_406),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_483),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_586),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_L g728 ( 
.A1(n_495),
.A2(n_441),
.B1(n_429),
.B2(n_426),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_487),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_495),
.B(n_498),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_495),
.B(n_410),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_524),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_498),
.B(n_410),
.Y(n_733)
);

OAI22xp33_ASAP7_75t_L g734 ( 
.A1(n_533),
.A2(n_544),
.B1(n_576),
.B2(n_239),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_498),
.B(n_410),
.Y(n_735)
);

INVx1_ASAP7_75t_SL g736 ( 
.A(n_513),
.Y(n_736)
);

NOR3xp33_ASAP7_75t_L g737 ( 
.A(n_470),
.B(n_285),
.C(n_299),
.Y(n_737)
);

OR2x2_ASAP7_75t_L g738 ( 
.A(n_467),
.B(n_334),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_451),
.B(n_410),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_478),
.B(n_411),
.Y(n_740)
);

INVx8_ASAP7_75t_L g741 ( 
.A(n_586),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_500),
.B(n_411),
.Y(n_742)
);

INVxp67_ASAP7_75t_L g743 ( 
.A(n_562),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_487),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_460),
.B(n_507),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_482),
.B(n_411),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_523),
.B(n_411),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_586),
.Y(n_748)
);

AND2x6_ASAP7_75t_L g749 ( 
.A(n_577),
.B(n_423),
.Y(n_749)
);

AO22x2_ASAP7_75t_L g750 ( 
.A1(n_542),
.A2(n_289),
.B1(n_287),
.B2(n_297),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_586),
.B(n_414),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_500),
.B(n_414),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_493),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_493),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_586),
.B(n_414),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_SL g756 ( 
.A(n_586),
.B(n_335),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_588),
.B(n_414),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_526),
.B(n_415),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_588),
.B(n_415),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_588),
.B(n_547),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_531),
.B(n_415),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_566),
.B(n_415),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_623),
.Y(n_763)
);

NAND3xp33_ASAP7_75t_SL g764 ( 
.A(n_737),
.B(n_622),
.C(n_601),
.Y(n_764)
);

BUFx2_ASAP7_75t_L g765 ( 
.A(n_604),
.Y(n_765)
);

NOR3xp33_ASAP7_75t_L g766 ( 
.A(n_659),
.B(n_243),
.C(n_241),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_624),
.B(n_588),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_660),
.B(n_480),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_730),
.A2(n_519),
.B(n_463),
.Y(n_769)
);

O2A1O1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_601),
.A2(n_624),
.B(n_637),
.C(n_622),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_660),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_660),
.B(n_585),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_720),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_603),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_607),
.B(n_588),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_607),
.B(n_588),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_599),
.B(n_589),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_632),
.B(n_594),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_618),
.A2(n_558),
.B1(n_576),
.B2(n_577),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_632),
.B(n_416),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_750),
.A2(n_429),
.B1(n_416),
.B2(n_422),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_660),
.Y(n_782)
);

AOI21x1_ASAP7_75t_L g783 ( 
.A1(n_724),
.A2(n_472),
.B(n_452),
.Y(n_783)
);

NAND2xp33_ASAP7_75t_L g784 ( 
.A(n_655),
.B(n_500),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_L g785 ( 
.A1(n_699),
.A2(n_577),
.B1(n_509),
.B2(n_537),
.Y(n_785)
);

AOI21x1_ASAP7_75t_L g786 ( 
.A1(n_724),
.A2(n_472),
.B(n_452),
.Y(n_786)
);

O2A1O1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_637),
.A2(n_429),
.B(n_426),
.C(n_422),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_599),
.B(n_509),
.Y(n_788)
);

O2A1O1Ixp33_ASAP7_75t_SL g789 ( 
.A1(n_628),
.A2(n_538),
.B(n_568),
.C(n_567),
.Y(n_789)
);

BUFx4f_ASAP7_75t_L g790 ( 
.A(n_719),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_619),
.B(n_422),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_716),
.A2(n_519),
.B(n_463),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_634),
.B(n_509),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_634),
.B(n_537),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_719),
.B(n_500),
.Y(n_795)
);

INVxp67_ASAP7_75t_L g796 ( 
.A(n_641),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_716),
.A2(n_519),
.B(n_517),
.Y(n_797)
);

BUFx8_ASAP7_75t_L g798 ( 
.A(n_640),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_716),
.A2(n_517),
.B(n_477),
.Y(n_799)
);

OAI21xp33_ASAP7_75t_L g800 ( 
.A1(n_619),
.A2(n_278),
.B(n_275),
.Y(n_800)
);

BUFx2_ASAP7_75t_L g801 ( 
.A(n_625),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_696),
.B(n_617),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_650),
.A2(n_562),
.B1(n_568),
.B2(n_567),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_627),
.Y(n_804)
);

O2A1O1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_651),
.A2(n_422),
.B(n_426),
.C(n_269),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_716),
.A2(n_699),
.B(n_602),
.Y(n_806)
);

NOR3xp33_ASAP7_75t_L g807 ( 
.A(n_606),
.B(n_261),
.C(n_241),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_741),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_697),
.B(n_423),
.Y(n_809)
);

NOR2x1_ASAP7_75t_L g810 ( 
.A(n_643),
.B(n_537),
.Y(n_810)
);

OAI321xp33_ASAP7_75t_L g811 ( 
.A1(n_734),
.A2(n_289),
.A3(n_297),
.B1(n_230),
.B2(n_387),
.C(n_383),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_697),
.B(n_701),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_701),
.B(n_546),
.Y(n_813)
);

BUFx12f_ASAP7_75t_L g814 ( 
.A(n_620),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_598),
.A2(n_477),
.B(n_476),
.Y(n_815)
);

INVx1_ASAP7_75t_SL g816 ( 
.A(n_653),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_679),
.B(n_500),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_677),
.B(n_423),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_629),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_628),
.A2(n_731),
.B(n_725),
.Y(n_820)
);

O2A1O1Ixp33_ASAP7_75t_SL g821 ( 
.A1(n_613),
.A2(n_508),
.B(n_476),
.C(n_484),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_661),
.B(n_546),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_693),
.B(n_561),
.Y(n_823)
);

OAI21xp5_ASAP7_75t_L g824 ( 
.A1(n_718),
.A2(n_488),
.B(n_484),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_656),
.B(n_423),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_683),
.B(n_546),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_711),
.B(n_233),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_735),
.A2(n_508),
.B(n_496),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_635),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_690),
.A2(n_703),
.B(n_700),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_741),
.Y(n_831)
);

BUFx2_ASAP7_75t_L g832 ( 
.A(n_657),
.Y(n_832)
);

AOI21x1_ASAP7_75t_L g833 ( 
.A1(n_739),
.A2(n_496),
.B(n_538),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_683),
.B(n_552),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_741),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_732),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_694),
.B(n_290),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_713),
.B(n_293),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_667),
.A2(n_492),
.B(n_488),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_670),
.B(n_552),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_610),
.A2(n_492),
.B1(n_550),
.B2(n_551),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_621),
.Y(n_842)
);

A2O1A1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_663),
.A2(n_552),
.B(n_527),
.C(n_499),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_684),
.A2(n_550),
.B(n_551),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_666),
.B(n_554),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_644),
.A2(n_577),
.B1(n_554),
.B2(n_557),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_750),
.A2(n_215),
.B1(n_189),
.B2(n_227),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_685),
.B(n_561),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_615),
.B(n_557),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_682),
.B(n_303),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_608),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_671),
.B(n_577),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_615),
.B(n_499),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_722),
.B(n_511),
.Y(n_854)
);

A2O1A1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_663),
.A2(n_536),
.B(n_511),
.C(n_540),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_732),
.Y(n_856)
);

NOR2xp67_ASAP7_75t_L g857 ( 
.A(n_702),
.B(n_386),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_732),
.Y(n_858)
);

OAI21xp33_ASAP7_75t_L g859 ( 
.A1(n_630),
.A2(n_230),
.B(n_518),
.Y(n_859)
);

NOR3xp33_ASAP7_75t_L g860 ( 
.A(n_737),
.B(n_540),
.C(n_518),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_722),
.B(n_527),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_718),
.A2(n_669),
.B(n_747),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_686),
.A2(n_539),
.B(n_536),
.C(n_530),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_717),
.B(n_530),
.Y(n_864)
);

O2A1O1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_648),
.A2(n_638),
.B(n_636),
.C(n_642),
.Y(n_865)
);

AOI21x1_ASAP7_75t_L g866 ( 
.A1(n_733),
.A2(n_539),
.B(n_382),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_686),
.B(n_524),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_611),
.B(n_532),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_614),
.B(n_532),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_672),
.B(n_534),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_705),
.B(n_386),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_688),
.A2(n_565),
.B(n_561),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_610),
.A2(n_534),
.B1(n_565),
.B2(n_561),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_734),
.A2(n_565),
.B1(n_561),
.B2(n_191),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_689),
.B(n_565),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_616),
.B(n_565),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_695),
.A2(n_187),
.B1(n_171),
.B2(n_173),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_646),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_720),
.Y(n_879)
);

INVx4_ASAP7_75t_L g880 ( 
.A(n_720),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_712),
.B(n_468),
.Y(n_881)
);

OR2x6_ASAP7_75t_L g882 ( 
.A(n_639),
.B(n_382),
.Y(n_882)
);

A2O1A1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_712),
.A2(n_382),
.B(n_263),
.C(n_221),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_706),
.B(n_545),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_705),
.B(n_545),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_708),
.B(n_386),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_681),
.A2(n_502),
.B(n_468),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_647),
.A2(n_502),
.B(n_468),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_652),
.A2(n_502),
.B(n_468),
.Y(n_889)
);

OR2x6_ASAP7_75t_L g890 ( 
.A(n_654),
.B(n_189),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_678),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_708),
.B(n_468),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_745),
.B(n_502),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_662),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_714),
.A2(n_502),
.B(n_545),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_665),
.B(n_386),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_680),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_673),
.Y(n_898)
);

A2O1A1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_709),
.A2(n_263),
.B(n_209),
.C(n_214),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_631),
.B(n_174),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_736),
.B(n_640),
.Y(n_901)
);

O2A1O1Ixp5_ASAP7_75t_L g902 ( 
.A1(n_609),
.A2(n_386),
.B(n_387),
.C(n_383),
.Y(n_902)
);

AOI33xp33_ASAP7_75t_L g903 ( 
.A1(n_633),
.A2(n_387),
.A3(n_383),
.B1(n_221),
.B2(n_214),
.B3(n_209),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_674),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_747),
.A2(n_179),
.B(n_180),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_664),
.B(n_386),
.Y(n_906)
);

INVx1_ASAP7_75t_SL g907 ( 
.A(n_738),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_691),
.Y(n_908)
);

OAI21xp33_ASAP7_75t_L g909 ( 
.A1(n_675),
.A2(n_230),
.B(n_295),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_758),
.A2(n_249),
.B(n_186),
.Y(n_910)
);

NOR3xp33_ASAP7_75t_L g911 ( 
.A(n_665),
.B(n_203),
.C(n_295),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_676),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_645),
.Y(n_913)
);

AOI21x1_ASAP7_75t_L g914 ( 
.A1(n_742),
.A2(n_203),
.B(n_270),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_750),
.B(n_227),
.Y(n_915)
);

INVxp67_ASAP7_75t_L g916 ( 
.A(n_756),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_668),
.B(n_185),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_758),
.A2(n_254),
.B(n_196),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_761),
.A2(n_255),
.B(n_197),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_761),
.A2(n_256),
.B(n_211),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_762),
.A2(n_262),
.B(n_228),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_762),
.A2(n_265),
.B(n_235),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_723),
.A2(n_192),
.B(n_240),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_760),
.A2(n_274),
.B1(n_238),
.B2(n_283),
.Y(n_924)
);

INVxp33_ASAP7_75t_L g925 ( 
.A(n_633),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_710),
.B(n_242),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_692),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_612),
.B(n_655),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_740),
.A2(n_276),
.B(n_245),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_612),
.B(n_248),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_605),
.A2(n_281),
.B(n_280),
.Y(n_931)
);

BUFx4f_ASAP7_75t_L g932 ( 
.A(n_749),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_732),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_748),
.B(n_298),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_649),
.A2(n_272),
.B1(n_251),
.B2(n_294),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_740),
.A2(n_270),
.B(n_294),
.Y(n_936)
);

OAI21xp33_ASAP7_75t_L g937 ( 
.A1(n_658),
.A2(n_294),
.B(n_217),
.Y(n_937)
);

INVxp67_ASAP7_75t_L g938 ( 
.A(n_749),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_655),
.B(n_270),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_760),
.B(n_743),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_743),
.B(n_6),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_742),
.A2(n_294),
.B(n_217),
.Y(n_942)
);

NOR2xp67_ASAP7_75t_SL g943 ( 
.A(n_814),
.B(n_832),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_812),
.B(n_749),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_770),
.B(n_749),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_796),
.B(n_749),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_796),
.B(n_727),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_SL g948 ( 
.A(n_790),
.B(n_727),
.Y(n_948)
);

AO32x1_ASAP7_75t_L g949 ( 
.A1(n_846),
.A2(n_626),
.A3(n_728),
.B1(n_753),
.B2(n_744),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_802),
.B(n_600),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_778),
.A2(n_600),
.B1(n_757),
.B2(n_755),
.Y(n_951)
);

O2A1O1Ixp33_ASAP7_75t_SL g952 ( 
.A1(n_764),
.A2(n_752),
.B(n_759),
.C(n_751),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_774),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_784),
.A2(n_687),
.B(n_655),
.Y(n_954)
);

INVx4_ASAP7_75t_L g955 ( 
.A(n_790),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_771),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_932),
.B(n_715),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_932),
.B(n_655),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_798),
.Y(n_959)
);

INVx1_ASAP7_75t_SL g960 ( 
.A(n_765),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_851),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_835),
.Y(n_962)
);

HB1xp67_ASAP7_75t_L g963 ( 
.A(n_801),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_835),
.Y(n_964)
);

CKINVDCx16_ASAP7_75t_R g965 ( 
.A(n_890),
.Y(n_965)
);

NAND3xp33_ASAP7_75t_L g966 ( 
.A(n_807),
.B(n_746),
.C(n_752),
.Y(n_966)
);

OAI21xp33_ASAP7_75t_L g967 ( 
.A1(n_800),
.A2(n_746),
.B(n_726),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_825),
.A2(n_754),
.B1(n_729),
.B2(n_721),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_880),
.B(n_655),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_798),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_816),
.B(n_707),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_779),
.A2(n_861),
.B(n_854),
.Y(n_972)
);

AO32x1_ASAP7_75t_L g973 ( 
.A1(n_896),
.A2(n_704),
.A3(n_698),
.B1(n_12),
.B2(n_14),
.Y(n_973)
);

O2A1O1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_764),
.A2(n_8),
.B(n_10),
.C(n_15),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_880),
.B(n_18),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_850),
.B(n_18),
.Y(n_976)
);

NAND3xp33_ASAP7_75t_L g977 ( 
.A(n_807),
.B(n_202),
.C(n_217),
.Y(n_977)
);

NAND2xp33_ASAP7_75t_SL g978 ( 
.A(n_835),
.B(n_687),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_806),
.A2(n_687),
.B(n_294),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_766),
.B(n_687),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_791),
.A2(n_687),
.B(n_217),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_766),
.B(n_687),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_771),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_925),
.B(n_19),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_879),
.B(n_20),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_777),
.A2(n_217),
.B(n_202),
.C(n_270),
.Y(n_986)
);

OR2x6_ASAP7_75t_L g987 ( 
.A(n_940),
.B(n_202),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_780),
.A2(n_202),
.B1(n_21),
.B2(n_25),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_SL g989 ( 
.A(n_938),
.B(n_202),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_904),
.B(n_270),
.Y(n_990)
);

CKINVDCx6p67_ASAP7_75t_R g991 ( 
.A(n_890),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_777),
.A2(n_270),
.B(n_31),
.C(n_34),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_767),
.A2(n_20),
.B1(n_31),
.B2(n_35),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_771),
.B(n_270),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_SL g995 ( 
.A(n_938),
.B(n_35),
.Y(n_995)
);

INVx1_ASAP7_75t_SL g996 ( 
.A(n_907),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_763),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_912),
.B(n_38),
.Y(n_998)
);

NAND2x1p5_ASAP7_75t_L g999 ( 
.A(n_835),
.B(n_81),
.Y(n_999)
);

AOI21xp33_ASAP7_75t_L g1000 ( 
.A1(n_847),
.A2(n_38),
.B(n_40),
.Y(n_1000)
);

A2O1A1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_813),
.A2(n_40),
.B(n_43),
.C(n_44),
.Y(n_1001)
);

BUFx4f_ASAP7_75t_L g1002 ( 
.A(n_890),
.Y(n_1002)
);

BUFx12f_ASAP7_75t_L g1003 ( 
.A(n_827),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_849),
.A2(n_853),
.B(n_776),
.Y(n_1004)
);

OR2x6_ASAP7_75t_L g1005 ( 
.A(n_773),
.B(n_901),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_871),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_775),
.A2(n_96),
.B(n_142),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_901),
.Y(n_1008)
);

NAND2x1p5_ASAP7_75t_L g1009 ( 
.A(n_808),
.B(n_93),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_804),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_771),
.B(n_46),
.Y(n_1011)
);

O2A1O1Ixp5_ASAP7_75t_L g1012 ( 
.A1(n_862),
.A2(n_49),
.B(n_51),
.C(n_55),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_809),
.B(n_51),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_773),
.B(n_67),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_813),
.B(n_69),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_819),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_810),
.B(n_85),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_865),
.A2(n_92),
.B(n_117),
.C(n_119),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_837),
.B(n_148),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_829),
.Y(n_1020)
);

OAI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_830),
.A2(n_129),
.B(n_130),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_866),
.A2(n_133),
.B(n_135),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_911),
.A2(n_941),
.B(n_794),
.C(n_793),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_878),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_894),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_911),
.A2(n_788),
.B(n_794),
.C(n_793),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_916),
.B(n_818),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_916),
.B(n_886),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_782),
.B(n_924),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_915),
.B(n_788),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_795),
.B(n_808),
.Y(n_1031)
);

BUFx2_ASAP7_75t_L g1032 ( 
.A(n_882),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_882),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_831),
.B(n_782),
.Y(n_1034)
);

BUFx2_ASAP7_75t_L g1035 ( 
.A(n_882),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_842),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_891),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_847),
.B(n_838),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_820),
.A2(n_939),
.B(n_785),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_934),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_782),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_913),
.B(n_898),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_782),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_892),
.B(n_874),
.Y(n_1044)
);

CKINVDCx11_ASAP7_75t_R g1045 ( 
.A(n_836),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_SL g1046 ( 
.A(n_936),
.B(n_831),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_897),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_R g1048 ( 
.A(n_856),
.B(n_858),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_939),
.A2(n_852),
.B(n_769),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_917),
.B(n_929),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_781),
.B(n_903),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_900),
.B(n_856),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_858),
.B(n_933),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_836),
.Y(n_1054)
);

AO32x2_ASAP7_75t_L g1055 ( 
.A1(n_935),
.A2(n_883),
.A3(n_811),
.B1(n_781),
.B2(n_821),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_852),
.A2(n_815),
.B(n_895),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_905),
.B(n_910),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_933),
.B(n_826),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_792),
.A2(n_828),
.B(n_772),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_867),
.A2(n_887),
.B(n_881),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_836),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_836),
.B(n_877),
.Y(n_1062)
);

AOI21x1_ASAP7_75t_L g1063 ( 
.A1(n_914),
.A2(n_783),
.B(n_786),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_841),
.A2(n_876),
.B1(n_834),
.B2(n_873),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_787),
.A2(n_805),
.B(n_845),
.C(n_860),
.Y(n_1065)
);

AOI21x1_ASAP7_75t_L g1066 ( 
.A1(n_833),
.A2(n_857),
.B(n_893),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_855),
.A2(n_863),
.B(n_843),
.Y(n_1067)
);

AOI33xp33_ASAP7_75t_L g1068 ( 
.A1(n_789),
.A2(n_803),
.A3(n_934),
.B1(n_927),
.B2(n_908),
.B3(n_860),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_868),
.A2(n_869),
.B1(n_864),
.B2(n_845),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_906),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_930),
.B(n_823),
.Y(n_1071)
);

INVx4_ASAP7_75t_L g1072 ( 
.A(n_885),
.Y(n_1072)
);

AOI21x1_ASAP7_75t_L g1073 ( 
.A1(n_823),
.A2(n_942),
.B(n_768),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_840),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_822),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_926),
.B(n_921),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_918),
.A2(n_920),
.B(n_919),
.C(n_922),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_928),
.A2(n_824),
.B(n_844),
.Y(n_1078)
);

AOI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_870),
.A2(n_822),
.B1(n_875),
.B2(n_817),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_870),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_848),
.Y(n_1081)
);

CKINVDCx8_ASAP7_75t_R g1082 ( 
.A(n_899),
.Y(n_1082)
);

AND2x4_ASAP7_75t_SL g1083 ( 
.A(n_902),
.B(n_872),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_839),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_902),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_923),
.B(n_931),
.Y(n_1086)
);

OR2x2_ASAP7_75t_L g1087 ( 
.A(n_960),
.B(n_909),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_954),
.A2(n_799),
.B(n_797),
.Y(n_1088)
);

AOI21x1_ASAP7_75t_L g1089 ( 
.A1(n_1049),
.A2(n_884),
.B(n_888),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_1045),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_960),
.B(n_859),
.Y(n_1091)
);

AO31x2_ASAP7_75t_L g1092 ( 
.A1(n_1060),
.A2(n_889),
.A3(n_937),
.B(n_972),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_1059),
.A2(n_1056),
.B(n_1039),
.Y(n_1093)
);

NAND3xp33_ASAP7_75t_SL g1094 ( 
.A(n_974),
.B(n_995),
.C(n_992),
.Y(n_1094)
);

O2A1O1Ixp33_ASAP7_75t_SL g1095 ( 
.A1(n_1026),
.A2(n_1023),
.B(n_1050),
.C(n_945),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_955),
.Y(n_1096)
);

O2A1O1Ixp5_ASAP7_75t_L g1097 ( 
.A1(n_1086),
.A2(n_1076),
.B(n_1021),
.C(n_1067),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1015),
.A2(n_1004),
.B(n_979),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_981),
.A2(n_1057),
.B(n_980),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1065),
.A2(n_945),
.B(n_966),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_1064),
.A2(n_944),
.B(n_1013),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_982),
.A2(n_1064),
.B(n_1021),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_997),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_965),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_955),
.B(n_1005),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_1063),
.A2(n_1078),
.B(n_1073),
.Y(n_1106)
);

NOR2xp67_ASAP7_75t_L g1107 ( 
.A(n_1008),
.B(n_1003),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_989),
.A2(n_949),
.B(n_952),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_989),
.A2(n_949),
.B(n_1069),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1030),
.A2(n_984),
.B1(n_998),
.B2(n_988),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_1066),
.A2(n_1022),
.B(n_968),
.Y(n_1111)
);

AO31x2_ASAP7_75t_L g1112 ( 
.A1(n_951),
.A2(n_968),
.A3(n_1069),
.B(n_986),
.Y(n_1112)
);

BUFx4f_ASAP7_75t_L g1113 ( 
.A(n_991),
.Y(n_1113)
);

AOI221x1_ASAP7_75t_L g1114 ( 
.A1(n_1000),
.A2(n_988),
.B1(n_993),
.B2(n_1001),
.C(n_1018),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1010),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_SL g1116 ( 
.A(n_1002),
.B(n_995),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_963),
.B(n_985),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1016),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1070),
.B(n_1080),
.Y(n_1119)
);

AO21x2_ASAP7_75t_L g1120 ( 
.A1(n_951),
.A2(n_990),
.B(n_1044),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_1007),
.A2(n_1084),
.B(n_990),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1046),
.A2(n_1077),
.B(n_958),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_1071),
.A2(n_1019),
.B(n_1068),
.C(n_1038),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1085),
.A2(n_1058),
.B(n_1012),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1075),
.A2(n_993),
.B1(n_976),
.B2(n_1020),
.Y(n_1125)
);

OR2x6_ASAP7_75t_L g1126 ( 
.A(n_1005),
.B(n_1040),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1009),
.A2(n_969),
.B(n_1080),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_950),
.A2(n_1006),
.B1(n_946),
.B2(n_947),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_1054),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_1009),
.A2(n_994),
.B(n_999),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1024),
.Y(n_1131)
);

O2A1O1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_975),
.A2(n_1011),
.B(n_957),
.C(n_1028),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_1048),
.Y(n_1133)
);

AO21x2_ASAP7_75t_L g1134 ( 
.A1(n_1062),
.A2(n_967),
.B(n_1029),
.Y(n_1134)
);

A2O1A1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_1052),
.A2(n_1017),
.B(n_1042),
.C(n_1014),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1025),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_L g1137 ( 
.A1(n_1002),
.A2(n_971),
.B1(n_1047),
.B2(n_1036),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_985),
.B(n_1027),
.Y(n_1138)
);

NAND3xp33_ASAP7_75t_L g1139 ( 
.A(n_1082),
.B(n_977),
.C(n_1074),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_999),
.A2(n_1041),
.B(n_1079),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_948),
.B(n_1072),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_959),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1041),
.A2(n_964),
.B(n_962),
.Y(n_1143)
);

NOR2x1_ASAP7_75t_SL g1144 ( 
.A(n_956),
.B(n_983),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_1051),
.A2(n_1046),
.B(n_1031),
.C(n_1053),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_970),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_978),
.A2(n_1032),
.B(n_1035),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_996),
.Y(n_1148)
);

OAI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1033),
.A2(n_1031),
.B(n_1034),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_949),
.A2(n_1083),
.B(n_948),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1037),
.B(n_1074),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_962),
.A2(n_964),
.B(n_1055),
.Y(n_1152)
);

AO31x2_ASAP7_75t_L g1153 ( 
.A1(n_1055),
.A2(n_973),
.A3(n_1072),
.B(n_987),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_SL g1154 ( 
.A1(n_987),
.A2(n_1074),
.B(n_1034),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1061),
.B(n_956),
.Y(n_1155)
);

INVx3_ASAP7_75t_L g1156 ( 
.A(n_956),
.Y(n_1156)
);

AOI21x1_ASAP7_75t_L g1157 ( 
.A1(n_987),
.A2(n_1055),
.B(n_973),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1081),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_973),
.A2(n_983),
.B(n_1043),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_943),
.A2(n_738),
.B1(n_907),
.B2(n_337),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_961),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_955),
.B(n_880),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_954),
.A2(n_451),
.B(n_812),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1049),
.A2(n_1059),
.B(n_1056),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_1008),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_972),
.A2(n_812),
.B(n_770),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_953),
.Y(n_1167)
);

INVx2_ASAP7_75t_SL g1168 ( 
.A(n_1002),
.Y(n_1168)
);

AO31x2_ASAP7_75t_L g1169 ( 
.A1(n_1060),
.A2(n_972),
.A3(n_951),
.B(n_1056),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_944),
.B(n_812),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_944),
.B(n_812),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_954),
.A2(n_451),
.B(n_812),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_953),
.Y(n_1173)
);

O2A1O1Ixp33_ASAP7_75t_SL g1174 ( 
.A1(n_1026),
.A2(n_812),
.B(n_1023),
.C(n_764),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_944),
.B(n_812),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_960),
.B(n_696),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_954),
.A2(n_451),
.B(n_812),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_953),
.Y(n_1178)
);

INVx8_ASAP7_75t_L g1179 ( 
.A(n_1003),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1049),
.A2(n_1059),
.B(n_1056),
.Y(n_1180)
);

OAI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_972),
.A2(n_812),
.B(n_770),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_SL g1182 ( 
.A(n_1002),
.B(n_533),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_944),
.B(n_812),
.Y(n_1183)
);

NOR2xp67_ASAP7_75t_L g1184 ( 
.A(n_1008),
.B(n_955),
.Y(n_1184)
);

AO31x2_ASAP7_75t_L g1185 ( 
.A1(n_1060),
.A2(n_972),
.A3(n_951),
.B(n_1056),
.Y(n_1185)
);

AO31x2_ASAP7_75t_L g1186 ( 
.A1(n_1060),
.A2(n_972),
.A3(n_951),
.B(n_1056),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_954),
.A2(n_451),
.B(n_812),
.Y(n_1187)
);

AO31x2_ASAP7_75t_L g1188 ( 
.A1(n_1060),
.A2(n_972),
.A3(n_951),
.B(n_1056),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_953),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_954),
.A2(n_451),
.B(n_812),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1049),
.A2(n_1059),
.B(n_1056),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_944),
.B(n_812),
.Y(n_1192)
);

AO31x2_ASAP7_75t_L g1193 ( 
.A1(n_1060),
.A2(n_972),
.A3(n_951),
.B(n_1056),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1049),
.A2(n_1059),
.B(n_1056),
.Y(n_1194)
);

OR2x2_ASAP7_75t_L g1195 ( 
.A(n_960),
.B(n_625),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1049),
.A2(n_1059),
.B(n_1056),
.Y(n_1196)
);

INVx2_ASAP7_75t_SL g1197 ( 
.A(n_1002),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_954),
.A2(n_451),
.B(n_812),
.Y(n_1198)
);

AOI221xp5_ASAP7_75t_L g1199 ( 
.A1(n_1000),
.A2(n_812),
.B1(n_770),
.B2(n_315),
.C(n_340),
.Y(n_1199)
);

INVx3_ASAP7_75t_SL g1200 ( 
.A(n_959),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_961),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_944),
.B(n_812),
.Y(n_1202)
);

OAI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_972),
.A2(n_812),
.B(n_770),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_961),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_960),
.B(n_696),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1049),
.A2(n_1059),
.B(n_1056),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_963),
.B(n_309),
.Y(n_1207)
);

AOI221xp5_ASAP7_75t_SL g1208 ( 
.A1(n_988),
.A2(n_770),
.B1(n_974),
.B2(n_993),
.C(n_1001),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_944),
.B(n_812),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_954),
.A2(n_451),
.B(n_812),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_953),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1049),
.A2(n_1059),
.B(n_1056),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_954),
.A2(n_451),
.B(n_812),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1015),
.A2(n_451),
.B(n_812),
.Y(n_1214)
);

NAND2x1p5_ASAP7_75t_L g1215 ( 
.A(n_955),
.B(n_790),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1015),
.A2(n_451),
.B(n_812),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_972),
.A2(n_812),
.B(n_770),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_953),
.Y(n_1218)
);

OAI22x1_ASAP7_75t_L g1219 ( 
.A1(n_985),
.A2(n_583),
.B1(n_528),
.B2(n_738),
.Y(n_1219)
);

INVx2_ASAP7_75t_SL g1220 ( 
.A(n_1002),
.Y(n_1220)
);

OR2x2_ASAP7_75t_L g1221 ( 
.A(n_960),
.B(n_625),
.Y(n_1221)
);

NOR2xp67_ASAP7_75t_L g1222 ( 
.A(n_1008),
.B(n_955),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1015),
.A2(n_451),
.B(n_812),
.Y(n_1223)
);

CKINVDCx6p67_ASAP7_75t_R g1224 ( 
.A(n_1200),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1176),
.B(n_1205),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1116),
.A2(n_1207),
.B1(n_1199),
.B2(n_1135),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_1165),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_1179),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1199),
.A2(n_1219),
.B1(n_1110),
.B2(n_1125),
.Y(n_1229)
);

OAI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1116),
.A2(n_1114),
.B1(n_1125),
.B2(n_1110),
.Y(n_1230)
);

CKINVDCx6p67_ASAP7_75t_R g1231 ( 
.A(n_1179),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_SL g1232 ( 
.A1(n_1109),
.A2(n_1100),
.B1(n_1182),
.B2(n_1091),
.Y(n_1232)
);

INVx6_ASAP7_75t_L g1233 ( 
.A(n_1096),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_1129),
.Y(n_1234)
);

CKINVDCx6p67_ASAP7_75t_R g1235 ( 
.A(n_1090),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1094),
.A2(n_1195),
.B1(n_1221),
.B2(n_1160),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_SL g1237 ( 
.A1(n_1109),
.A2(n_1100),
.B1(n_1182),
.B2(n_1128),
.Y(n_1237)
);

INVx3_ASAP7_75t_L g1238 ( 
.A(n_1215),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1103),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1115),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1118),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_SL g1242 ( 
.A1(n_1128),
.A2(n_1181),
.B1(n_1217),
.B2(n_1203),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1138),
.A2(n_1137),
.B1(n_1101),
.B2(n_1166),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_1133),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_SL g1245 ( 
.A1(n_1166),
.A2(n_1181),
.B1(n_1217),
.B2(n_1203),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1102),
.A2(n_1192),
.B1(n_1170),
.B2(n_1209),
.Y(n_1246)
);

CKINVDCx11_ASAP7_75t_R g1247 ( 
.A(n_1090),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1148),
.B(n_1119),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1117),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_1104),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_SL g1251 ( 
.A1(n_1101),
.A2(n_1120),
.B1(n_1134),
.B2(n_1087),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1119),
.B(n_1170),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1120),
.A2(n_1209),
.B1(n_1192),
.B2(n_1171),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1171),
.B(n_1175),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1175),
.A2(n_1183),
.B1(n_1202),
.B2(n_1123),
.Y(n_1255)
);

INVx8_ASAP7_75t_L g1256 ( 
.A(n_1090),
.Y(n_1256)
);

BUFx2_ASAP7_75t_SL g1257 ( 
.A(n_1107),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1208),
.A2(n_1141),
.B1(n_1222),
.B2(n_1184),
.Y(n_1258)
);

CKINVDCx11_ASAP7_75t_R g1259 ( 
.A(n_1096),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1167),
.A2(n_1218),
.B1(n_1173),
.B2(n_1178),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1131),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1136),
.Y(n_1262)
);

INVx6_ASAP7_75t_L g1263 ( 
.A(n_1096),
.Y(n_1263)
);

INVx6_ASAP7_75t_L g1264 ( 
.A(n_1162),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1189),
.A2(n_1211),
.B1(n_1151),
.B2(n_1158),
.Y(n_1265)
);

INVx1_ASAP7_75t_SL g1266 ( 
.A(n_1146),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1161),
.A2(n_1204),
.B1(n_1201),
.B2(n_1134),
.Y(n_1267)
);

INVx6_ASAP7_75t_L g1268 ( 
.A(n_1105),
.Y(n_1268)
);

CKINVDCx6p67_ASAP7_75t_R g1269 ( 
.A(n_1155),
.Y(n_1269)
);

BUFx12f_ASAP7_75t_L g1270 ( 
.A(n_1142),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_SL g1271 ( 
.A1(n_1208),
.A2(n_1108),
.B1(n_1150),
.B2(n_1105),
.Y(n_1271)
);

BUFx10_ASAP7_75t_L g1272 ( 
.A(n_1168),
.Y(n_1272)
);

INVxp67_ASAP7_75t_L g1273 ( 
.A(n_1152),
.Y(n_1273)
);

INVxp67_ASAP7_75t_L g1274 ( 
.A(n_1149),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1126),
.A2(n_1139),
.B1(n_1197),
.B2(n_1220),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1126),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1156),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1108),
.A2(n_1149),
.B1(n_1126),
.B2(n_1113),
.Y(n_1278)
);

OAI21xp5_ASAP7_75t_SL g1279 ( 
.A1(n_1132),
.A2(n_1124),
.B(n_1157),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1124),
.A2(n_1223),
.B1(n_1216),
.B2(n_1214),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1145),
.A2(n_1223),
.B1(n_1216),
.B2(n_1214),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1147),
.B(n_1144),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1147),
.A2(n_1098),
.B1(n_1174),
.B2(n_1140),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1095),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1143),
.Y(n_1285)
);

INVxp67_ASAP7_75t_SL g1286 ( 
.A(n_1106),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1127),
.Y(n_1287)
);

INVxp67_ASAP7_75t_SL g1288 ( 
.A(n_1093),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1159),
.Y(n_1289)
);

INVx6_ASAP7_75t_L g1290 ( 
.A(n_1154),
.Y(n_1290)
);

CKINVDCx11_ASAP7_75t_R g1291 ( 
.A(n_1153),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1112),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1121),
.A2(n_1099),
.B1(n_1130),
.B2(n_1122),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1112),
.Y(n_1294)
);

CKINVDCx11_ASAP7_75t_R g1295 ( 
.A(n_1153),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1112),
.Y(n_1296)
);

BUFx8_ASAP7_75t_SL g1297 ( 
.A(n_1089),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1163),
.A2(n_1187),
.B1(n_1210),
.B2(n_1198),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1169),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1172),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1169),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1177),
.A2(n_1213),
.B1(n_1190),
.B2(n_1111),
.Y(n_1302)
);

CKINVDCx20_ASAP7_75t_R g1303 ( 
.A(n_1088),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_SL g1304 ( 
.A1(n_1097),
.A2(n_1188),
.B1(n_1193),
.B2(n_1169),
.Y(n_1304)
);

OAI21xp33_ASAP7_75t_L g1305 ( 
.A1(n_1164),
.A2(n_1212),
.B(n_1180),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_SL g1306 ( 
.A1(n_1191),
.A2(n_1206),
.B1(n_1196),
.B2(n_1194),
.Y(n_1306)
);

CKINVDCx20_ASAP7_75t_R g1307 ( 
.A(n_1193),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1185),
.Y(n_1308)
);

CKINVDCx11_ASAP7_75t_R g1309 ( 
.A(n_1185),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_SL g1310 ( 
.A1(n_1186),
.A2(n_1188),
.B1(n_1193),
.B2(n_1092),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1186),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1186),
.Y(n_1312)
);

CKINVDCx20_ASAP7_75t_R g1313 ( 
.A(n_1188),
.Y(n_1313)
);

INVx6_ASAP7_75t_L g1314 ( 
.A(n_1092),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1092),
.A2(n_460),
.B1(n_745),
.B2(n_750),
.Y(n_1315)
);

OAI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1116),
.A2(n_995),
.B1(n_812),
.B2(n_1000),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1129),
.Y(n_1317)
);

CKINVDCx6p67_ASAP7_75t_R g1318 ( 
.A(n_1200),
.Y(n_1318)
);

INVx6_ASAP7_75t_L g1319 ( 
.A(n_1096),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_1165),
.Y(n_1320)
);

BUFx12f_ASAP7_75t_L g1321 ( 
.A(n_1090),
.Y(n_1321)
);

CKINVDCx11_ASAP7_75t_R g1322 ( 
.A(n_1200),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1176),
.B(n_1205),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_SL g1324 ( 
.A1(n_1116),
.A2(n_460),
.B1(n_1038),
.B2(n_1125),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1176),
.B(n_1205),
.Y(n_1325)
);

CKINVDCx20_ASAP7_75t_R g1326 ( 
.A(n_1104),
.Y(n_1326)
);

CKINVDCx11_ASAP7_75t_R g1327 ( 
.A(n_1200),
.Y(n_1327)
);

OAI22xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1116),
.A2(n_1038),
.B1(n_738),
.B2(n_1125),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_SL g1329 ( 
.A1(n_1116),
.A2(n_460),
.B1(n_1038),
.B2(n_1125),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1176),
.B(n_1205),
.Y(n_1330)
);

INVx6_ASAP7_75t_L g1331 ( 
.A(n_1096),
.Y(n_1331)
);

AOI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1116),
.A2(n_657),
.B1(n_1207),
.B2(n_528),
.Y(n_1332)
);

CKINVDCx20_ASAP7_75t_R g1333 ( 
.A(n_1104),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_1179),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1215),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1179),
.Y(n_1336)
);

BUFx10_ASAP7_75t_L g1337 ( 
.A(n_1165),
.Y(n_1337)
);

CKINVDCx11_ASAP7_75t_R g1338 ( 
.A(n_1200),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1219),
.A2(n_738),
.B1(n_907),
.B2(n_460),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1129),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_1104),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_1215),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1292),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1294),
.B(n_1312),
.Y(n_1344)
);

AO31x2_ASAP7_75t_L g1345 ( 
.A1(n_1281),
.A2(n_1301),
.A3(n_1299),
.B(n_1308),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1248),
.B(n_1296),
.Y(n_1346)
);

AO21x2_ASAP7_75t_L g1347 ( 
.A1(n_1279),
.A2(n_1311),
.B(n_1230),
.Y(n_1347)
);

CKINVDCx20_ASAP7_75t_R g1348 ( 
.A(n_1322),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1245),
.B(n_1242),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1254),
.B(n_1252),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1302),
.A2(n_1298),
.B(n_1293),
.Y(n_1351)
);

OAI222xp33_ASAP7_75t_L g1352 ( 
.A1(n_1324),
.A2(n_1329),
.B1(n_1226),
.B2(n_1229),
.C1(n_1339),
.C2(n_1230),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1285),
.Y(n_1353)
);

INVx3_ASAP7_75t_L g1354 ( 
.A(n_1297),
.Y(n_1354)
);

OA21x2_ASAP7_75t_L g1355 ( 
.A1(n_1305),
.A2(n_1280),
.B(n_1298),
.Y(n_1355)
);

AO21x2_ASAP7_75t_L g1356 ( 
.A1(n_1311),
.A2(n_1316),
.B(n_1288),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1239),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1245),
.B(n_1242),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1323),
.B(n_1330),
.Y(n_1359)
);

AO21x1_ASAP7_75t_L g1360 ( 
.A1(n_1316),
.A2(n_1328),
.B(n_1255),
.Y(n_1360)
);

CKINVDCx12_ASAP7_75t_R g1361 ( 
.A(n_1282),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1240),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1241),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1261),
.Y(n_1364)
);

AND2x4_ASAP7_75t_L g1365 ( 
.A(n_1276),
.B(n_1274),
.Y(n_1365)
);

OR2x2_ASAP7_75t_L g1366 ( 
.A(n_1225),
.B(n_1325),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1262),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1253),
.B(n_1267),
.Y(n_1368)
);

OR2x2_ASAP7_75t_L g1369 ( 
.A(n_1253),
.B(n_1267),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1303),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1280),
.A2(n_1283),
.B(n_1288),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1249),
.B(n_1246),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1274),
.B(n_1307),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1287),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1289),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1313),
.B(n_1309),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1300),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1273),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1314),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1273),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1237),
.B(n_1251),
.Y(n_1381)
);

AO21x2_ASAP7_75t_L g1382 ( 
.A1(n_1286),
.A2(n_1258),
.B(n_1284),
.Y(n_1382)
);

AOI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1277),
.A2(n_1340),
.B(n_1317),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1234),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1251),
.B(n_1243),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1237),
.B(n_1271),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1304),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1286),
.Y(n_1388)
);

INVx11_ASAP7_75t_L g1389 ( 
.A(n_1270),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1310),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1244),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1243),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1271),
.Y(n_1393)
);

OAI21xp5_ASAP7_75t_SL g1394 ( 
.A1(n_1324),
.A2(n_1329),
.B(n_1332),
.Y(n_1394)
);

BUFx4f_ASAP7_75t_L g1395 ( 
.A(n_1231),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1283),
.B(n_1278),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1315),
.A2(n_1291),
.B1(n_1295),
.B2(n_1236),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1278),
.A2(n_1238),
.B(n_1335),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1236),
.B(n_1232),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1264),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1315),
.A2(n_1265),
.B(n_1260),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1306),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1290),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1233),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1233),
.Y(n_1405)
);

INVx1_ASAP7_75t_SL g1406 ( 
.A(n_1266),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1290),
.A2(n_1275),
.B1(n_1269),
.B2(n_1268),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1290),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1256),
.B(n_1235),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1342),
.Y(n_1410)
);

INVx2_ASAP7_75t_SL g1411 ( 
.A(n_1264),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1263),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1256),
.B(n_1224),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1319),
.Y(n_1414)
);

AO21x2_ASAP7_75t_L g1415 ( 
.A1(n_1319),
.A2(n_1331),
.B(n_1272),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_R g1416 ( 
.A(n_1250),
.B(n_1341),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1331),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1272),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1257),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1256),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1365),
.B(n_1373),
.Y(n_1421)
);

A2O1A1Ixp33_ASAP7_75t_L g1422 ( 
.A1(n_1394),
.A2(n_1228),
.B(n_1336),
.C(n_1334),
.Y(n_1422)
);

NOR2x1_ASAP7_75t_SL g1423 ( 
.A(n_1415),
.B(n_1372),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1365),
.B(n_1227),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1370),
.B(n_1337),
.Y(n_1425)
);

NAND4xp25_ASAP7_75t_L g1426 ( 
.A(n_1349),
.B(n_1337),
.C(n_1338),
.D(n_1327),
.Y(n_1426)
);

OAI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1349),
.A2(n_1326),
.B(n_1333),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1370),
.B(n_1247),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1350),
.B(n_1318),
.Y(n_1429)
);

A2O1A1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1399),
.A2(n_1358),
.B(n_1381),
.C(n_1385),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1373),
.B(n_1320),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1364),
.B(n_1259),
.Y(n_1432)
);

NAND2x1_ASAP7_75t_L g1433 ( 
.A(n_1377),
.B(n_1321),
.Y(n_1433)
);

A2O1A1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1399),
.A2(n_1358),
.B(n_1381),
.C(n_1385),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1366),
.B(n_1359),
.Y(n_1435)
);

OAI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1386),
.A2(n_1387),
.B(n_1392),
.Y(n_1436)
);

NAND2xp33_ASAP7_75t_R g1437 ( 
.A(n_1416),
.B(n_1354),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1377),
.B(n_1391),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1360),
.A2(n_1397),
.B1(n_1386),
.B2(n_1376),
.Y(n_1439)
);

INVx4_ASAP7_75t_L g1440 ( 
.A(n_1377),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1406),
.B(n_1413),
.Y(n_1441)
);

BUFx4f_ASAP7_75t_SL g1442 ( 
.A(n_1348),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1384),
.B(n_1376),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1354),
.B(n_1387),
.Y(n_1444)
);

AO32x2_ASAP7_75t_L g1445 ( 
.A1(n_1400),
.A2(n_1411),
.A3(n_1383),
.B1(n_1346),
.B2(n_1390),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1344),
.B(n_1383),
.Y(n_1446)
);

OA21x2_ASAP7_75t_L g1447 ( 
.A1(n_1351),
.A2(n_1371),
.B(n_1402),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1344),
.B(n_1404),
.Y(n_1448)
);

OA21x2_ASAP7_75t_L g1449 ( 
.A1(n_1351),
.A2(n_1371),
.B(n_1402),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1405),
.B(n_1412),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1414),
.Y(n_1451)
);

BUFx5_ASAP7_75t_L g1452 ( 
.A(n_1353),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1378),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1357),
.B(n_1362),
.Y(n_1454)
);

OAI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1352),
.A2(n_1393),
.B(n_1396),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1363),
.B(n_1367),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1414),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1375),
.Y(n_1458)
);

O2A1O1Ixp33_ASAP7_75t_L g1459 ( 
.A1(n_1419),
.A2(n_1347),
.B(n_1418),
.C(n_1396),
.Y(n_1459)
);

OAI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1396),
.A2(n_1369),
.B(n_1368),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1419),
.B(n_1409),
.Y(n_1461)
);

NOR2x1_ASAP7_75t_SL g1462 ( 
.A(n_1382),
.B(n_1356),
.Y(n_1462)
);

OAI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1396),
.A2(n_1368),
.B(n_1369),
.Y(n_1463)
);

OAI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1374),
.A2(n_1398),
.B(n_1380),
.Y(n_1464)
);

AND2x2_ASAP7_75t_SL g1465 ( 
.A(n_1361),
.B(n_1407),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1343),
.B(n_1353),
.Y(n_1466)
);

AOI221xp5_ASAP7_75t_L g1467 ( 
.A1(n_1343),
.A2(n_1356),
.B1(n_1388),
.B2(n_1418),
.C(n_1410),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1452),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1447),
.B(n_1355),
.Y(n_1469)
);

INVxp67_ASAP7_75t_SL g1470 ( 
.A(n_1453),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1458),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1454),
.B(n_1382),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1447),
.B(n_1355),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1449),
.B(n_1355),
.Y(n_1474)
);

INVxp67_ASAP7_75t_SL g1475 ( 
.A(n_1462),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1449),
.B(n_1355),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1455),
.A2(n_1401),
.B1(n_1408),
.B2(n_1403),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1455),
.A2(n_1401),
.B1(n_1408),
.B2(n_1403),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1466),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1446),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1421),
.B(n_1388),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1421),
.B(n_1345),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1448),
.B(n_1345),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1452),
.B(n_1345),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1456),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1443),
.B(n_1379),
.Y(n_1486)
);

INVx3_ASAP7_75t_L g1487 ( 
.A(n_1440),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1451),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1426),
.B(n_1417),
.Y(n_1489)
);

BUFx2_ASAP7_75t_L g1490 ( 
.A(n_1440),
.Y(n_1490)
);

AOI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1477),
.A2(n_1439),
.B1(n_1430),
.B2(n_1434),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1471),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1469),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1469),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1480),
.B(n_1450),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1471),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1480),
.B(n_1445),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1471),
.Y(n_1498)
);

A2O1A1Ixp33_ASAP7_75t_L g1499 ( 
.A1(n_1477),
.A2(n_1459),
.B(n_1427),
.C(n_1436),
.Y(n_1499)
);

INVxp67_ASAP7_75t_SL g1500 ( 
.A(n_1470),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1469),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1483),
.B(n_1445),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1469),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1476),
.Y(n_1504)
);

AOI221xp5_ASAP7_75t_L g1505 ( 
.A1(n_1472),
.A2(n_1427),
.B1(n_1463),
.B2(n_1460),
.C(n_1467),
.Y(n_1505)
);

OAI211xp5_ASAP7_75t_L g1506 ( 
.A1(n_1475),
.A2(n_1426),
.B(n_1422),
.C(n_1429),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1483),
.B(n_1445),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1470),
.B(n_1435),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1483),
.B(n_1423),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1475),
.Y(n_1510)
);

INVx4_ASAP7_75t_L g1511 ( 
.A(n_1487),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1486),
.B(n_1438),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1486),
.B(n_1481),
.Y(n_1513)
);

INVxp67_ASAP7_75t_L g1514 ( 
.A(n_1488),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1481),
.B(n_1457),
.Y(n_1515)
);

NAND3xp33_ASAP7_75t_L g1516 ( 
.A(n_1476),
.B(n_1463),
.C(n_1460),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1489),
.B(n_1432),
.Y(n_1517)
);

INVx2_ASAP7_75t_SL g1518 ( 
.A(n_1490),
.Y(n_1518)
);

OAI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1478),
.A2(n_1465),
.B(n_1464),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1473),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1473),
.Y(n_1521)
);

AOI21xp33_ASAP7_75t_SL g1522 ( 
.A1(n_1489),
.A2(n_1437),
.B(n_1428),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1473),
.Y(n_1523)
);

NAND4xp25_ASAP7_75t_L g1524 ( 
.A(n_1478),
.B(n_1425),
.C(n_1461),
.D(n_1431),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1492),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1497),
.B(n_1488),
.Y(n_1526)
);

INVx2_ASAP7_75t_SL g1527 ( 
.A(n_1510),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1500),
.B(n_1485),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1497),
.B(n_1481),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1492),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1500),
.B(n_1485),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1498),
.Y(n_1532)
);

INVxp67_ASAP7_75t_SL g1533 ( 
.A(n_1514),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1514),
.B(n_1479),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1497),
.B(n_1484),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1493),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1508),
.B(n_1493),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1498),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1513),
.B(n_1493),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1513),
.B(n_1484),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1496),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1513),
.B(n_1484),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1496),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1494),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1508),
.B(n_1479),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1494),
.B(n_1479),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1501),
.B(n_1482),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1511),
.B(n_1482),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1511),
.B(n_1468),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1533),
.B(n_1505),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1525),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1539),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1525),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1544),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1540),
.B(n_1495),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1530),
.Y(n_1556)
);

OAI211xp5_ASAP7_75t_SL g1557 ( 
.A1(n_1533),
.A2(n_1506),
.B(n_1499),
.C(n_1517),
.Y(n_1557)
);

NOR2x1p5_ASAP7_75t_SL g1558 ( 
.A(n_1544),
.B(n_1503),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1548),
.B(n_1522),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1539),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1530),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1540),
.B(n_1495),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1532),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1532),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1540),
.B(n_1495),
.Y(n_1565)
);

INVx2_ASAP7_75t_SL g1566 ( 
.A(n_1548),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1538),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1534),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1545),
.B(n_1505),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1545),
.B(n_1512),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1534),
.B(n_1503),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1538),
.Y(n_1572)
);

INVxp67_ASAP7_75t_L g1573 ( 
.A(n_1528),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1548),
.B(n_1510),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1541),
.Y(n_1575)
);

NOR2x1_ASAP7_75t_L g1576 ( 
.A(n_1528),
.B(n_1524),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1541),
.Y(n_1577)
);

OAI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1527),
.A2(n_1499),
.B(n_1516),
.Y(n_1578)
);

AND2x2_ASAP7_75t_SL g1579 ( 
.A(n_1526),
.B(n_1510),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1543),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1539),
.Y(n_1581)
);

BUFx2_ASAP7_75t_L g1582 ( 
.A(n_1527),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1531),
.B(n_1504),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1531),
.B(n_1504),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1543),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1526),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1547),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1547),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1542),
.B(n_1515),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1537),
.B(n_1504),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1548),
.B(n_1511),
.Y(n_1591)
);

NAND2x1p5_ASAP7_75t_L g1592 ( 
.A(n_1576),
.B(n_1395),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1550),
.B(n_1537),
.Y(n_1593)
);

NOR3xp33_ASAP7_75t_L g1594 ( 
.A(n_1557),
.B(n_1506),
.C(n_1522),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1569),
.B(n_1537),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1555),
.B(n_1542),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1568),
.B(n_1546),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_SL g1598 ( 
.A(n_1579),
.B(n_1527),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1551),
.Y(n_1599)
);

INVx3_ASAP7_75t_L g1600 ( 
.A(n_1579),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1551),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1555),
.B(n_1542),
.Y(n_1602)
);

NAND4xp75_ASAP7_75t_L g1603 ( 
.A(n_1576),
.B(n_1519),
.C(n_1491),
.D(n_1507),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1573),
.B(n_1526),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1578),
.B(n_1562),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1562),
.B(n_1529),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1565),
.B(n_1529),
.Y(n_1607)
);

NAND4xp75_ASAP7_75t_L g1608 ( 
.A(n_1579),
.B(n_1558),
.C(n_1519),
.D(n_1491),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1565),
.B(n_1529),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1589),
.B(n_1548),
.Y(n_1610)
);

INVx1_ASAP7_75t_SL g1611 ( 
.A(n_1582),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1586),
.B(n_1535),
.Y(n_1612)
);

NOR2x1_ASAP7_75t_L g1613 ( 
.A(n_1582),
.B(n_1524),
.Y(n_1613)
);

NAND2x1p5_ASAP7_75t_L g1614 ( 
.A(n_1559),
.B(n_1395),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1589),
.B(n_1535),
.Y(n_1615)
);

INVxp67_ASAP7_75t_SL g1616 ( 
.A(n_1554),
.Y(n_1616)
);

INVxp67_ASAP7_75t_L g1617 ( 
.A(n_1553),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1570),
.B(n_1442),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1552),
.B(n_1535),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1552),
.B(n_1547),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1560),
.B(n_1546),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1553),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1560),
.B(n_1546),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1566),
.B(n_1517),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1581),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1556),
.Y(n_1626)
);

NOR3xp33_ASAP7_75t_L g1627 ( 
.A(n_1603),
.B(n_1608),
.C(n_1594),
.Y(n_1627)
);

OAI21x1_ASAP7_75t_SL g1628 ( 
.A1(n_1613),
.A2(n_1566),
.B(n_1581),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1615),
.B(n_1587),
.Y(n_1629)
);

INVxp67_ASAP7_75t_SL g1630 ( 
.A(n_1592),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1595),
.B(n_1611),
.Y(n_1631)
);

NOR2x1_ASAP7_75t_L g1632 ( 
.A(n_1608),
.B(n_1574),
.Y(n_1632)
);

O2A1O1Ixp33_ASAP7_75t_SL g1633 ( 
.A1(n_1598),
.A2(n_1518),
.B(n_1433),
.C(n_1588),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1595),
.B(n_1587),
.Y(n_1634)
);

AOI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1603),
.A2(n_1502),
.B1(n_1507),
.B2(n_1516),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1599),
.Y(n_1636)
);

AOI21xp33_ASAP7_75t_SL g1637 ( 
.A1(n_1592),
.A2(n_1574),
.B(n_1591),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1593),
.B(n_1588),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1592),
.B(n_1574),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1593),
.B(n_1558),
.Y(n_1640)
);

NAND2x1_ASAP7_75t_L g1641 ( 
.A(n_1600),
.B(n_1574),
.Y(n_1641)
);

OAI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1605),
.A2(n_1509),
.B1(n_1507),
.B2(n_1502),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1601),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1618),
.B(n_1389),
.Y(n_1644)
);

OAI211xp5_ASAP7_75t_L g1645 ( 
.A1(n_1600),
.A2(n_1617),
.B(n_1604),
.C(n_1624),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1622),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1626),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1596),
.Y(n_1648)
);

NOR3xp33_ASAP7_75t_L g1649 ( 
.A(n_1600),
.B(n_1554),
.C(n_1563),
.Y(n_1649)
);

AOI211xp5_ASAP7_75t_L g1650 ( 
.A1(n_1619),
.A2(n_1583),
.B(n_1584),
.C(n_1590),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1625),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_SL g1652 ( 
.A(n_1614),
.B(n_1591),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1627),
.B(n_1616),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1648),
.B(n_1615),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1631),
.B(n_1607),
.Y(n_1655)
);

OAI221xp5_ASAP7_75t_SL g1656 ( 
.A1(n_1635),
.A2(n_1612),
.B1(n_1597),
.B2(n_1619),
.C(n_1623),
.Y(n_1656)
);

OAI22xp33_ASAP7_75t_L g1657 ( 
.A1(n_1642),
.A2(n_1614),
.B1(n_1509),
.B2(n_1609),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1643),
.Y(n_1658)
);

OAI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1642),
.A2(n_1614),
.B1(n_1502),
.B2(n_1625),
.Y(n_1659)
);

OAI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1640),
.A2(n_1521),
.B1(n_1523),
.B2(n_1520),
.Y(n_1660)
);

AOI32xp33_ASAP7_75t_L g1661 ( 
.A1(n_1632),
.A2(n_1620),
.A3(n_1606),
.B1(n_1596),
.B2(n_1602),
.Y(n_1661)
);

INVx1_ASAP7_75t_SL g1662 ( 
.A(n_1634),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1643),
.Y(n_1663)
);

OAI21xp33_ASAP7_75t_L g1664 ( 
.A1(n_1645),
.A2(n_1606),
.B(n_1602),
.Y(n_1664)
);

OAI31xp33_ASAP7_75t_L g1665 ( 
.A1(n_1649),
.A2(n_1597),
.A3(n_1620),
.B(n_1474),
.Y(n_1665)
);

NAND3xp33_ASAP7_75t_SL g1666 ( 
.A(n_1650),
.B(n_1610),
.C(n_1621),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1638),
.B(n_1621),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1651),
.Y(n_1668)
);

NOR2xp67_ASAP7_75t_L g1669 ( 
.A(n_1637),
.B(n_1623),
.Y(n_1669)
);

NOR3xp33_ASAP7_75t_L g1670 ( 
.A(n_1630),
.B(n_1554),
.C(n_1572),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1641),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1662),
.B(n_1629),
.Y(n_1672)
);

AO22x1_ASAP7_75t_L g1673 ( 
.A1(n_1653),
.A2(n_1630),
.B1(n_1644),
.B2(n_1646),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1654),
.Y(n_1674)
);

NAND2xp33_ASAP7_75t_SL g1675 ( 
.A(n_1653),
.B(n_1636),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1662),
.Y(n_1676)
);

CKINVDCx14_ASAP7_75t_R g1677 ( 
.A(n_1658),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1663),
.Y(n_1678)
);

OAI21xp33_ASAP7_75t_L g1679 ( 
.A1(n_1664),
.A2(n_1639),
.B(n_1652),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1667),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1668),
.Y(n_1681)
);

AOI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1675),
.A2(n_1628),
.B(n_1656),
.Y(n_1682)
);

OAI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1675),
.A2(n_1666),
.B(n_1669),
.Y(n_1683)
);

NAND4xp25_ASAP7_75t_L g1684 ( 
.A(n_1679),
.B(n_1661),
.C(n_1655),
.D(n_1671),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1672),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1674),
.B(n_1644),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1673),
.B(n_1670),
.Y(n_1687)
);

NAND3xp33_ASAP7_75t_SL g1688 ( 
.A(n_1676),
.B(n_1665),
.C(n_1647),
.Y(n_1688)
);

NOR3xp33_ASAP7_75t_SL g1689 ( 
.A(n_1680),
.B(n_1657),
.C(n_1659),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1677),
.B(n_1610),
.Y(n_1690)
);

OAI221xp5_ASAP7_75t_L g1691 ( 
.A1(n_1683),
.A2(n_1681),
.B1(n_1678),
.B2(n_1633),
.C(n_1677),
.Y(n_1691)
);

INVxp67_ASAP7_75t_L g1692 ( 
.A(n_1686),
.Y(n_1692)
);

OAI221xp5_ASAP7_75t_SL g1693 ( 
.A1(n_1682),
.A2(n_1660),
.B1(n_1590),
.B2(n_1583),
.C(n_1584),
.Y(n_1693)
);

AND4x2_ASAP7_75t_L g1694 ( 
.A(n_1684),
.B(n_1389),
.C(n_1591),
.D(n_1395),
.Y(n_1694)
);

NOR2xp67_ASAP7_75t_L g1695 ( 
.A(n_1690),
.B(n_1556),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1692),
.Y(n_1696)
);

NAND4xp25_ASAP7_75t_L g1697 ( 
.A(n_1691),
.B(n_1685),
.C(n_1687),
.D(n_1688),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1695),
.B(n_1689),
.Y(n_1698)
);

AOI222xp33_ASAP7_75t_L g1699 ( 
.A1(n_1693),
.A2(n_1474),
.B1(n_1563),
.B2(n_1561),
.C1(n_1572),
.C2(n_1567),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1694),
.B(n_1561),
.Y(n_1700)
);

AOI221x1_ASAP7_75t_L g1701 ( 
.A1(n_1694),
.A2(n_1567),
.B1(n_1564),
.B2(n_1585),
.C(n_1580),
.Y(n_1701)
);

NOR2x1_ASAP7_75t_L g1702 ( 
.A(n_1697),
.B(n_1591),
.Y(n_1702)
);

NOR2x1_ASAP7_75t_L g1703 ( 
.A(n_1696),
.B(n_1564),
.Y(n_1703)
);

NOR2x1_ASAP7_75t_L g1704 ( 
.A(n_1698),
.B(n_1575),
.Y(n_1704)
);

OAI211xp5_ASAP7_75t_L g1705 ( 
.A1(n_1700),
.A2(n_1585),
.B(n_1580),
.C(n_1577),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1701),
.B(n_1431),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1704),
.Y(n_1707)
);

BUFx6f_ASAP7_75t_L g1708 ( 
.A(n_1706),
.Y(n_1708)
);

NAND3xp33_ASAP7_75t_L g1709 ( 
.A(n_1702),
.B(n_1699),
.C(n_1577),
.Y(n_1709)
);

INVxp67_ASAP7_75t_L g1710 ( 
.A(n_1708),
.Y(n_1710)
);

INVx1_ASAP7_75t_SL g1711 ( 
.A(n_1710),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1711),
.B(n_1707),
.Y(n_1712)
);

BUFx2_ASAP7_75t_L g1713 ( 
.A(n_1711),
.Y(n_1713)
);

AOI22x1_ASAP7_75t_L g1714 ( 
.A1(n_1713),
.A2(n_1703),
.B1(n_1709),
.B2(n_1705),
.Y(n_1714)
);

AOI21xp5_ASAP7_75t_L g1715 ( 
.A1(n_1712),
.A2(n_1575),
.B(n_1571),
.Y(n_1715)
);

OAI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1714),
.A2(n_1571),
.B1(n_1544),
.B2(n_1536),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1715),
.Y(n_1717)
);

AOI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1717),
.A2(n_1716),
.B1(n_1544),
.B2(n_1536),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1718),
.B(n_1441),
.Y(n_1719)
);

CKINVDCx20_ASAP7_75t_R g1720 ( 
.A(n_1719),
.Y(n_1720)
);

OAI221xp5_ASAP7_75t_R g1721 ( 
.A1(n_1720),
.A2(n_1518),
.B1(n_1536),
.B2(n_1549),
.C(n_1409),
.Y(n_1721)
);

AOI211xp5_ASAP7_75t_L g1722 ( 
.A1(n_1721),
.A2(n_1444),
.B(n_1420),
.C(n_1424),
.Y(n_1722)
);


endmodule