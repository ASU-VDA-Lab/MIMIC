module fake_jpeg_31914_n_100 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_100);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_100;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_15),
.B(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_8),
.B(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_45),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_42),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_47),
.B(n_50),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_36),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_1),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

AND2x4_ASAP7_75t_SL g53 ( 
.A(n_45),
.B(n_39),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_4),
.C(n_5),
.Y(n_72)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_50),
.B(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_6),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_48),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_3),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_48),
.A2(n_49),
.B1(n_46),
.B2(n_35),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_60),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_68)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_43),
.B1(n_38),
.B2(n_34),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_65),
.B1(n_25),
.B2(n_32),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_SL g65 ( 
.A1(n_53),
.A2(n_39),
.B(n_16),
.C(n_19),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_59),
.A2(n_37),
.B1(n_39),
.B2(n_14),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_68),
.B1(n_9),
.B2(n_10),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_1),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_72),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_21),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_54),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_74),
.A2(n_62),
.B1(n_61),
.B2(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_7),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_78),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_80),
.A2(n_83),
.B(n_75),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

AND2x6_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_27),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_58),
.C(n_61),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_64),
.C(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_87),
.B(n_90),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_82),
.Y(n_93)
);

OA21x2_ASAP7_75t_SL g94 ( 
.A1(n_93),
.A2(n_65),
.B(n_83),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_92),
.B(n_76),
.Y(n_95)
);

AOI322xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_81),
.A3(n_88),
.B1(n_78),
.B2(n_93),
.C1(n_89),
.C2(n_86),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_20),
.Y(n_97)
);

AOI322xp5_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_22),
.A3(n_28),
.B1(n_30),
.B2(n_79),
.C1(n_9),
.C2(n_11),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_98),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_11),
.Y(n_100)
);


endmodule