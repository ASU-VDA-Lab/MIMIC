module fake_jpeg_680_n_135 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_135);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_24),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_22),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_48),
.Y(n_57)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_53),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_52),
.A2(n_45),
.B1(n_42),
.B2(n_47),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_48),
.A2(n_39),
.B1(n_44),
.B2(n_42),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_43),
.B1(n_47),
.B2(n_49),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_44),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_62),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_51),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_35),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_41),
.Y(n_76)
);

O2A1O1Ixp33_ASAP7_75t_SL g65 ( 
.A1(n_59),
.A2(n_53),
.B(n_49),
.C(n_54),
.Y(n_65)
);

OAI32xp33_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_58),
.A3(n_61),
.B1(n_6),
.B2(n_7),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_46),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_55),
.B(n_36),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_68),
.B(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_37),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_72),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_37),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_43),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_77),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_58),
.B1(n_61),
.B2(n_6),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_39),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_56),
.C(n_57),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_57),
.B(n_3),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_80),
.C(n_84),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_64),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_76),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_83),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_58),
.C(n_61),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_90),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_34),
.B1(n_29),
.B2(n_28),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_18),
.C(n_33),
.Y(n_90)
);

OAI22x1_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_71),
.B1(n_19),
.B2(n_20),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_93),
.B1(n_96),
.B2(n_104),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_16),
.B1(n_31),
.B2(n_30),
.Y(n_93)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_99),
.Y(n_106)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_88),
.A2(n_4),
.B(n_5),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_15),
.B(n_25),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_4),
.B(n_5),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_102),
.A2(n_11),
.B(n_12),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_82),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_103),
.B(n_14),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_27),
.Y(n_104)
);

NOR3xp33_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_15),
.C(n_17),
.Y(n_113)
);

AOI322xp5_ASAP7_75t_SL g105 ( 
.A1(n_94),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_11),
.C1(n_12),
.C2(n_14),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_105),
.B(n_108),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_98),
.B(n_26),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_91),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_9),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_112),
.B(n_113),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_110),
.Y(n_118)
);

BUFx24_ASAP7_75t_SL g111 ( 
.A(n_102),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_111),
.A2(n_114),
.B(n_117),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_115),
.A2(n_116),
.B1(n_101),
.B2(n_98),
.Y(n_123)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_101),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_122),
.B(n_123),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_107),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_122),
.C(n_118),
.Y(n_127)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_126),
.C(n_120),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_121),
.B(n_109),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_124),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_130),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

BUFx24_ASAP7_75t_SL g133 ( 
.A(n_132),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_127),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_128),
.Y(n_135)
);


endmodule