module fake_jpeg_7990_n_275 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_275);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_275;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_27),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_43),
.B(n_34),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_33),
.B1(n_32),
.B2(n_31),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_45),
.A2(n_50),
.B(n_53),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_24),
.B(n_33),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_30),
.Y(n_68)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_33),
.B1(n_32),
.B2(n_31),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_31),
.B1(n_21),
.B2(n_24),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_57),
.B1(n_42),
.B2(n_29),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_52),
.B(n_54),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_30),
.B1(n_29),
.B2(n_26),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_43),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_30),
.B1(n_29),
.B2(n_26),
.Y(n_57)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_61),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_34),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_63),
.Y(n_67)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_64),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_66),
.A2(n_71),
.B1(n_81),
.B2(n_83),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_68),
.A2(n_82),
.B(n_85),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_40),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_69),
.B(n_72),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_41),
.B1(n_26),
.B2(n_18),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_70),
.A2(n_92),
.B1(n_100),
.B2(n_36),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_59),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_40),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_74),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_61),
.Y(n_74)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_77),
.Y(n_103)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_78),
.B(n_79),
.Y(n_121)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_49),
.A2(n_17),
.B1(n_18),
.B2(n_20),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_41),
.C(n_38),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_87),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_41),
.C(n_38),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_25),
.Y(n_87)
);

AO22x1_ASAP7_75t_SL g88 ( 
.A1(n_45),
.A2(n_50),
.B1(n_57),
.B2(n_53),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_88),
.A2(n_93),
.B1(n_95),
.B2(n_0),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_20),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_90),
.Y(n_105)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_49),
.A2(n_23),
.B1(n_19),
.B2(n_28),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_60),
.A2(n_25),
.B1(n_22),
.B2(n_28),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_40),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_99),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_62),
.A2(n_22),
.B1(n_17),
.B2(n_23),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_60),
.A2(n_23),
.B1(n_28),
.B2(n_19),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_27),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_98),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_46),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_63),
.A2(n_28),
.B1(n_19),
.B2(n_27),
.Y(n_100)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_111),
.Y(n_144)
);

NOR2x1_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_70),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_108),
.A2(n_89),
.B(n_65),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_89),
.A2(n_19),
.B1(n_46),
.B2(n_36),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_110),
.A2(n_118),
.B1(n_115),
.B2(n_128),
.Y(n_153)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_114),
.B(n_112),
.Y(n_143)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_119),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_68),
.A2(n_40),
.B(n_27),
.C(n_36),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_92),
.B(n_78),
.C(n_40),
.Y(n_147)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_122),
.B1(n_126),
.B2(n_105),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_88),
.A2(n_36),
.B1(n_40),
.B2(n_56),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_68),
.B(n_56),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_96),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_88),
.A2(n_40),
.B1(n_16),
.B2(n_3),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_72),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_127),
.A2(n_73),
.B1(n_75),
.B2(n_77),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_128),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_129),
.A2(n_104),
.B(n_5),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_85),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_132),
.C(n_134),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_131),
.A2(n_133),
.B1(n_139),
.B2(n_101),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_82),
.C(n_76),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_76),
.B1(n_97),
.B2(n_90),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_65),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_136),
.Y(n_166)
);

NOR3xp33_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_97),
.C(n_74),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_137),
.A2(n_145),
.B(n_147),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_121),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_146),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_108),
.B(n_93),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_157),
.C(n_101),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_152),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_112),
.A2(n_99),
.B(n_100),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_84),
.Y(n_148)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_79),
.Y(n_149)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_149),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_153),
.B1(n_126),
.B2(n_120),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_91),
.Y(n_151)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_1),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_113),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_155),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_103),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_109),
.Y(n_156)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_156),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_111),
.B(n_64),
.C(n_80),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_161),
.A2(n_163),
.B1(n_131),
.B2(n_147),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_127),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_162),
.B(n_167),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_141),
.A2(n_110),
.B1(n_125),
.B2(n_118),
.Y(n_163)
);

OAI32xp33_ASAP7_75t_L g198 ( 
.A1(n_168),
.A2(n_153),
.A3(n_155),
.B1(n_133),
.B2(n_150),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_129),
.A2(n_102),
.B1(n_106),
.B2(n_123),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_169),
.A2(n_138),
.B1(n_157),
.B2(n_83),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_142),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_176),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_132),
.B(n_102),
.C(n_123),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_177),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_109),
.Y(n_173)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_119),
.C(n_117),
.Y(n_177)
);

A2O1A1O1Ixp25_ASAP7_75t_L g179 ( 
.A1(n_145),
.A2(n_3),
.B(n_4),
.C(n_5),
.D(n_6),
.Y(n_179)
);

A2O1A1O1Ixp25_ASAP7_75t_L g196 ( 
.A1(n_179),
.A2(n_180),
.B(n_4),
.C(n_6),
.D(n_7),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_144),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_183),
.Y(n_186)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_140),
.Y(n_187)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_188),
.A2(n_205),
.B1(n_171),
.B2(n_159),
.Y(n_216)
);

INVxp33_ASAP7_75t_SL g189 ( 
.A(n_158),
.Y(n_189)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_166),
.B(n_154),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_191),
.B(n_193),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_156),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_178),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_195),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_146),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_179),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_161),
.A2(n_163),
.B1(n_169),
.B2(n_137),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_197),
.A2(n_165),
.B1(n_177),
.B2(n_175),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_198),
.A2(n_199),
.B1(n_180),
.B2(n_172),
.Y(n_208)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_201),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_109),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_204),
.Y(n_221)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_164),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_165),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_9),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_162),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_192),
.Y(n_224)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_199),
.A2(n_158),
.B1(n_183),
.B2(n_160),
.Y(n_209)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_211),
.B(n_191),
.Y(n_226)
);

AOI21x1_ASAP7_75t_L g213 ( 
.A1(n_190),
.A2(n_171),
.B(n_167),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_197),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_216),
.A2(n_219),
.B1(n_206),
.B2(n_202),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_217),
.A2(n_188),
.B1(n_198),
.B2(n_205),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_190),
.A2(n_174),
.B(n_175),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_9),
.C(n_11),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_222),
.C(n_185),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_9),
.C(n_11),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_12),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_230),
.C(n_235),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_226),
.Y(n_242)
);

NAND3xp33_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_194),
.C(n_200),
.Y(n_227)
);

AOI21xp33_ASAP7_75t_L g249 ( 
.A1(n_227),
.A2(n_210),
.B(n_219),
.Y(n_249)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_212),
.B(n_186),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_229),
.B(n_232),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_216),
.A2(n_204),
.B1(n_196),
.B2(n_14),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_233),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_221),
.Y(n_234)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_15),
.C(n_12),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_236),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_217),
.A2(n_13),
.B1(n_15),
.B2(n_214),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_238),
.A2(n_222),
.B1(n_210),
.B2(n_220),
.Y(n_248)
);

FAx1_ASAP7_75t_SL g241 ( 
.A(n_230),
.B(n_221),
.CI(n_223),
.CON(n_241),
.SN(n_241)
);

OAI321xp33_ASAP7_75t_L g256 ( 
.A1(n_241),
.A2(n_249),
.A3(n_237),
.B1(n_234),
.B2(n_211),
.C(n_235),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_231),
.A2(n_214),
.B1(n_215),
.B2(n_218),
.Y(n_246)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_246),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_248),
.Y(n_252)
);

NAND3xp33_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_238),
.C(n_225),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_250),
.B(n_251),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_224),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_236),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_255),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_244),
.B(n_232),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_256),
.A2(n_243),
.B(n_248),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_13),
.C(n_245),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_13),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_260),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_253),
.A2(n_243),
.B1(n_247),
.B2(n_245),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_252),
.C(n_239),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_241),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_242),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_259),
.Y(n_264)
);

INVxp33_ASAP7_75t_L g270 ( 
.A(n_264),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_258),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_266),
.B(n_263),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_268),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_269),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_271),
.B(n_267),
.C(n_270),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_272),
.C(n_250),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_241),
.Y(n_275)
);


endmodule