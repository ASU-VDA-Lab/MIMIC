module fake_jpeg_24525_n_220 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_220);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_220;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_4),
.B(n_2),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_35),
.B(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_21),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx2_ASAP7_75t_SL g49 ( 
.A(n_37),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_38),
.B(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_44),
.A2(n_26),
.B1(n_18),
.B2(n_27),
.Y(n_48)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_48),
.A2(n_44),
.B1(n_40),
.B2(n_34),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_27),
.B1(n_18),
.B2(n_24),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_50),
.A2(n_51),
.B1(n_36),
.B2(n_21),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_27),
.B1(n_26),
.B2(n_24),
.Y(n_51)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_33),
.Y(n_55)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_69),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_29),
.Y(n_57)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_32),
.B1(n_19),
.B2(n_28),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_59),
.A2(n_64),
.B1(n_23),
.B2(n_25),
.Y(n_92)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_66),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_43),
.A2(n_32),
.B1(n_19),
.B2(n_28),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_70),
.Y(n_100)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_35),
.B(n_21),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_42),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_86),
.C(n_89),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_31),
.B(n_34),
.C(n_22),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_75),
.A2(n_97),
.B1(n_61),
.B2(n_46),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_41),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_84),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_77),
.A2(n_80),
.B1(n_87),
.B2(n_92),
.Y(n_119)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_83),
.Y(n_120)
);

NOR2x1_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_22),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_81),
.B(n_93),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_53),
.B(n_16),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_82),
.B(n_85),
.Y(n_115)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_41),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_36),
.C(n_41),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_39),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_99),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_39),
.C(n_16),
.Y(n_89)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_67),
.A2(n_29),
.B1(n_25),
.B2(n_23),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_98),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_17),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_30),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_124),
.Y(n_132)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_106),
.Y(n_145)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_65),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_78),
.B(n_80),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_110),
.B(n_128),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_100),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_117),
.Y(n_146)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_121),
.Y(n_147)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_126),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_92),
.A2(n_61),
.B1(n_46),
.B2(n_65),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_85),
.B1(n_74),
.B2(n_86),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_65),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_17),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_30),
.Y(n_140)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_127),
.Y(n_138)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_129),
.A2(n_134),
.B1(n_137),
.B2(n_109),
.Y(n_151)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_131),
.B(n_133),
.Y(n_166)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_106),
.A2(n_76),
.B1(n_89),
.B2(n_97),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_135),
.A2(n_110),
.B(n_115),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_105),
.B(n_90),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_140),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_125),
.A2(n_78),
.B1(n_83),
.B2(n_79),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_124),
.A2(n_17),
.B1(n_30),
.B2(n_91),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_139),
.A2(n_123),
.B1(n_109),
.B2(n_128),
.Y(n_152)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_142),
.Y(n_163)
);

AND2x6_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_1),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_148),
.Y(n_162)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_102),
.B(n_3),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_108),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_112),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_151),
.A2(n_148),
.B1(n_143),
.B2(n_133),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_152),
.A2(n_156),
.B1(n_137),
.B2(n_147),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_149),
.A2(n_120),
.B(n_112),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_153),
.A2(n_161),
.B(n_130),
.Y(n_171)
);

BUFx24_ASAP7_75t_SL g154 ( 
.A(n_141),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_154),
.B(n_167),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_145),
.A2(n_142),
.B1(n_135),
.B2(n_138),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_157),
.A2(n_160),
.B(n_165),
.Y(n_176)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_119),
.B(n_113),
.Y(n_160)
);

AO22x1_ASAP7_75t_L g161 ( 
.A1(n_129),
.A2(n_122),
.B1(n_114),
.B2(n_103),
.Y(n_161)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_132),
.A2(n_104),
.B(n_117),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_138),
.B(n_15),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_168),
.A2(n_170),
.B1(n_171),
.B2(n_177),
.Y(n_190)
);

NAND3xp33_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_131),
.C(n_140),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_164),
.Y(n_182)
);

AND3x1_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_130),
.C(n_134),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_136),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_175),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_174),
.A2(n_179),
.B1(n_181),
.B2(n_170),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_139),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_161),
.A2(n_146),
.B1(n_144),
.B2(n_150),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_156),
.A2(n_150),
.B1(n_144),
.B2(n_15),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_13),
.C(n_12),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_167),
.C(n_157),
.Y(n_192)
);

AO22x1_ASAP7_75t_L g198 ( 
.A1(n_182),
.A2(n_175),
.B1(n_5),
.B2(n_6),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_162),
.C(n_153),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_186),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_184),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_162),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_152),
.C(n_158),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_188),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_158),
.C(n_166),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_178),
.B(n_155),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_189),
.A2(n_192),
.B(n_163),
.Y(n_193)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_191),
.B(n_179),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_193),
.A2(n_196),
.B(n_199),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_194),
.B(n_200),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_L g196 ( 
.A1(n_190),
.A2(n_172),
.B(n_155),
.Y(n_196)
);

NOR2xp67_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_6),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_183),
.A2(n_173),
.B(n_5),
.Y(n_199)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_192),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_185),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_203),
.C(n_196),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_185),
.C(n_186),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_205),
.A2(n_203),
.B1(n_206),
.B2(n_204),
.Y(n_211)
);

OAI21x1_ASAP7_75t_L g208 ( 
.A1(n_207),
.A2(n_198),
.B(n_201),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_208),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_209),
.A2(n_211),
.B(n_8),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_7),
.C(n_8),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_210),
.A2(n_8),
.B(n_9),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_213),
.B(n_9),
.C(n_10),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_214),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_215),
.A2(n_11),
.B1(n_208),
.B2(n_212),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_212),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_217),
.B(n_218),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_217),
.Y(n_220)
);


endmodule