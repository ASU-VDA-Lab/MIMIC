module fake_netlist_6_3967_n_542 (n_52, n_16, n_1, n_46, n_18, n_21, n_3, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_77, n_42, n_8, n_24, n_54, n_0, n_32, n_66, n_85, n_78, n_84, n_13, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_45, n_34, n_70, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_61, n_81, n_59, n_76, n_36, n_26, n_55, n_58, n_64, n_48, n_65, n_25, n_40, n_80, n_41, n_86, n_9, n_10, n_71, n_74, n_6, n_14, n_72, n_60, n_35, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_542);

input n_52;
input n_16;
input n_1;
input n_46;
input n_18;
input n_21;
input n_3;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_77;
input n_42;
input n_8;
input n_24;
input n_54;
input n_0;
input n_32;
input n_66;
input n_85;
input n_78;
input n_84;
input n_13;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_45;
input n_34;
input n_70;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_61;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_55;
input n_58;
input n_64;
input n_48;
input n_65;
input n_25;
input n_40;
input n_80;
input n_41;
input n_86;
input n_9;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_72;
input n_60;
input n_35;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_542;

wire n_435;
wire n_91;
wire n_326;
wire n_256;
wire n_440;
wire n_507;
wire n_209;
wire n_367;
wire n_465;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_144;
wire n_365;
wire n_125;
wire n_168;
wire n_384;
wire n_297;
wire n_524;
wire n_342;
wire n_106;
wire n_358;
wire n_160;
wire n_449;
wire n_131;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_495;
wire n_350;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_108;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_389;
wire n_415;
wire n_230;
wire n_461;
wire n_141;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_114;
wire n_198;
wire n_104;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_229;
wire n_305;
wire n_532;
wire n_173;
wire n_535;
wire n_250;
wire n_372;
wire n_468;
wire n_111;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_338;
wire n_522;
wire n_466;
wire n_506;
wire n_360;
wire n_119;
wire n_235;
wire n_536;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_428;
wire n_432;
wire n_101;
wire n_167;
wire n_174;
wire n_127;
wire n_516;
wire n_153;
wire n_525;
wire n_156;
wire n_491;
wire n_145;
wire n_133;
wire n_96;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_109;
wire n_529;
wire n_445;
wire n_425;
wire n_122;
wire n_454;
wire n_218;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_112;
wire n_172;
wire n_472;
wire n_270;
wire n_239;
wire n_126;
wire n_414;
wire n_97;
wire n_490;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_93;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_460;
wire n_107;
wire n_417;
wire n_446;
wire n_498;
wire n_89;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_103;
wire n_272;
wire n_526;
wire n_185;
wire n_348;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_154;
wire n_456;
wire n_98;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_503;
wire n_152;
wire n_92;
wire n_513;
wire n_321;
wire n_331;
wire n_105;
wire n_227;
wire n_132;
wire n_406;
wire n_483;
wire n_102;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_130;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_100;
wire n_121;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_477;
wire n_533;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_243;
wire n_124;
wire n_94;
wire n_282;
wire n_436;
wire n_116;
wire n_211;
wire n_523;
wire n_117;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_505;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_537;
wire n_273;
wire n_95;
wire n_311;
wire n_403;
wire n_253;
wire n_123;
wire n_136;
wire n_249;
wire n_201;
wire n_386;
wire n_159;
wire n_157;
wire n_162;
wire n_115;
wire n_487;
wire n_128;
wire n_241;
wire n_275;
wire n_276;
wire n_441;
wire n_221;
wire n_444;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_88;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_113;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_453;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_431;
wire n_90;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_87;
wire n_195;
wire n_285;
wire n_497;
wire n_99;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_489;
wire n_205;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_151;
wire n_110;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_514;
wire n_528;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_73),
.Y(n_87)
);

NOR2xp67_ASAP7_75t_L g88 ( 
.A(n_44),
.B(n_49),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_16),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_52),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

BUFx10_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_22),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_80),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_6),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_31),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g103 ( 
.A(n_26),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_38),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_20),
.B(n_14),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_42),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_54),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_25),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_21),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_15),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_14),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_37),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

NOR2xp67_ASAP7_75t_L g116 ( 
.A(n_4),
.B(n_50),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_16),
.Y(n_120)
);

INVx4_ASAP7_75t_R g121 ( 
.A(n_7),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_51),
.Y(n_122)
);

INVxp33_ASAP7_75t_SL g123 ( 
.A(n_8),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_2),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_17),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_0),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_35),
.Y(n_128)
);

NOR2xp67_ASAP7_75t_L g129 ( 
.A(n_12),
.B(n_63),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_33),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_15),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_2),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_10),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_27),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_85),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_39),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_47),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_9),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_3),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_60),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_28),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_29),
.Y(n_145)
);

NOR2xp67_ASAP7_75t_L g146 ( 
.A(n_48),
.B(n_78),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_75),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_8),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_3),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_7),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_40),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_6),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_20),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_57),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_72),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_84),
.Y(n_157)
);

INVxp67_ASAP7_75t_SL g158 ( 
.A(n_0),
.Y(n_158)
);

INVxp33_ASAP7_75t_SL g159 ( 
.A(n_45),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_79),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_12),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_11),
.Y(n_162)
);

INVxp33_ASAP7_75t_L g163 ( 
.A(n_13),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_41),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_82),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_36),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_113),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_113),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_118),
.B(n_1),
.Y(n_171)
);

AND2x4_ASAP7_75t_L g172 ( 
.A(n_102),
.B(n_24),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_127),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_126),
.B(n_1),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_92),
.B(n_4),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_87),
.Y(n_180)
);

NOR2x1_ASAP7_75t_L g181 ( 
.A(n_92),
.B(n_43),
.Y(n_181)
);

OAI22x1_ASAP7_75t_L g182 ( 
.A1(n_149),
.A2(n_133),
.B1(n_141),
.B2(n_135),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_92),
.B(n_5),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_89),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_5),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_97),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_126),
.Y(n_188)
);

AND2x6_ASAP7_75t_L g189 ( 
.A(n_147),
.B(n_100),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_112),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_142),
.A2(n_9),
.B1(n_11),
.B2(n_13),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_101),
.B(n_17),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_120),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_100),
.B(n_18),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_134),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_111),
.B(n_150),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_125),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_133),
.Y(n_199)
);

NAND2xp33_ASAP7_75t_L g200 ( 
.A(n_106),
.B(n_18),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_109),
.B(n_19),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_153),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_141),
.A2(n_55),
.B1(n_56),
.B2(n_65),
.Y(n_203)
);

AND2x4_ASAP7_75t_L g204 ( 
.A(n_102),
.B(n_74),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_111),
.B(n_76),
.Y(n_205)
);

AND2x4_ASAP7_75t_L g206 ( 
.A(n_150),
.B(n_155),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_142),
.A2(n_77),
.B1(n_83),
.B2(n_123),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

AND2x4_ASAP7_75t_L g209 ( 
.A(n_155),
.B(n_107),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_123),
.A2(n_110),
.B1(n_91),
.B2(n_140),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_162),
.Y(n_211)
);

BUFx8_ASAP7_75t_L g212 ( 
.A(n_125),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_135),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_119),
.B(n_117),
.Y(n_214)
);

AND2x4_ASAP7_75t_L g215 ( 
.A(n_90),
.B(n_130),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_94),
.B(n_158),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_91),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_94),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_161),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_147),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_96),
.A2(n_110),
.B1(n_138),
.B2(n_140),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_93),
.B(n_131),
.Y(n_222)
);

AND2x4_ASAP7_75t_L g223 ( 
.A(n_98),
.B(n_132),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_147),
.Y(n_224)
);

NOR2x1_ASAP7_75t_L g225 ( 
.A(n_88),
.B(n_146),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_99),
.Y(n_226)
);

AND2x4_ASAP7_75t_L g227 ( 
.A(n_104),
.B(n_136),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g228 ( 
.A(n_94),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_116),
.B(n_129),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_108),
.Y(n_230)
);

NAND2xp33_ASAP7_75t_L g231 ( 
.A(n_95),
.B(n_156),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_114),
.Y(n_232)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_159),
.Y(n_233)
);

AND2x6_ASAP7_75t_L g234 ( 
.A(n_115),
.B(n_143),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_124),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_128),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_96),
.A2(n_138),
.B1(n_159),
.B2(n_105),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_139),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_192),
.A2(n_201),
.B1(n_200),
.B2(n_206),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_192),
.B(n_95),
.Y(n_240)
);

AND2x4_ASAP7_75t_L g241 ( 
.A(n_172),
.B(n_152),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_171),
.A2(n_165),
.B(n_164),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_178),
.Y(n_243)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_170),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_169),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_179),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_169),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_180),
.B(n_166),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_177),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_201),
.B(n_103),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_179),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_204),
.B(n_157),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_199),
.B(n_219),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_177),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_170),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_204),
.B(n_122),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_220),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_179),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_L g262 ( 
.A1(n_176),
.A2(n_103),
.B1(n_105),
.B2(n_160),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_137),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_229),
.B(n_137),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_214),
.B(n_144),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_220),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_224),
.Y(n_267)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_235),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_226),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_233),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_232),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_225),
.B(n_144),
.Y(n_272)
);

OR2x6_ASAP7_75t_L g273 ( 
.A(n_182),
.B(n_121),
.Y(n_273)
);

AO21x2_ASAP7_75t_L g274 ( 
.A1(n_184),
.A2(n_145),
.B(n_156),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_235),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_186),
.B(n_145),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_172),
.B(n_160),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_172),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_179),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_222),
.B(n_197),
.Y(n_280)
);

INVx6_ASAP7_75t_L g281 ( 
.A(n_212),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_219),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_194),
.B(n_236),
.Y(n_283)
);

AND2x6_ASAP7_75t_L g284 ( 
.A(n_181),
.B(n_206),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_216),
.B(n_233),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_236),
.B(n_218),
.Y(n_286)
);

OR2x6_ASAP7_75t_L g287 ( 
.A(n_228),
.B(n_191),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_200),
.A2(n_206),
.B1(n_209),
.B2(n_223),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_228),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_233),
.B(n_215),
.Y(n_290)
);

AND2x6_ASAP7_75t_L g291 ( 
.A(n_215),
.B(n_223),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_183),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_167),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_233),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_234),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_265),
.B(n_231),
.Y(n_296)
);

O2A1O1Ixp5_ASAP7_75t_L g297 ( 
.A1(n_242),
.A2(n_227),
.B(n_223),
.C(n_215),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_239),
.A2(n_205),
.B1(n_237),
.B2(n_174),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_234),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_239),
.A2(n_168),
.B1(n_173),
.B2(n_203),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_234),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_257),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_234),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_289),
.Y(n_304)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_291),
.Y(n_305)
);

NAND2xp33_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_189),
.Y(n_306)
);

AND2x6_ASAP7_75t_L g307 ( 
.A(n_278),
.B(n_227),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_246),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_269),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_246),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_271),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_R g312 ( 
.A(n_248),
.B(n_231),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_240),
.A2(n_210),
.B1(n_207),
.B2(n_221),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_278),
.B(n_227),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_288),
.B(n_209),
.Y(n_315)
);

AND2x4_ASAP7_75t_L g316 ( 
.A(n_241),
.B(n_196),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_293),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_257),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_286),
.B(n_209),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_275),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_266),
.Y(n_321)
);

AND3x1_ASAP7_75t_L g322 ( 
.A(n_283),
.B(n_193),
.C(n_211),
.Y(n_322)
);

AND2x4_ASAP7_75t_L g323 ( 
.A(n_241),
.B(n_195),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g324 ( 
.A1(n_288),
.A2(n_190),
.B1(n_198),
.B2(n_213),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_252),
.B(n_189),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_263),
.B(n_185),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_286),
.B(n_213),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_256),
.B(n_189),
.Y(n_328)
);

A2O1A1Ixp33_ASAP7_75t_L g329 ( 
.A1(n_263),
.A2(n_187),
.B(n_202),
.C(n_208),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_284),
.B(n_217),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_284),
.B(n_175),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_290),
.B(n_285),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_285),
.B(n_188),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_266),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_274),
.B(n_277),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_267),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_250),
.B(n_262),
.Y(n_337)
);

A2O1A1Ixp33_ASAP7_75t_L g338 ( 
.A1(n_296),
.A2(n_277),
.B(n_276),
.C(n_253),
.Y(n_338)
);

A2O1A1Ixp33_ASAP7_75t_L g339 ( 
.A1(n_296),
.A2(n_276),
.B(n_264),
.C(n_272),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_315),
.B(n_270),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_316),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_326),
.B(n_282),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_302),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_315),
.B(n_270),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_294),
.B(n_273),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_326),
.B(n_264),
.Y(n_346)
);

O2A1O1Ixp33_ASAP7_75t_L g347 ( 
.A1(n_298),
.A2(n_259),
.B(n_261),
.C(n_260),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_302),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_R g349 ( 
.A(n_304),
.B(n_281),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_318),
.Y(n_350)
);

CKINVDCx11_ASAP7_75t_R g351 ( 
.A(n_300),
.Y(n_351)
);

A2O1A1Ixp33_ASAP7_75t_L g352 ( 
.A1(n_297),
.A2(n_335),
.B(n_295),
.C(n_337),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_314),
.A2(n_268),
.B(n_258),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_319),
.B(n_273),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_R g355 ( 
.A(n_306),
.B(n_281),
.Y(n_355)
);

O2A1O1Ixp33_ASAP7_75t_L g356 ( 
.A1(n_329),
.A2(n_243),
.B(n_255),
.C(n_245),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_316),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_332),
.A2(n_268),
.B(n_246),
.Y(n_358)
);

O2A1O1Ixp5_ASAP7_75t_SL g359 ( 
.A1(n_320),
.A2(n_247),
.B(n_249),
.C(n_244),
.Y(n_359)
);

BUFx8_ASAP7_75t_L g360 ( 
.A(n_309),
.Y(n_360)
);

OR2x6_ASAP7_75t_SL g361 ( 
.A(n_331),
.B(n_287),
.Y(n_361)
);

AND2x4_ASAP7_75t_L g362 ( 
.A(n_323),
.B(n_292),
.Y(n_362)
);

NOR2xp67_ASAP7_75t_L g363 ( 
.A(n_305),
.B(n_254),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_327),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_307),
.Y(n_365)
);

A2O1A1Ixp33_ASAP7_75t_L g366 ( 
.A1(n_313),
.A2(n_325),
.B(n_328),
.C(n_311),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_318),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_299),
.A2(n_251),
.B(n_258),
.Y(n_368)
);

INVx3_ASAP7_75t_SL g369 ( 
.A(n_317),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_321),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_301),
.A2(n_279),
.B(n_303),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_330),
.Y(n_372)
);

NAND3xp33_ASAP7_75t_SL g373 ( 
.A(n_312),
.B(n_324),
.C(n_322),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_305),
.A2(n_321),
.B1(n_334),
.B2(n_336),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_307),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_305),
.A2(n_334),
.B(n_336),
.Y(n_376)
);

NOR2xp67_ASAP7_75t_L g377 ( 
.A(n_308),
.B(n_310),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_310),
.B(n_296),
.Y(n_378)
);

NAND2x1p5_ASAP7_75t_L g379 ( 
.A(n_310),
.B(n_315),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_310),
.B(n_296),
.Y(n_380)
);

AO21x1_ASAP7_75t_L g381 ( 
.A1(n_335),
.A2(n_296),
.B(n_298),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_296),
.A2(n_335),
.B1(n_298),
.B2(n_337),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_315),
.A2(n_314),
.B(n_332),
.Y(n_383)
);

A2O1A1Ixp33_ASAP7_75t_L g384 ( 
.A1(n_296),
.A2(n_242),
.B(n_326),
.C(n_297),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_315),
.A2(n_314),
.B(n_332),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_315),
.A2(n_314),
.B(n_332),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g387 ( 
.A(n_327),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_304),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_296),
.B(n_315),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g390 ( 
.A(n_364),
.B(n_342),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_382),
.B(n_380),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_343),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_348),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_341),
.B(n_357),
.Y(n_394)
);

CKINVDCx11_ASAP7_75t_R g395 ( 
.A(n_361),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_L g396 ( 
.A1(n_381),
.A2(n_351),
.B1(n_373),
.B2(n_387),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_338),
.B(n_372),
.Y(n_397)
);

A2O1A1Ixp33_ASAP7_75t_L g398 ( 
.A1(n_384),
.A2(n_339),
.B(n_352),
.C(n_385),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_350),
.Y(n_399)
);

NAND2x1p5_ASAP7_75t_L g400 ( 
.A(n_365),
.B(n_375),
.Y(n_400)
);

A2O1A1Ixp33_ASAP7_75t_L g401 ( 
.A1(n_383),
.A2(n_386),
.B(n_366),
.C(n_347),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_378),
.A2(n_354),
.B1(n_345),
.B2(n_379),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_367),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_370),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_340),
.A2(n_344),
.B(n_371),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_369),
.B(n_341),
.Y(n_406)
);

INVxp33_ASAP7_75t_SL g407 ( 
.A(n_388),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_365),
.B(n_341),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_356),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_357),
.Y(n_410)
);

OAI21x1_ASAP7_75t_L g411 ( 
.A1(n_368),
.A2(n_376),
.B(n_358),
.Y(n_411)
);

OAI21x1_ASAP7_75t_L g412 ( 
.A1(n_359),
.A2(n_353),
.B(n_374),
.Y(n_412)
);

INVx6_ASAP7_75t_L g413 ( 
.A(n_360),
.Y(n_413)
);

AO31x2_ASAP7_75t_L g414 ( 
.A1(n_377),
.A2(n_363),
.A3(n_355),
.B(n_360),
.Y(n_414)
);

CKINVDCx8_ASAP7_75t_R g415 ( 
.A(n_349),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_377),
.A2(n_221),
.B1(n_188),
.B2(n_210),
.Y(n_416)
);

AO31x2_ASAP7_75t_L g417 ( 
.A1(n_363),
.A2(n_381),
.A3(n_352),
.B(n_384),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_341),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_L g419 ( 
.A1(n_381),
.A2(n_382),
.B1(n_296),
.B2(n_337),
.Y(n_419)
);

O2A1O1Ixp33_ASAP7_75t_L g420 ( 
.A1(n_346),
.A2(n_338),
.B(n_384),
.C(n_339),
.Y(n_420)
);

AO32x2_ASAP7_75t_L g421 ( 
.A1(n_381),
.A2(n_298),
.A3(n_300),
.B1(n_374),
.B2(n_387),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_381),
.A2(n_382),
.B1(n_389),
.B2(n_351),
.Y(n_422)
);

AO32x2_ASAP7_75t_L g423 ( 
.A1(n_381),
.A2(n_298),
.A3(n_300),
.B1(n_374),
.B2(n_387),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_389),
.A2(n_315),
.B(n_383),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_346),
.B(n_333),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_388),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_346),
.B(n_217),
.Y(n_427)
);

O2A1O1Ixp33_ASAP7_75t_L g428 ( 
.A1(n_346),
.A2(n_338),
.B(n_384),
.C(n_339),
.Y(n_428)
);

O2A1O1Ixp5_ASAP7_75t_L g429 ( 
.A1(n_378),
.A2(n_296),
.B(n_381),
.C(n_384),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_342),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_389),
.A2(n_315),
.B(n_383),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_341),
.B(n_357),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_343),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_342),
.Y(n_434)
);

AO22x2_ASAP7_75t_L g435 ( 
.A1(n_373),
.A2(n_298),
.B1(n_337),
.B2(n_346),
.Y(n_435)
);

INVx2_ASAP7_75t_SL g436 ( 
.A(n_362),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_346),
.B(n_217),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_382),
.A2(n_239),
.B1(n_346),
.B2(n_384),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_388),
.Y(n_439)
);

A2O1A1Ixp33_ASAP7_75t_L g440 ( 
.A1(n_420),
.A2(n_428),
.B(n_422),
.C(n_419),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_409),
.Y(n_441)
);

CKINVDCx6p67_ASAP7_75t_R g442 ( 
.A(n_426),
.Y(n_442)
);

OA21x2_ASAP7_75t_L g443 ( 
.A1(n_398),
.A2(n_429),
.B(n_401),
.Y(n_443)
);

OAI21x1_ASAP7_75t_SL g444 ( 
.A1(n_438),
.A2(n_424),
.B(n_431),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_392),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_393),
.Y(n_446)
);

CKINVDCx11_ASAP7_75t_R g447 ( 
.A(n_415),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_425),
.B(n_391),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_394),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_407),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_391),
.A2(n_397),
.B(n_405),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_435),
.B(n_422),
.Y(n_452)
);

A2O1A1Ixp33_ASAP7_75t_L g453 ( 
.A1(n_427),
.A2(n_437),
.B(n_402),
.C(n_396),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_399),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_403),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_421),
.B(n_423),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_404),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_433),
.Y(n_458)
);

AO21x2_ASAP7_75t_L g459 ( 
.A1(n_412),
.A2(n_402),
.B(n_411),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_406),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_430),
.B(n_434),
.Y(n_461)
);

OAI222xp33_ASAP7_75t_L g462 ( 
.A1(n_390),
.A2(n_418),
.B1(n_394),
.B2(n_432),
.C1(n_416),
.C2(n_436),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_421),
.B(n_423),
.Y(n_463)
);

OAI322xp33_ASAP7_75t_L g464 ( 
.A1(n_416),
.A2(n_408),
.A3(n_423),
.B1(n_421),
.B2(n_418),
.C1(n_410),
.C2(n_400),
.Y(n_464)
);

AOI22xp33_ASAP7_75t_SL g465 ( 
.A1(n_439),
.A2(n_432),
.B1(n_410),
.B2(n_413),
.Y(n_465)
);

BUFx4f_ASAP7_75t_SL g466 ( 
.A(n_413),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_395),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_417),
.Y(n_468)
);

BUFx8_ASAP7_75t_L g469 ( 
.A(n_414),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_435),
.A2(n_351),
.B1(n_381),
.B2(n_296),
.Y(n_470)
);

OR2x6_ASAP7_75t_L g471 ( 
.A(n_444),
.B(n_451),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_441),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g473 ( 
.A(n_460),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_448),
.B(n_470),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_449),
.B(n_455),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_452),
.B(n_440),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_468),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_453),
.B(n_463),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_456),
.B(n_463),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_456),
.B(n_443),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_469),
.Y(n_481)
);

OA21x2_ASAP7_75t_L g482 ( 
.A1(n_462),
.A2(n_458),
.B(n_445),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_461),
.A2(n_465),
.B1(n_446),
.B2(n_458),
.Y(n_483)
);

AO21x2_ASAP7_75t_L g484 ( 
.A1(n_459),
.A2(n_457),
.B(n_446),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_454),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_477),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_474),
.B(n_450),
.Y(n_487)
);

AOI211xp5_ASAP7_75t_L g488 ( 
.A1(n_474),
.A2(n_464),
.B(n_450),
.C(n_454),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_476),
.B(n_442),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_481),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_477),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_475),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_476),
.B(n_442),
.Y(n_493)
);

OR2x2_ASAP7_75t_SL g494 ( 
.A(n_476),
.B(n_466),
.Y(n_494)
);

OR2x6_ASAP7_75t_L g495 ( 
.A(n_471),
.B(n_469),
.Y(n_495)
);

NOR2xp67_ASAP7_75t_L g496 ( 
.A(n_483),
.B(n_469),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_473),
.B(n_447),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_490),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_488),
.B(n_478),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_494),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_486),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_492),
.B(n_479),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_495),
.B(n_480),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_495),
.B(n_484),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_491),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_488),
.B(n_478),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_505),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_503),
.B(n_495),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_503),
.B(n_495),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_501),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_502),
.B(n_495),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_502),
.B(n_506),
.Y(n_512)
);

NAND2x1_ASAP7_75t_L g513 ( 
.A(n_505),
.B(n_496),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_511),
.B(n_504),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_510),
.Y(n_515)
);

AOI21xp33_ASAP7_75t_L g516 ( 
.A1(n_513),
.A2(n_489),
.B(n_493),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_507),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_511),
.B(n_504),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_507),
.Y(n_519)
);

NAND2xp33_ASAP7_75t_SL g520 ( 
.A(n_512),
.B(n_506),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_508),
.A2(n_494),
.B1(n_496),
.B2(n_500),
.Y(n_521)
);

OAI21xp33_ASAP7_75t_L g522 ( 
.A1(n_516),
.A2(n_487),
.B(n_499),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_519),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_515),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_520),
.B(n_500),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_520),
.A2(n_471),
.B(n_499),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_525),
.B(n_518),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_526),
.B(n_518),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_522),
.B(n_497),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_529),
.A2(n_525),
.B(n_521),
.Y(n_530)
);

AOI211xp5_ASAP7_75t_L g531 ( 
.A1(n_528),
.A2(n_500),
.B(n_498),
.C(n_524),
.Y(n_531)
);

AOI221xp5_ASAP7_75t_L g532 ( 
.A1(n_530),
.A2(n_527),
.B1(n_498),
.B2(n_523),
.C(n_517),
.Y(n_532)
);

AOI221xp5_ASAP7_75t_L g533 ( 
.A1(n_531),
.A2(n_473),
.B1(n_509),
.B2(n_508),
.C(n_514),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_467),
.Y(n_534)
);

NOR3xp33_ASAP7_75t_L g535 ( 
.A(n_532),
.B(n_490),
.C(n_483),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_534),
.B(n_509),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_536),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_537),
.A2(n_535),
.B(n_481),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_538),
.A2(n_519),
.B1(n_481),
.B2(n_504),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_539),
.B(n_514),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_540),
.A2(n_469),
.B1(n_504),
.B2(n_472),
.Y(n_541)
);

AOI21xp33_ASAP7_75t_SL g542 ( 
.A1(n_541),
.A2(n_485),
.B(n_482),
.Y(n_542)
);


endmodule