module real_jpeg_30957_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_663, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_663;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_611;
wire n_221;
wire n_489;
wire n_393;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_653;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_497;
wire n_633;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_604;
wire n_420;
wire n_357;
wire n_431;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_586;
wire n_572;
wire n_548;
wire n_319;
wire n_487;
wire n_93;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_602;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_636;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_0),
.Y(n_129)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_0),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_0),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_0),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_1),
.Y(n_174)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_1),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_2),
.A2(n_160),
.B1(n_161),
.B2(n_166),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_2),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_2),
.A2(n_160),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_2),
.A2(n_160),
.B1(n_292),
.B2(n_296),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_2),
.A2(n_160),
.B1(n_403),
.B2(n_406),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_3),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_3),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_L g259 ( 
.A1(n_3),
.A2(n_186),
.B1(n_260),
.B2(n_262),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_3),
.A2(n_186),
.B1(n_372),
.B2(n_375),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_3),
.A2(n_186),
.B1(n_463),
.B2(n_466),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_4),
.A2(n_113),
.B1(n_120),
.B2(n_121),
.Y(n_112)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_4),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_4),
.A2(n_120),
.B1(n_146),
.B2(n_151),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_4),
.A2(n_120),
.B1(n_284),
.B2(n_286),
.Y(n_283)
);

AO22x1_ASAP7_75t_L g628 ( 
.A1(n_4),
.A2(n_120),
.B1(n_629),
.B2(n_631),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_5),
.A2(n_239),
.B1(n_240),
.B2(n_243),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_5),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_5),
.A2(n_239),
.B1(n_341),
.B2(n_345),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g433 ( 
.A1(n_5),
.A2(n_239),
.B1(n_434),
.B2(n_437),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_SL g533 ( 
.A1(n_5),
.A2(n_239),
.B1(n_534),
.B2(n_536),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_6),
.A2(n_72),
.B1(n_77),
.B2(n_78),
.Y(n_71)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_6),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_6),
.A2(n_77),
.B1(n_138),
.B2(n_141),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_6),
.A2(n_77),
.B1(n_637),
.B2(n_638),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_7),
.B(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_7),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_7),
.B(n_170),
.Y(n_408)
);

OAI32xp33_ASAP7_75t_L g441 ( 
.A1(n_7),
.A2(n_442),
.A3(n_445),
.B1(n_447),
.B2(n_452),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_SL g483 ( 
.A1(n_7),
.A2(n_368),
.B1(n_484),
.B2(n_487),
.Y(n_483)
);

OAI21xp33_ASAP7_75t_L g515 ( 
.A1(n_7),
.A2(n_220),
.B(n_516),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_8),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_8),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_8),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_9),
.Y(n_88)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_9),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_10),
.Y(n_133)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_10),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_11),
.A2(n_103),
.B1(n_108),
.B2(n_109),
.Y(n_102)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_11),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_11),
.A2(n_108),
.B1(n_206),
.B2(n_209),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g328 ( 
.A1(n_11),
.A2(n_108),
.B1(n_329),
.B2(n_332),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g601 ( 
.A1(n_11),
.A2(n_108),
.B1(n_317),
.B2(n_602),
.Y(n_601)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_13),
.B(n_646),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_13),
.B(n_645),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_14),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_15),
.A2(n_271),
.B1(n_272),
.B2(n_278),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_15),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_15),
.A2(n_271),
.B1(n_383),
.B2(n_389),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_SL g489 ( 
.A1(n_15),
.A2(n_271),
.B1(n_490),
.B2(n_492),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_15),
.A2(n_271),
.B1(n_504),
.B2(n_508),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_16),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_16),
.Y(n_107)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_16),
.Y(n_119)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_17),
.A2(n_60),
.B1(n_215),
.B2(n_218),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_17),
.A2(n_60),
.B1(n_611),
.B2(n_614),
.Y(n_610)
);

INVxp33_ASAP7_75t_L g646 ( 
.A(n_18),
.Y(n_646)
);

OAI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.A3(n_592),
.B1(n_643),
.B2(n_654),
.C(n_658),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2x1_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_422),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_347),
.B(n_418),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_25),
.B(n_589),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_246),
.B(n_297),
.Y(n_25)
);

NOR2x1_ASAP7_75t_L g420 ( 
.A(n_26),
.B(n_246),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_26),
.B(n_246),
.Y(n_421)
);

XOR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_202),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_124),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g653 ( 
.A(n_28),
.Y(n_653)
);

OA21x2_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_83),
.B(n_123),
.Y(n_28)
);

NAND2x1_ASAP7_75t_L g123 ( 
.A(n_29),
.B(n_83),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_58),
.B1(n_71),
.B2(n_81),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_30),
.A2(n_371),
.B1(n_377),
.B2(n_378),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_30),
.B(n_566),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_30),
.A2(n_81),
.B1(n_371),
.B2(n_576),
.Y(n_575)
);

OA21x2_ASAP7_75t_L g607 ( 
.A1(n_30),
.A2(n_71),
.B(n_81),
.Y(n_607)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_31),
.A2(n_59),
.B1(n_145),
.B2(n_154),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_31),
.A2(n_145),
.B1(n_154),
.B2(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_31),
.A2(n_154),
.B1(n_205),
.B2(n_291),
.Y(n_290)
);

OAI21xp33_ASAP7_75t_SL g432 ( 
.A1(n_31),
.A2(n_433),
.B(n_439),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_31),
.A2(n_154),
.B1(n_433),
.B2(n_489),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_46),
.Y(n_31)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

OAI22x1_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_36),
.B1(n_40),
.B2(n_43),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g510 ( 
.A(n_34),
.Y(n_510)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_39),
.Y(n_551)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_41),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_43),
.Y(n_467)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_45),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_45),
.Y(n_465)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_45),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_51),
.B1(n_52),
.B2(n_55),
.Y(n_46)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_47),
.Y(n_446)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_48),
.Y(n_376)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_54),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_54),
.Y(n_438)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B(n_65),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g491 ( 
.A(n_64),
.Y(n_491)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_69),
.Y(n_212)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_69),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_70),
.Y(n_374)
);

BUFx5_ASAP7_75t_L g557 ( 
.A(n_70),
.Y(n_557)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_76),
.Y(n_208)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_76),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_76),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_80),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_81),
.B(n_371),
.Y(n_439)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_82),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_82),
.B(n_368),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_102),
.B1(n_111),
.B2(n_112),
.Y(n_83)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_84),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_84),
.A2(n_380),
.B1(n_381),
.B2(n_382),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_84),
.B(n_414),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_84),
.A2(n_112),
.B1(n_381),
.B2(n_610),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_84),
.A2(n_111),
.B1(n_610),
.B2(n_636),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_92),
.Y(n_84)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_88),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_89),
.A2(n_93),
.B1(n_97),
.B2(n_101),
.Y(n_92)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_93),
.Y(n_345)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

INVx4_ASAP7_75t_L g614 ( 
.A(n_95),
.Y(n_614)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_102),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_105),
.Y(n_261)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_106),
.Y(n_231)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_107),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_107),
.Y(n_182)
);

BUFx4f_ASAP7_75t_L g309 ( 
.A(n_109),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_110),
.Y(n_228)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_110),
.Y(n_344)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_110),
.Y(n_613)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_111),
.Y(n_232)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_111),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_111),
.B(n_259),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_111),
.B(n_382),
.Y(n_411)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_118),
.Y(n_390)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_118),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_119),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_119),
.Y(n_388)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_123),
.Y(n_617)
);

XOR2xp5_ASAP7_75t_L g650 ( 
.A(n_123),
.B(n_598),
.Y(n_650)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_124),
.Y(n_652)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_155),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g618 ( 
.A1(n_125),
.A2(n_199),
.B(n_619),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_144),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_126),
.Y(n_252)
);

OA21x2_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_130),
.B(n_137),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_127),
.Y(n_460)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_130),
.A2(n_137),
.B(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_130),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_130),
.A2(n_223),
.B1(n_283),
.B2(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_130),
.B(n_462),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_130),
.A2(n_288),
.B1(n_531),
.B2(n_532),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.Y(n_130)
);

BUFx4f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_133),
.Y(n_217)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_133),
.Y(n_285)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_133),
.Y(n_527)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_134),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_136),
.Y(n_513)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_137),
.Y(n_221)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_140),
.Y(n_219)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_142),
.Y(n_286)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_142),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_143),
.Y(n_331)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_143),
.Y(n_405)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_143),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_144),
.A2(n_198),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_144),
.Y(n_253)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_SL g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx4f_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_154),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_198),
.B2(n_199),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_157),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_183),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_170),
.Y(n_158)
);

AO22x1_ASAP7_75t_L g599 ( 
.A1(n_159),
.A2(n_600),
.B1(n_601),
.B2(n_604),
.Y(n_599)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_163),
.A2(n_167),
.B1(n_192),
.B2(n_194),
.Y(n_191)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_164),
.Y(n_242)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_165),
.Y(n_245)
);

INVx6_ASAP7_75t_L g315 ( 
.A(n_165),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_165),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx4_ASAP7_75t_SL g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_170),
.B(n_184),
.Y(n_236)
);

AO22x1_ASAP7_75t_L g269 ( 
.A1(n_170),
.A2(n_190),
.B1(n_238),
.B2(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_170),
.B(n_270),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_170),
.Y(n_604)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_175),
.B1(n_177),
.B2(n_180),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_174),
.Y(n_179)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_174),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_174),
.Y(n_324)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_176),
.Y(n_486)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_180),
.Y(n_321)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_182),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_182),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_183),
.B(n_337),
.Y(n_336)
);

NAND2x1_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_190),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g603 ( 
.A(n_189),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_SL g237 ( 
.A(n_190),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_190),
.B(n_363),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_190),
.Y(n_600)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_193),
.Y(n_311)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_201),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_201),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_R g651 ( 
.A(n_202),
.B(n_652),
.C(n_653),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_224),
.C(n_234),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_203),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_213),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_204),
.B(n_213),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_208),
.Y(n_296)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_214),
.A2(n_220),
.B1(n_282),
.B2(n_287),
.Y(n_281)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_217),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

OAI22x1_ASAP7_75t_L g397 ( 
.A1(n_220),
.A2(n_328),
.B1(n_398),
.B2(n_402),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g573 ( 
.A1(n_220),
.A2(n_516),
.B(n_533),
.Y(n_573)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_224),
.A2(n_234),
.B1(n_235),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_224),
.Y(n_249)
);

OA22x2_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_232),
.B2(n_233),
.Y(n_224)
);

OAI22x1_ASAP7_75t_L g257 ( 
.A1(n_225),
.A2(n_226),
.B1(n_258),
.B2(n_267),
.Y(n_257)
);

OA21x2_ASAP7_75t_L g339 ( 
.A1(n_225),
.A2(n_340),
.B(n_346),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_225),
.A2(n_346),
.B(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_236),
.B(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_245),
.Y(n_279)
);

MAJx2_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_250),
.C(n_254),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_247),
.B(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_251),
.B(n_255),
.Y(n_299)
);

INVxp33_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_268),
.C(n_280),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_257),
.B(n_269),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_258),
.Y(n_414)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_263),
.Y(n_454)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_267),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_267),
.B(n_368),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_275),
.Y(n_632)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_303),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_290),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_281),
.B(n_290),
.Y(n_358)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx5_ASAP7_75t_L g524 ( 
.A(n_289),
.Y(n_524)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_291),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_298),
.B(n_300),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_304),
.C(n_305),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_301),
.A2(n_302),
.B1(n_304),
.B2(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_304),
.Y(n_352)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_305),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_335),
.C(n_338),
.Y(n_305)
);

XNOR2x1_ASAP7_75t_SL g354 ( 
.A(n_306),
.B(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_325),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_307),
.A2(n_308),
.B1(n_325),
.B2(n_326),
.Y(n_415)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

AOI32xp33_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_310),
.A3(n_312),
.B1(n_316),
.B2(n_319),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_315),
.Y(n_367)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_315),
.Y(n_630)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_316),
.Y(n_369)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NAND2xp33_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_322),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_333),
.Y(n_538)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_335),
.A2(n_336),
.B1(n_339),
.B2(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_339),
.Y(n_356)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_340),
.Y(n_380)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_353),
.C(n_391),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g589 ( 
.A1(n_349),
.A2(n_590),
.B(n_591),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_353),
.Y(n_590)
);

MAJx2_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_357),
.C(n_359),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_354),
.B(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_358),
.B(n_360),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

MAJx2_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_370),
.C(n_379),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_361),
.B(n_394),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_364),
.A2(n_368),
.B(n_369),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_368),
.B(n_448),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_368),
.B(n_524),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_368),
.B(n_554),
.Y(n_553)
);

OAI21xp33_ASAP7_75t_SL g566 ( 
.A1(n_368),
.A2(n_553),
.B(n_567),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_370),
.B(n_379),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_374),
.Y(n_496)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_416),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_392),
.B(n_416),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_395),
.C(n_415),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_393),
.B(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_396),
.A2(n_415),
.B1(n_470),
.B2(n_471),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_408),
.B1(n_409),
.B2(n_412),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_397),
.B(n_408),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_397),
.B(n_408),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_397),
.A2(n_408),
.B1(n_409),
.B2(n_412),
.Y(n_472)
);

INVx3_ASAP7_75t_SL g398 ( 
.A(n_399),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_402),
.A2(n_460),
.B(n_461),
.Y(n_459)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_411),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_411),
.B(n_413),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_415),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_419),
.A2(n_420),
.B(n_421),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_588),
.Y(n_422)
);

OAI21x1_ASAP7_75t_L g423 ( 
.A1(n_424),
.A2(n_473),
.B(n_586),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_468),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_426),
.B(n_587),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_431),
.C(n_440),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_428),
.B(n_476),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_431),
.A2(n_432),
.B1(n_440),
.B2(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx2_ASAP7_75t_SL g434 ( 
.A(n_435),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_436),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_439),
.B(n_565),
.Y(n_564)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_440),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_459),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_441),
.B(n_459),
.Y(n_480)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_451),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_455),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_461),
.A2(n_503),
.B(n_511),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_462),
.B(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_468),
.Y(n_587)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_474),
.A2(n_497),
.B(n_585),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_475),
.B(n_478),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_475),
.B(n_478),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_481),
.C(n_488),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_480),
.B(n_571),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_482),
.B(n_488),
.Y(n_571)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_489),
.Y(n_576)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

OAI321xp33_ASAP7_75t_L g497 ( 
.A1(n_498),
.A2(n_569),
.A3(n_578),
.B1(n_583),
.B2(n_584),
.C(n_663),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_499),
.A2(n_529),
.B(n_568),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_500),
.A2(n_514),
.B(n_528),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_502),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_501),
.B(n_502),
.Y(n_528)
);

INVxp33_ASAP7_75t_L g531 ( 
.A(n_503),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

BUFx2_ASAP7_75t_SL g506 ( 
.A(n_507),
.Y(n_506)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_515),
.B(n_522),
.Y(n_514)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_523),
.B(n_525),
.Y(n_522)
);

INVx5_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_530),
.B(n_539),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_530),
.B(n_539),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_564),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_540),
.B(n_564),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_541),
.A2(n_552),
.B1(n_558),
.B2(n_563),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_542),
.B(n_546),
.Y(n_541)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_542),
.Y(n_563)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

INVx6_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_559),
.B(n_561),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_560),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

AND2x2_ASAP7_75t_SL g569 ( 
.A(n_570),
.B(n_572),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g584 ( 
.A(n_570),
.B(n_572),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_573),
.B(n_574),
.C(n_577),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_573),
.B(n_581),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_574),
.A2(n_575),
.B1(n_577),
.B2(n_582),
.Y(n_581)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_577),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_579),
.B(n_580),
.Y(n_578)
);

NAND2xp33_ASAP7_75t_SL g583 ( 
.A(n_579),
.B(n_580),
.Y(n_583)
);

NAND3xp33_ASAP7_75t_L g654 ( 
.A(n_592),
.B(n_644),
.C(n_655),
.Y(n_654)
);

AOI221xp5_ASAP7_75t_L g658 ( 
.A1(n_592),
.A2(n_593),
.B1(n_659),
.B2(n_660),
.C(n_661),
.Y(n_658)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_593),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_594),
.B(n_642),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_595),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_596),
.B(n_621),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_596),
.B(n_621),
.Y(n_642)
);

OAI21xp5_ASAP7_75t_L g596 ( 
.A1(n_597),
.A2(n_616),
.B(n_620),
.Y(n_596)
);

INVxp33_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

XNOR2x1_ASAP7_75t_L g598 ( 
.A(n_599),
.B(n_605),
.Y(n_598)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_599),
.Y(n_623)
);

AO22x1_ASAP7_75t_SL g627 ( 
.A1(n_600),
.A2(n_601),
.B1(n_604),
.B2(n_628),
.Y(n_627)
);

INVx5_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

AOI21x1_ASAP7_75t_L g605 ( 
.A1(n_606),
.A2(n_608),
.B(n_615),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_606),
.A2(n_607),
.B1(n_634),
.B2(n_635),
.Y(n_633)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_607),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_607),
.B(n_609),
.Y(n_615)
);

MAJx2_ASAP7_75t_L g622 ( 
.A(n_607),
.B(n_608),
.C(n_623),
.Y(n_622)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_609),
.Y(n_608)
);

INVx1_ASAP7_75t_SL g611 ( 
.A(n_612),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_613),
.Y(n_612)
);

INVx3_ASAP7_75t_SL g637 ( 
.A(n_614),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_617),
.B(n_618),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_617),
.B(n_618),
.Y(n_620)
);

XNOR2xp5_ASAP7_75t_L g649 ( 
.A(n_618),
.B(n_650),
.Y(n_649)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_622),
.B(n_624),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_623),
.B(n_625),
.Y(n_624)
);

XOR2xp5_ASAP7_75t_L g625 ( 
.A(n_626),
.B(n_633),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_627),
.Y(n_626)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_630),
.Y(n_629)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_632),
.Y(n_631)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_635),
.Y(n_634)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_639),
.Y(n_638)
);

HB1xp67_ASAP7_75t_L g639 ( 
.A(n_640),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_641),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_643),
.B(n_655),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_644),
.B(n_647),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_645),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_645),
.B(n_647),
.Y(n_660)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_648),
.Y(n_647)
);

NOR2xp67_ASAP7_75t_L g648 ( 
.A(n_649),
.B(n_651),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_649),
.B(n_651),
.Y(n_657)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_656),
.Y(n_655)
);

INVxp33_ASAP7_75t_SL g656 ( 
.A(n_657),
.Y(n_656)
);


endmodule