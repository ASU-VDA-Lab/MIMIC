module real_jpeg_32702_n_2 (n_14, n_1, n_0, n_2);

input n_14;
input n_1;
input n_0;

output n_2;

wire n_5;
wire n_4;
wire n_8;
wire n_12;
wire n_11;
wire n_6;
wire n_7;
wire n_3;
wire n_10;
wire n_9;

INVxp67_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_4),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

AO21x1_ASAP7_75t_L g2 ( 
.A1(n_3),
.A2(n_10),
.B(n_11),
.Y(n_2)
);

INVxp33_ASAP7_75t_L g3 ( 
.A(n_4),
.Y(n_3)
);

NOR2xp33_ASAP7_75t_L g4 ( 
.A(n_5),
.B(n_6),
.Y(n_4)
);

INVx5_ASAP7_75t_L g6 ( 
.A(n_7),
.Y(n_6)
);

INVx3_ASAP7_75t_L g7 ( 
.A(n_8),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_9),
.Y(n_8)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g5 ( 
.A(n_14),
.Y(n_5)
);


endmodule