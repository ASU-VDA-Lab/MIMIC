module fake_jpeg_15703_n_289 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_289);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_12),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_33),
.B(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx12f_ASAP7_75t_SL g36 ( 
.A(n_19),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_38),
.Y(n_46)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_15),
.Y(n_40)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_27),
.B1(n_18),
.B2(n_16),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_44),
.A2(n_51),
.B1(n_20),
.B2(n_22),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_14),
.B1(n_16),
.B2(n_18),
.Y(n_51)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_33),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_56),
.B(n_59),
.Y(n_78)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_14),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_56),
.A2(n_37),
.B1(n_34),
.B2(n_40),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_60),
.A2(n_54),
.B1(n_43),
.B2(n_30),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_62),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_51),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_84),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_46),
.A2(n_39),
.B(n_38),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_75),
.B(n_39),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_40),
.B1(n_37),
.B2(n_34),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_68),
.A2(n_79),
.B1(n_80),
.B2(n_48),
.Y(n_97)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

BUFx8_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_41),
.A2(n_27),
.B1(n_22),
.B2(n_18),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_74),
.A2(n_81),
.B(n_83),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_27),
.B1(n_22),
.B2(n_40),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_37),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_55),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_27),
.B1(n_30),
.B2(n_40),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_49),
.A2(n_30),
.B1(n_35),
.B2(n_32),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_50),
.A2(n_16),
.B1(n_26),
.B2(n_17),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_50),
.A2(n_17),
.B1(n_26),
.B2(n_23),
.Y(n_83)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_100),
.Y(n_114)
);

HAxp5_ASAP7_75t_SL g121 ( 
.A(n_86),
.B(n_71),
.CON(n_121),
.SN(n_121)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

XNOR2x1_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_66),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_103),
.C(n_107),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_25),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_102),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_23),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_94),
.B(n_96),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_62),
.B(n_26),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_97),
.A2(n_65),
.B1(n_35),
.B2(n_32),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_53),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_101),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_75),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_25),
.Y(n_104)
);

INVxp33_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

MAJx2_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_48),
.C(n_30),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_108),
.A2(n_73),
.B1(n_67),
.B2(n_80),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_84),
.A2(n_32),
.B1(n_31),
.B2(n_35),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_109),
.A2(n_73),
.B1(n_67),
.B2(n_70),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_60),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_84),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_111),
.A2(n_102),
.B(n_96),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_113),
.A2(n_117),
.B1(n_126),
.B2(n_133),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_106),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_134),
.Y(n_141)
);

OAI32xp33_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_65),
.A3(n_71),
.B1(n_61),
.B2(n_17),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_109),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_71),
.Y(n_119)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_110),
.A2(n_73),
.B1(n_72),
.B2(n_70),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_129),
.B1(n_131),
.B2(n_132),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_93),
.B(n_95),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_70),
.Y(n_124)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_65),
.B1(n_57),
.B2(n_52),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_100),
.A2(n_32),
.B1(n_35),
.B2(n_47),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_105),
.A2(n_57),
.B1(n_52),
.B2(n_47),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_87),
.A2(n_10),
.B1(n_13),
.B2(n_11),
.Y(n_133)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_88),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_105),
.A2(n_28),
.B1(n_21),
.B2(n_42),
.Y(n_135)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_107),
.C(n_106),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_137),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_130),
.B(n_94),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_139),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_130),
.B(n_97),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_119),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_145),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_106),
.C(n_108),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_144),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_99),
.C(n_95),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_115),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_99),
.Y(n_146)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_116),
.Y(n_147)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_148),
.A2(n_151),
.B1(n_156),
.B2(n_155),
.Y(n_161)
);

AND2x6_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_93),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_149),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_124),
.Y(n_150)
);

XOR2x2_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_127),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_111),
.A2(n_90),
.B1(n_25),
.B2(n_28),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_154),
.A2(n_148),
.B1(n_123),
.B2(n_141),
.Y(n_172)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_112),
.Y(n_157)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_125),
.A2(n_89),
.B(n_19),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_29),
.Y(n_180)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_115),
.Y(n_160)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_161),
.A2(n_167),
.B1(n_178),
.B2(n_152),
.Y(n_202)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_157),
.Y(n_163)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_160),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_168),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_155),
.A2(n_127),
.B1(n_129),
.B2(n_133),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_159),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_144),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_156),
.A2(n_113),
.B1(n_126),
.B2(n_132),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_171),
.A2(n_173),
.B1(n_176),
.B2(n_177),
.Y(n_206)
);

AO21x1_ASAP7_75t_L g198 ( 
.A1(n_172),
.A2(n_180),
.B(n_158),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_153),
.A2(n_120),
.B1(n_135),
.B2(n_123),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_153),
.A2(n_125),
.B1(n_131),
.B2(n_117),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_149),
.A2(n_89),
.B1(n_28),
.B2(n_21),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_152),
.A2(n_143),
.B1(n_140),
.B2(n_151),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_140),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_185),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_145),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_136),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_188),
.C(n_175),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_150),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_195),
.Y(n_208)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_184),
.Y(n_191)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_162),
.B(n_138),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_197),
.Y(n_221)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_184),
.Y(n_193)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_201),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_142),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_139),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_198),
.A2(n_204),
.B1(n_172),
.B2(n_183),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_203),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_137),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_202),
.A2(n_190),
.B1(n_205),
.B2(n_206),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_162),
.B(n_154),
.Y(n_203)
);

BUFx4f_ASAP7_75t_SL g204 ( 
.A(n_182),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_178),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_205),
.A2(n_171),
.B1(n_180),
.B2(n_174),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_164),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_177),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_209),
.A2(n_206),
.B1(n_198),
.B2(n_199),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_188),
.B(n_169),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_218),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_217),
.C(n_224),
.Y(n_232)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_215),
.A2(n_220),
.B(n_196),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_216),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_164),
.C(n_183),
.Y(n_217)
);

OAI322xp33_ASAP7_75t_L g218 ( 
.A1(n_195),
.A2(n_174),
.A3(n_89),
.B1(n_19),
.B2(n_28),
.C1(n_21),
.C2(n_10),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_202),
.A2(n_0),
.B(n_2),
.Y(n_220)
);

A2O1A1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_200),
.A2(n_13),
.B(n_11),
.C(n_9),
.Y(n_223)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_223),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_201),
.B(n_13),
.Y(n_224)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_229),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_231),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_187),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_233),
.Y(n_246)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_237),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_194),
.C(n_204),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_239),
.C(n_211),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_208),
.A2(n_204),
.B1(n_21),
.B2(n_3),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_236),
.B(n_238),
.Y(n_250)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_225),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_42),
.C(n_29),
.Y(n_239)
);

BUFx24_ASAP7_75t_SL g241 ( 
.A(n_240),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_252),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_249),
.C(n_251),
.Y(n_263)
);

A2O1A1O1Ixp25_ASAP7_75t_L g243 ( 
.A1(n_240),
.A2(n_222),
.B(n_219),
.C(n_224),
.D(n_223),
.Y(n_243)
);

OAI21x1_ASAP7_75t_L g255 ( 
.A1(n_243),
.A2(n_226),
.B(n_231),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_219),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_215),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_210),
.C(n_225),
.Y(n_252)
);

AOI21xp33_ASAP7_75t_L g253 ( 
.A1(n_244),
.A2(n_228),
.B(n_227),
.Y(n_253)
);

NOR2xp67_ASAP7_75t_SL g271 ( 
.A(n_253),
.B(n_255),
.Y(n_271)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_247),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_258),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_249),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_261),
.C(n_29),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_246),
.B(n_230),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_236),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_260),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_230),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_248),
.A2(n_234),
.B(n_220),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_214),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_239),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_269),
.Y(n_276)
);

AOI322xp5_ASAP7_75t_L g267 ( 
.A1(n_261),
.A2(n_243),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_0),
.Y(n_267)
);

OAI21x1_ASAP7_75t_L g273 ( 
.A1(n_267),
.A2(n_4),
.B(n_5),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_7),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_256),
.Y(n_269)
);

AOI31xp67_ASAP7_75t_L g270 ( 
.A1(n_263),
.A2(n_0),
.A3(n_2),
.B(n_4),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_272),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_29),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_273),
.A2(n_275),
.B(n_277),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_271),
.A2(n_5),
.B(n_6),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_274),
.A2(n_8),
.B(n_279),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_264),
.A2(n_6),
.B(n_7),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_29),
.C(n_7),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_278),
.B(n_267),
.C(n_8),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_282),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_276),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_283),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_8),
.Y(n_284)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_286),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_287),
.A2(n_285),
.B(n_281),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_284),
.Y(n_289)
);


endmodule