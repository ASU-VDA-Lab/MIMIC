module fake_jpeg_16145_n_148 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_148);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx8_ASAP7_75t_SL g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_20),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_33),
.Y(n_52)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

OAI21xp33_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_28),
.B(n_23),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_14),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_35),
.A2(n_16),
.B1(n_28),
.B2(n_27),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_16),
.B1(n_38),
.B2(n_31),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_27),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_44),
.Y(n_75)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_21),
.B(n_17),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_14),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_47),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_31),
.B(n_21),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_51),
.B(n_17),
.Y(n_64)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_20),
.Y(n_56)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_49),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_61),
.Y(n_80)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_38),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_62),
.A2(n_42),
.B1(n_36),
.B2(n_32),
.Y(n_91)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_67),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_64),
.B(n_68),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_39),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_39),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_47),
.B(n_25),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_71),
.A2(n_9),
.B1(n_6),
.B2(n_7),
.Y(n_92)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_0),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_36),
.Y(n_73)
);

AND2x6_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_28),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_74),
.A2(n_24),
.B(n_48),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_81),
.A2(n_72),
.B1(n_76),
.B2(n_75),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_76),
.A2(n_37),
.B(n_42),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_73),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_50),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_89),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_50),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_91),
.A2(n_66),
.B1(n_67),
.B2(n_69),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_9),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_50),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_89),
.Y(n_104)
);

INVxp33_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_100),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_98),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_82),
.B(n_84),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_90),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_88),
.B1(n_85),
.B2(n_93),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_99),
.A2(n_105),
.B1(n_63),
.B2(n_61),
.Y(n_118)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_70),
.Y(n_103)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_106),
.Y(n_116)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_68),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_83),
.Y(n_112)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_105),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_78),
.C(n_75),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_96),
.C(n_99),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_86),
.B(n_58),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_115),
.A2(n_117),
.B(n_98),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_86),
.B(n_75),
.Y(n_117)
);

NAND2xp33_ASAP7_75t_SL g126 ( 
.A(n_118),
.B(n_74),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_113),
.A2(n_106),
.B1(n_102),
.B2(n_104),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_119),
.A2(n_122),
.B1(n_126),
.B2(n_111),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_121),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_102),
.C(n_101),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_124),
.A2(n_115),
.B(n_117),
.Y(n_127)
);

AO221x1_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_77),
.B1(n_83),
.B2(n_65),
.C(n_59),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_125),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_129),
.C(n_121),
.Y(n_133)
);

BUFx24_ASAP7_75t_SL g129 ( 
.A(n_123),
.Y(n_129)
);

NOR3xp33_ASAP7_75t_SL g130 ( 
.A(n_120),
.B(n_109),
.C(n_110),
.Y(n_130)
);

OA21x2_ASAP7_75t_SL g135 ( 
.A1(n_130),
.A2(n_81),
.B(n_119),
.Y(n_135)
);

AO21x1_ASAP7_75t_SL g137 ( 
.A1(n_132),
.A2(n_81),
.B(n_37),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_134),
.Y(n_138)
);

OAI21x1_ASAP7_75t_L g134 ( 
.A1(n_131),
.A2(n_124),
.B(n_122),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_135),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_116),
.C(n_29),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_131),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_137),
.A2(n_77),
.B1(n_29),
.B2(n_32),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_139),
.A2(n_1),
.B(n_8),
.Y(n_144)
);

AOI322xp5_ASAP7_75t_L g142 ( 
.A1(n_140),
.A2(n_29),
.A3(n_15),
.B1(n_5),
.B2(n_1),
.C1(n_3),
.C2(n_13),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_142),
.Y(n_145)
);

AOI322xp5_ASAP7_75t_L g143 ( 
.A1(n_139),
.A2(n_6),
.A3(n_8),
.B1(n_15),
.B2(n_1),
.C1(n_3),
.C2(n_5),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_143),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_138),
.Y(n_147)
);

OAI32xp33_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_141),
.A3(n_145),
.B1(n_144),
.B2(n_140),
.Y(n_148)
);


endmodule