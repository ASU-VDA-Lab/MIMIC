module fake_jpeg_5364_n_229 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_2),
.B(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_35),
.Y(n_55)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_36),
.B(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_28),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_21),
.Y(n_51)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx4f_ASAP7_75t_SL g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_41),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_39),
.B(n_21),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_40),
.C(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_51),
.Y(n_57)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_49),
.Y(n_83)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_49),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_29),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_36),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_59),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_60),
.B(n_63),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_61),
.A2(n_71),
.B(n_51),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_56),
.B1(n_38),
.B2(n_52),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_62),
.A2(n_45),
.B1(n_29),
.B2(n_24),
.Y(n_93)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_64),
.B(n_65),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_20),
.B1(n_18),
.B2(n_33),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_68),
.Y(n_102)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_47),
.B(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_54),
.B(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_69),
.B(n_75),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_34),
.B(n_18),
.Y(n_71)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_76),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_36),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_82),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_46),
.B(n_17),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_50),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_52),
.A2(n_38),
.B1(n_18),
.B2(n_20),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_78),
.A2(n_80),
.B1(n_84),
.B2(n_25),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_42),
.A2(n_33),
.B1(n_35),
.B2(n_30),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_48),
.B(n_22),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_52),
.A2(n_33),
.B1(n_35),
.B2(n_30),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_35),
.B1(n_40),
.B2(n_37),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_85),
.A2(n_95),
.B1(n_96),
.B2(n_99),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_51),
.B(n_37),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_87),
.B(n_89),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_37),
.B(n_31),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_93),
.B(n_98),
.Y(n_120)
);

OR2x2_ASAP7_75t_SL g94 ( 
.A(n_59),
.B(n_1),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_94),
.A2(n_26),
.B(n_83),
.C(n_3),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_62),
.A2(n_32),
.B1(n_23),
.B2(n_31),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_61),
.A2(n_32),
.B1(n_23),
.B2(n_22),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_50),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_74),
.A2(n_57),
.B1(n_71),
.B2(n_67),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_57),
.B(n_21),
.Y(n_101)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

NOR3xp33_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_24),
.C(n_25),
.Y(n_127)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_107),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_58),
.B(n_21),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_83),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_111),
.A2(n_116),
.B(n_118),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_75),
.B(n_82),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_89),
.B(n_90),
.Y(n_142)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_117),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_81),
.B(n_70),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_58),
.B(n_72),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_99),
.A2(n_64),
.B1(n_72),
.B2(n_70),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_129),
.B1(n_131),
.B2(n_93),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_73),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_121),
.B(n_133),
.Y(n_135)
);

AND2x6_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_88),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_124),
.Y(n_144)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_128),
.Y(n_138)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_86),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_91),
.B(n_98),
.Y(n_125)
);

AOI221xp5_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_127),
.B1(n_132),
.B2(n_95),
.C(n_96),
.Y(n_147)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_85),
.A2(n_73),
.B1(n_76),
.B2(n_83),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_130),
.B(n_15),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_108),
.A2(n_27),
.B1(n_19),
.B2(n_26),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_91),
.A2(n_19),
.B(n_27),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_19),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_113),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_136),
.B(n_140),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_106),
.Y(n_137)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_106),
.Y(n_139)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_105),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_141),
.A2(n_153),
.B1(n_137),
.B2(n_152),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_142),
.B(n_145),
.Y(n_166)
);

OA21x2_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_103),
.B(n_107),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_143),
.A2(n_148),
.B(n_154),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_105),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_146),
.A2(n_149),
.B1(n_111),
.B2(n_5),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_147),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_94),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_19),
.C(n_27),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_120),
.C(n_110),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_1),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_152),
.B(n_130),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_114),
.A2(n_1),
.B(n_2),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_132),
.B(n_4),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_155),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_27),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_156),
.A2(n_136),
.B1(n_150),
.B2(n_148),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_174),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_120),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_162),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_138),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_161),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_126),
.C(n_131),
.Y(n_162)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_111),
.C(n_5),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_154),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_169),
.A2(n_175),
.B(n_168),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_134),
.Y(n_170)
);

BUFx24_ASAP7_75t_SL g180 ( 
.A(n_170),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_171),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_149),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_172)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_172),
.Y(n_183)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_143),
.Y(n_174)
);

OA21x2_ASAP7_75t_SL g177 ( 
.A1(n_160),
.A2(n_148),
.B(n_142),
.Y(n_177)
);

NAND3xp33_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_157),
.C(n_151),
.Y(n_196)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_187),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_185),
.A2(n_151),
.B(n_146),
.Y(n_197)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_156),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_162),
.C(n_167),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_158),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_189),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_178),
.C(n_184),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_188),
.A2(n_165),
.B1(n_159),
.B2(n_156),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_192),
.A2(n_181),
.B1(n_141),
.B2(n_166),
.Y(n_204)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_180),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_193),
.B(n_198),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_181),
.A2(n_165),
.B(n_176),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_195),
.A2(n_197),
.B(n_200),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_196),
.A2(n_179),
.B1(n_157),
.B2(n_164),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_186),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_159),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_199),
.B(n_183),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_207),
.C(n_12),
.Y(n_216)
);

XNOR2x1_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_184),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_203),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_215)
);

AOI322xp5_ASAP7_75t_L g210 ( 
.A1(n_204),
.A2(n_195),
.A3(n_143),
.B1(n_185),
.B2(n_192),
.C1(n_153),
.C2(n_191),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_206),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_135),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_13),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_210),
.A2(n_206),
.B(n_202),
.Y(n_217)
);

INVx11_ASAP7_75t_L g211 ( 
.A(n_208),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_9),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_190),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_213),
.A2(n_8),
.B(n_9),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_215),
.C(n_216),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_217),
.Y(n_225)
);

NAND2xp33_ASAP7_75t_SL g218 ( 
.A(n_211),
.B(n_13),
.Y(n_218)
);

OAI31xp33_ASAP7_75t_SL g223 ( 
.A1(n_218),
.A2(n_219),
.A3(n_10),
.B(n_11),
.Y(n_223)
);

INVxp33_ASAP7_75t_L g224 ( 
.A(n_221),
.Y(n_224)
);

NOR2x1_ASAP7_75t_L g222 ( 
.A(n_220),
.B(n_212),
.Y(n_222)
);

AOI21xp33_ASAP7_75t_L g227 ( 
.A1(n_222),
.A2(n_213),
.B(n_216),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_223),
.B(n_215),
.Y(n_226)
);

OAI221xp5_ASAP7_75t_L g228 ( 
.A1(n_226),
.A2(n_227),
.B1(n_225),
.B2(n_224),
.C(n_11),
.Y(n_228)
);

XOR2x2_ASAP7_75t_SL g229 ( 
.A(n_228),
.B(n_10),
.Y(n_229)
);


endmodule