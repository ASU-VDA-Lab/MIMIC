module fake_jpeg_5698_n_181 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_181);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_181;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_33),
.Y(n_39)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_32),
.A2(n_20),
.B1(n_16),
.B2(n_13),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_36),
.A2(n_37),
.B1(n_47),
.B2(n_48),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_32),
.A2(n_13),
.B1(n_15),
.B2(n_17),
.Y(n_37)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_28),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_17),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_39),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_32),
.A2(n_14),
.B1(n_15),
.B2(n_20),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_31),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_29),
.A2(n_19),
.B1(n_24),
.B2(n_22),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_49),
.A2(n_20),
.B(n_16),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_51),
.B(n_61),
.Y(n_74)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_53),
.Y(n_71)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_27),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_65),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_48),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_58),
.Y(n_75)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_31),
.Y(n_65)
);

FAx1_ASAP7_75t_SL g66 ( 
.A(n_47),
.B(n_33),
.CI(n_28),
.CON(n_66),
.SN(n_66)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_66),
.B(n_16),
.Y(n_80)
);

AOI32xp33_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_46),
.A3(n_28),
.B1(n_38),
.B2(n_26),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_68),
.A2(n_81),
.B(n_23),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_56),
.A2(n_35),
.B1(n_29),
.B2(n_50),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_76),
.B1(n_59),
.B2(n_65),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_50),
.B1(n_42),
.B2(n_26),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_82),
.Y(n_84)
);

AOI32xp33_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_35),
.A3(n_30),
.B1(n_34),
.B2(n_14),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_88),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_82),
.C(n_76),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_94),
.Y(n_114)
);

AO21x1_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_57),
.B(n_65),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_86),
.A2(n_95),
.B(n_96),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_87),
.A2(n_70),
.B1(n_64),
.B2(n_67),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_73),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_53),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_74),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_91),
.Y(n_110)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_93),
.Y(n_106)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_54),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_51),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_72),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_97),
.A2(n_98),
.B(n_67),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_72),
.A2(n_22),
.B(n_24),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_102),
.B(n_105),
.Y(n_119)
);

AOI22x1_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_35),
.B1(n_34),
.B2(n_30),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_111),
.B1(n_78),
.B2(n_41),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_113),
.Y(n_115)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_109),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_70),
.B1(n_78),
.B2(n_34),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_110),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_116),
.B(n_123),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_101),
.B1(n_108),
.B2(n_24),
.Y(n_135)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_107),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_94),
.C(n_93),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_127),
.C(n_128),
.Y(n_138)
);

AOI322xp5_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_95),
.A3(n_96),
.B1(n_84),
.B2(n_91),
.C1(n_85),
.C2(n_86),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_125),
.Y(n_134)
);

OAI21x1_ASAP7_75t_SL g122 ( 
.A1(n_103),
.A2(n_95),
.B(n_86),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_122),
.A2(n_103),
.B1(n_104),
.B2(n_100),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_99),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_105),
.Y(n_124)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_25),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_45),
.C(n_41),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_25),
.Y(n_128)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_136),
.B1(n_126),
.B2(n_118),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_129),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_132),
.A2(n_133),
.B(n_137),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_124),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_139),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_115),
.A2(n_22),
.B1(n_23),
.B2(n_45),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_1),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_140),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_120),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_144),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_119),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_145),
.A2(n_142),
.B1(n_149),
.B2(n_148),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_127),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_150),
.C(n_2),
.Y(n_158)
);

MAJx2_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_128),
.C(n_11),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_149),
.A2(n_10),
.B1(n_3),
.B2(n_4),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_140),
.C(n_139),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_141),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_156),
.C(n_158),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_135),
.Y(n_153)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_153),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_147),
.A2(n_45),
.B1(n_41),
.B2(n_4),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_155),
.Y(n_165)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_150),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_2),
.C(n_3),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_156),
.C(n_158),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_2),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_166),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_6),
.C(n_8),
.Y(n_170)
);

AOI31xp67_ASAP7_75t_SL g164 ( 
.A1(n_159),
.A2(n_3),
.A3(n_5),
.B(n_6),
.Y(n_164)
);

AO21x1_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_6),
.B(n_8),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_5),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_165),
.A2(n_157),
.B(n_7),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_168),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_170),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_8),
.C(n_9),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_9),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_167),
.B1(n_166),
.B2(n_10),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_173),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_176),
.B(n_173),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_178),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_R g180 ( 
.A1(n_179),
.A2(n_177),
.B(n_174),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_175),
.Y(n_181)
);


endmodule