module fake_jpeg_27539_n_167 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_167);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx4f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_26),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_31),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

INVx8_ASAP7_75t_SL g66 ( 
.A(n_15),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_73),
.Y(n_85)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_0),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_65),
.Y(n_75)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_84),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_75),
.B(n_44),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_70),
.A2(n_55),
.B1(n_49),
.B2(n_60),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_79),
.B1(n_80),
.B2(n_45),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_72),
.A2(n_55),
.B1(n_50),
.B2(n_54),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_68),
.A2(n_54),
.B1(n_57),
.B2(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_64),
.B(n_63),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_53),
.B(n_62),
.Y(n_98)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_89),
.B(n_98),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_103),
.B1(n_104),
.B2(n_106),
.Y(n_113)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_85),
.B(n_58),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_101),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_20),
.B(n_43),
.Y(n_101)
);

INVx6_ASAP7_75t_SL g102 ( 
.A(n_81),
.Y(n_102)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_76),
.A2(n_52),
.B1(n_48),
.B2(n_46),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_80),
.A2(n_52),
.B1(n_59),
.B2(n_56),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_105),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_85),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_47),
.B1(n_62),
.B2(n_17),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_107),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_105),
.A2(n_12),
.B1(n_41),
.B2(n_36),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_108),
.A2(n_93),
.B1(n_4),
.B2(n_5),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_107),
.B1(n_92),
.B2(n_5),
.Y(n_128)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_120),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_122),
.Y(n_131)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_127),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_100),
.C(n_91),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_97),
.C(n_109),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_90),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_114),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_94),
.Y(n_126)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_113),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_128),
.A2(n_129),
.B1(n_3),
.B2(n_6),
.Y(n_139)
);

INVxp67_ASAP7_75t_SL g130 ( 
.A(n_123),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_135),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_133),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_120),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_128),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_126),
.Y(n_136)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_125),
.A2(n_117),
.B(n_111),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_140),
.C(n_142),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_139),
.A2(n_134),
.B1(n_141),
.B2(n_142),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_109),
.C(n_18),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_145),
.Y(n_154)
);

OA21x2_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_13),
.B(n_35),
.Y(n_147)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_131),
.B1(n_7),
.B2(n_8),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_150),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_135),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_150)
);

FAx1_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_144),
.CI(n_148),
.CON(n_155),
.SN(n_155)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_155),
.B(n_156),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_151),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_146),
.B1(n_143),
.B2(n_152),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_146),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_153),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_147),
.C(n_22),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_19),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_163),
.A2(n_24),
.B(n_34),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_10),
.B(n_33),
.Y(n_165)
);

CKINVDCx12_ASAP7_75t_R g166 ( 
.A(n_165),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_9),
.Y(n_167)
);


endmodule