module fake_ariane_1880_n_116 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_30, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_116);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_30;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_116;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_106;
wire n_53;
wire n_111;
wire n_115;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_49;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_107;
wire n_72;
wire n_105;
wire n_44;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_112;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_61;
wire n_108;
wire n_102;
wire n_43;
wire n_81;
wire n_87;
wire n_41;
wire n_55;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_35;
wire n_54;

BUFx3_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_10),
.B(n_3),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

OAI21x1_ASAP7_75t_L g38 ( 
.A1(n_6),
.A2(n_21),
.B(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

AND2x4_ASAP7_75t_L g41 ( 
.A(n_7),
.B(n_5),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_4),
.B(n_13),
.Y(n_42)
);

NOR2x1_ASAP7_75t_L g43 ( 
.A(n_8),
.B(n_14),
.Y(n_43)
);

AND2x4_ASAP7_75t_L g44 ( 
.A(n_2),
.B(n_24),
.Y(n_44)
);

BUFx8_ASAP7_75t_SL g45 ( 
.A(n_1),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_11),
.A2(n_0),
.B1(n_23),
.B2(n_26),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

NAND3xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_46),
.C(n_35),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_SL g56 ( 
.A(n_50),
.B(n_16),
.C(n_27),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_30),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_33),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_53),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_31),
.B(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_31),
.B(n_53),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_51),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

AO221x1_ASAP7_75t_L g67 ( 
.A1(n_37),
.A2(n_52),
.B1(n_47),
.B2(n_39),
.C(n_45),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_52),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_57),
.B(n_58),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_52),
.Y(n_73)
);

NOR3xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_34),
.C(n_42),
.Y(n_74)
);

AND2x4_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_41),
.Y(n_75)
);

OAI21x1_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_38),
.B(n_43),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_48),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_41),
.Y(n_79)
);

OAI22x1_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_44),
.B1(n_34),
.B2(n_32),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

OAI21x1_ASAP7_75t_L g83 ( 
.A1(n_76),
.A2(n_59),
.B(n_61),
.Y(n_83)
);

AO21x1_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_44),
.B(n_61),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_80),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

NAND2x1p5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_39),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

AND2x4_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_59),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_69),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_80),
.B1(n_75),
.B2(n_79),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_75),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_86),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_86),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_93),
.B(n_84),
.Y(n_101)
);

NOR3xp33_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_85),
.C(n_87),
.Y(n_102)
);

XOR2x2_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_92),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g104 ( 
.A1(n_99),
.A2(n_92),
.B1(n_100),
.B2(n_85),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_96),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_102),
.A2(n_95),
.B1(n_100),
.B2(n_82),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_103),
.A2(n_83),
.B(n_88),
.Y(n_107)
);

NAND5xp2_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_78),
.C(n_96),
.D(n_84),
.E(n_88),
.Y(n_108)
);

NAND5xp2_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_88),
.C(n_37),
.D(n_47),
.E(n_52),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_106),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_47),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_111),
.Y(n_112)
);

AND4x1_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_97),
.C(n_98),
.D(n_39),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_112),
.A2(n_113),
.B1(n_70),
.B2(n_83),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_70),
.Y(n_115)
);

OR2x6_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_70),
.Y(n_116)
);


endmodule