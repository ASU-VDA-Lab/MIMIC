module fake_jpeg_6392_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_10),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_42),
.B(n_44),
.Y(n_87)
);

INVx2_ASAP7_75t_R g43 ( 
.A(n_32),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_46),
.Y(n_66)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_47),
.B1(n_17),
.B2(n_38),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_0),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_32),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_48),
.B(n_26),
.Y(n_109)
);

BUFx24_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_20),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_59),
.Y(n_72)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_52),
.B(n_54),
.Y(n_112)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_23),
.B(n_10),
.Y(n_56)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_57),
.B(n_65),
.Y(n_111)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_23),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_24),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_64),
.Y(n_73)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_24),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx11_ASAP7_75t_L g149 ( 
.A(n_67),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_17),
.B1(n_38),
.B2(n_16),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_68),
.A2(n_70),
.B1(n_74),
.B2(n_77),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_69),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_38),
.B1(n_16),
.B2(n_40),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_71),
.B(n_75),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_53),
.A2(n_40),
.B1(n_25),
.B2(n_30),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_30),
.B1(n_25),
.B2(n_33),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_45),
.A2(n_31),
.B1(n_28),
.B2(n_33),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_78),
.A2(n_82),
.B1(n_90),
.B2(n_98),
.Y(n_122)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_79),
.B(n_80),
.Y(n_131)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_64),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_81),
.B(n_92),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_47),
.A2(n_31),
.B1(n_28),
.B2(n_35),
.Y(n_82)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_84),
.B(n_86),
.Y(n_135)
);

BUFx16f_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_88),
.B(n_91),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_59),
.A2(n_18),
.B1(n_22),
.B2(n_27),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_95),
.B1(n_96),
.B2(n_101),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_61),
.A2(n_18),
.B1(n_22),
.B2(n_27),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_48),
.B(n_32),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_54),
.A2(n_39),
.B1(n_21),
.B2(n_29),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_58),
.A2(n_39),
.B1(n_21),
.B2(n_29),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_97),
.B(n_102),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_49),
.A2(n_29),
.B1(n_37),
.B2(n_41),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_49),
.A2(n_39),
.B1(n_21),
.B2(n_37),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_46),
.B(n_12),
.Y(n_102)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_43),
.A2(n_29),
.B1(n_37),
.B2(n_41),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_107),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_129)
);

AO21x1_ASAP7_75t_L g133 ( 
.A1(n_109),
.A2(n_9),
.B(n_14),
.Y(n_133)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_114),
.B(n_123),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_66),
.B(n_41),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_115),
.B(n_120),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_66),
.B(n_41),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_121),
.Y(n_177)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_72),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_127),
.Y(n_161)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_100),
.A2(n_36),
.B1(n_26),
.B2(n_10),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_128),
.A2(n_123),
.B1(n_125),
.B2(n_144),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_129),
.A2(n_99),
.B1(n_143),
.B2(n_127),
.Y(n_181)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_137),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_73),
.B(n_0),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_140),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_133),
.A2(n_76),
.B1(n_108),
.B2(n_109),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_100),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_134),
.A2(n_116),
.B1(n_145),
.B2(n_146),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_136),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_111),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_112),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_138),
.B(n_142),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_82),
.B(n_78),
.Y(n_140)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_145),
.Y(n_153)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_77),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_74),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_146),
.B(n_148),
.Y(n_154)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_70),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_104),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_87),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_152),
.B(n_155),
.Y(n_200)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_150),
.B(n_108),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_167),
.Y(n_196)
);

INVxp33_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_164),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_136),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_159),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_107),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_168),
.C(n_170),
.Y(n_190)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_165),
.B(n_166),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_121),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_139),
.B(n_126),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_69),
.Y(n_168)
);

XNOR2x1_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_98),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_101),
.C(n_110),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_119),
.C(n_136),
.Y(n_209)
);

O2A1O1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_118),
.A2(n_110),
.B(n_86),
.C(n_99),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_172),
.A2(n_183),
.B(n_15),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_173),
.A2(n_121),
.B(n_15),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_132),
.B(n_104),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_174),
.B(n_176),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_175),
.A2(n_185),
.B1(n_119),
.B2(n_142),
.Y(n_210)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_178),
.B(n_113),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_3),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_180),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_122),
.B(n_7),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_116),
.B(n_7),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_184),
.Y(n_207)
);

O2A1O1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_133),
.A2(n_103),
.B(n_11),
.C(n_13),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_113),
.B(n_9),
.Y(n_184)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_136),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_187),
.Y(n_218)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_189),
.Y(n_222)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_170),
.A2(n_125),
.B1(n_149),
.B2(n_103),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_191),
.A2(n_192),
.B1(n_216),
.B2(n_220),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_178),
.A2(n_182),
.B1(n_180),
.B2(n_163),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_193),
.B(n_194),
.Y(n_231)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_195),
.Y(n_223)
);

FAx1_ASAP7_75t_SL g197 ( 
.A(n_160),
.B(n_130),
.CI(n_149),
.CON(n_197),
.SN(n_197)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_211),
.Y(n_224)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_202),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g203 ( 
.A(n_164),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_203),
.Y(n_226)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_204),
.Y(n_230)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_215),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_210),
.A2(n_177),
.B1(n_211),
.B2(n_209),
.Y(n_242)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_173),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_153),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_163),
.B(n_121),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_214),
.Y(n_227)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_154),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_168),
.B(n_162),
.C(n_167),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_175),
.A2(n_114),
.B1(n_11),
.B2(n_14),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_154),
.B(n_9),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_176),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_221),
.A2(n_184),
.B(n_157),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_192),
.A2(n_172),
.B1(n_171),
.B2(n_153),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_233),
.A2(n_236),
.B1(n_237),
.B2(n_245),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_238),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_205),
.A2(n_152),
.B1(n_162),
.B2(n_165),
.Y(n_236)
);

AOI22x1_ASAP7_75t_SL g237 ( 
.A1(n_190),
.A2(n_185),
.B1(n_183),
.B2(n_179),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_194),
.B(n_151),
.Y(n_239)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_239),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_190),
.A2(n_151),
.B(n_159),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_166),
.Y(n_241)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_241),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_221),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_196),
.A2(n_177),
.B(n_215),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_244),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_196),
.A2(n_177),
.B(n_207),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_191),
.A2(n_216),
.B1(n_200),
.B2(n_210),
.Y(n_245)
);

NAND3xp33_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_197),
.C(n_207),
.Y(n_246)
);

BUFx12f_ASAP7_75t_SL g249 ( 
.A(n_246),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_197),
.B(n_198),
.Y(n_247)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_247),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_198),
.B(n_199),
.Y(n_248)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_248),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_208),
.C(n_218),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_250),
.B(n_253),
.C(n_256),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_251),
.A2(n_237),
.B(n_248),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_188),
.C(n_217),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_228),
.B(n_222),
.Y(n_255)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_255),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_201),
.C(n_205),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_195),
.Y(n_258)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_258),
.Y(n_287)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_220),
.C(n_212),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_261),
.B(n_246),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_222),
.B(n_189),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_262),
.B(n_265),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_203),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_263),
.A2(n_234),
.B(n_231),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_229),
.B(n_203),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_227),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_266),
.B(n_229),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_203),
.C(n_224),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_268),
.C(n_237),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_227),
.C(n_241),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_285),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_239),
.Y(n_272)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_275),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_269),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_279),
.C(n_280),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_242),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_249),
.A2(n_232),
.B1(n_245),
.B2(n_233),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_276),
.A2(n_283),
.B1(n_260),
.B2(n_257),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_249),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_286),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_252),
.Y(n_281)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_281),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_270),
.A2(n_232),
.B1(n_236),
.B2(n_231),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_253),
.B(n_225),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_279),
.C(n_250),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_293),
.C(n_274),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_256),
.C(n_268),
.Y(n_293)
);

A2O1A1O1Ixp25_ASAP7_75t_L g295 ( 
.A1(n_271),
.A2(n_257),
.B(n_261),
.C(n_267),
.D(n_263),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_275),
.Y(n_305)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_287),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_296),
.B(n_297),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_282),
.Y(n_297)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_283),
.A2(n_254),
.B1(n_236),
.B2(n_226),
.Y(n_300)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_300),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_276),
.A2(n_230),
.B1(n_223),
.B2(n_225),
.Y(n_301)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_301),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_296),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_310),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_290),
.B(n_287),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_306),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_307),
.C(n_311),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_299),
.B(n_284),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_289),
.A2(n_277),
.B1(n_273),
.B2(n_280),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_281),
.Y(n_311)
);

NOR2xp67_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_295),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_314),
.A2(n_291),
.B(n_298),
.Y(n_322)
);

NAND2xp67_ASAP7_75t_SL g315 ( 
.A(n_310),
.B(n_300),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_312),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_301),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_316),
.A2(n_294),
.B1(n_238),
.B2(n_223),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_292),
.C(n_293),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_291),
.C(n_305),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_302),
.B(n_272),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_320),
.A2(n_321),
.B(n_288),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_230),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_323),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_324),
.A2(n_325),
.B(n_317),
.Y(n_331)
);

NOR2xp67_ASAP7_75t_SL g330 ( 
.A(n_326),
.B(n_327),
.Y(n_330)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_313),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_319),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_329),
.B(n_331),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_330),
.B(n_318),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_328),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_332),
.Y(n_337)
);


endmodule