module real_jpeg_326_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_1),
.A2(n_59),
.B1(n_60),
.B2(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_1),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_1),
.A2(n_35),
.B1(n_37),
.B2(n_114),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_114),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_1),
.A2(n_46),
.B1(n_50),
.B2(n_114),
.Y(n_228)
);

BUFx4f_ASAP7_75t_L g104 ( 
.A(n_2),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_3),
.A2(n_59),
.B1(n_60),
.B2(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_3),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_3),
.A2(n_35),
.B1(n_37),
.B2(n_153),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_153),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_3),
.A2(n_46),
.B1(n_50),
.B2(n_153),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_4),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_4),
.A2(n_39),
.B1(n_59),
.B2(n_60),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_39),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_4),
.A2(n_39),
.B1(n_46),
.B2(n_50),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_5),
.B(n_59),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_5),
.B(n_85),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_5),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_5),
.A2(n_59),
.B(n_188),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_5),
.B(n_27),
.Y(n_250)
);

AOI21xp33_ASAP7_75t_L g257 ( 
.A1(n_5),
.A2(n_37),
.B(n_258),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_5),
.B(n_46),
.C(n_49),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_224),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_5),
.B(n_103),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_5),
.B(n_44),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_6),
.A2(n_35),
.B1(n_37),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_42),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_6),
.A2(n_42),
.B1(n_46),
.B2(n_50),
.Y(n_106)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_11),
.A2(n_59),
.B1(n_60),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_11),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_11),
.A2(n_35),
.B1(n_37),
.B2(n_69),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_69),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_11),
.A2(n_46),
.B1(n_50),
.B2(n_69),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_12),
.A2(n_59),
.B1(n_60),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_12),
.A2(n_35),
.B1(n_37),
.B2(n_72),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_72),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_L g215 ( 
.A1(n_12),
.A2(n_46),
.B1(n_50),
.B2(n_72),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_13),
.A2(n_59),
.B1(n_60),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_13),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_13),
.A2(n_35),
.B1(n_37),
.B2(n_198),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_198),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_13),
.A2(n_46),
.B1(n_50),
.B2(n_198),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_14),
.A2(n_59),
.B1(n_60),
.B2(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_14),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_14),
.A2(n_35),
.B1(n_37),
.B2(n_179),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_179),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_14),
.A2(n_46),
.B1(n_50),
.B2(n_179),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_16),
.A2(n_59),
.B1(n_60),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_16),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_16),
.A2(n_35),
.B1(n_37),
.B2(n_67),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_16),
.A2(n_28),
.B1(n_29),
.B2(n_67),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_16),
.A2(n_46),
.B1(n_50),
.B2(n_67),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_91),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_89),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_78),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_21),
.B(n_78),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_70),
.C(n_73),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_22),
.A2(n_70),
.B1(n_122),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_22),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_55),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_43),
.B2(n_54),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_25),
.B(n_43),
.C(n_55),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_25)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_26),
.A2(n_40),
.B1(n_119),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_26),
.A2(n_40),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_26),
.A2(n_40),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_26),
.A2(n_40),
.B1(n_194),
.B2(n_210),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_26),
.A2(n_40),
.B1(n_209),
.B2(n_257),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_34),
.Y(n_26)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_27),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_27),
.A2(n_76),
.B(n_81),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_27),
.A2(n_75),
.B1(n_76),
.B2(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_27),
.A2(n_76),
.B1(n_149),
.B2(n_176),
.Y(n_175)
);

AO22x2_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_28),
.A2(n_29),
.B1(n_48),
.B2(n_49),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_28),
.B(n_33),
.Y(n_225)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI32xp33_ASAP7_75t_L g222 ( 
.A1(n_29),
.A2(n_31),
.A3(n_37),
.B1(n_223),
.B2(n_225),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_29),
.B(n_266),
.Y(n_265)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_33),
.B1(n_35),
.B2(n_37),
.Y(n_34)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_35),
.A2(n_37),
.B1(n_62),
.B2(n_63),
.Y(n_65)
);

NAND2xp33_ASAP7_75t_SL g189 ( 
.A(n_35),
.B(n_62),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_35),
.B(n_224),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI32xp33_ASAP7_75t_L g187 ( 
.A1(n_37),
.A2(n_60),
.A3(n_63),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_38),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_41),
.Y(n_81)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_70),
.C(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_43),
.A2(n_54),
.B1(n_74),
.B2(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_51),
.B(n_53),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_44),
.A2(n_51),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_44),
.A2(n_51),
.B1(n_53),
.B2(n_110),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_44),
.A2(n_51),
.B1(n_109),
.B2(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_44),
.A2(n_51),
.B1(n_218),
.B2(n_220),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_44),
.A2(n_51),
.B1(n_220),
.B2(n_240),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_44),
.A2(n_51),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_44),
.A2(n_51),
.B1(n_248),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_45),
.A2(n_146),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_45),
.A2(n_172),
.B1(n_219),
.B2(n_260),
.Y(n_259)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_45)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_46),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_46),
.B(n_276),
.Y(n_275)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_51),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_56),
.A2(n_65),
.B1(n_66),
.B2(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_56),
.A2(n_65),
.B1(n_71),
.B2(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_56),
.A2(n_65),
.B1(n_113),
.B2(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_56),
.A2(n_65),
.B1(n_197),
.B2(n_199),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_56),
.A2(n_65),
.B1(n_197),
.B2(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_57),
.A2(n_85),
.B1(n_152),
.B2(n_178),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_65),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_68),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_70),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_73),
.B(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_88),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B1(n_86),
.B2(n_87),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_80),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AO21x1_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_159),
.B(n_316),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_154),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_128),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_95),
.B(n_128),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_115),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_96),
.B(n_121),
.C(n_126),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_111),
.B(n_112),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_97),
.A2(n_98),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_107),
.Y(n_98)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_99),
.A2(n_111),
.B1(n_112),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_99),
.A2(n_107),
.B1(n_108),
.B2(n_111),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_102),
.B(n_105),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_100),
.A2(n_102),
.B1(n_142),
.B2(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_100),
.A2(n_102),
.B1(n_227),
.B2(n_229),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_100),
.A2(n_102),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_101),
.A2(n_103),
.B1(n_106),
.B2(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_101),
.A2(n_103),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_101),
.A2(n_103),
.B1(n_191),
.B2(n_215),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_101),
.A2(n_103),
.B1(n_228),
.B2(n_252),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_101),
.A2(n_103),
.B1(n_224),
.B2(n_278),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_101),
.A2(n_103),
.B1(n_278),
.B2(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_121),
.B1(n_126),
.B2(n_127),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_116),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_117),
.B(n_120),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

INVxp33_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_121),
.Y(n_127)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_134),
.C(n_136),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_130),
.B1(n_134),
.B2(n_135),
.Y(n_162)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_147),
.C(n_150),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_137),
.A2(n_138),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_139),
.A2(n_140),
.B1(n_143),
.B2(n_144),
.Y(n_200)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_150),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_154),
.A2(n_317),
.B(n_318),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_158),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_155),
.B(n_158),
.Y(n_318)
);

AO21x1_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_180),
.B(n_315),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_161),
.B(n_163),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.C(n_168),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_167),
.Y(n_202)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_165),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_202),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_175),
.C(n_177),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_170),
.B(n_173),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_171),
.Y(n_240)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_177),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_176),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_203),
.B(n_314),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_201),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_182),
.B(n_201),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.C(n_200),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_183),
.B(n_200),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_185),
.B(n_301),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_193),
.C(n_196),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_186),
.B(n_304),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_187),
.B(n_190),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_193),
.B(n_196),
.Y(n_304)
);

AOI31xp33_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_298),
.A3(n_307),
.B(n_311),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_243),
.B(n_297),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_230),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_206),
.B(n_230),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_217),
.C(n_221),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_207),
.B(n_294),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_212),
.C(n_216),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_216),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_214),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_217),
.B(n_221),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_226),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_226),
.Y(n_254)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_223),
.Y(n_258)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_232),
.B(n_233),
.C(n_234),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_235),
.B(n_238),
.C(n_242),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_241),
.B2(n_242),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_238),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_239),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_292),
.B(n_296),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_261),
.B(n_291),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_253),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_246),
.B(n_253),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_250),
.C(n_251),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_250),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_249),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_271),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_252),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_254),
.B(n_256),
.C(n_259),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_259),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_272),
.B(n_290),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_270),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_270),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_267),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_264),
.A2(n_265),
.B1(n_267),
.B2(n_268),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_284),
.B(n_289),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_279),
.B(n_283),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_281),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_282),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_288),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_288),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_295),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_295),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_299),
.A2(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_302),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_302),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_305),
.C(n_306),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_310),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_306),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_309),
.Y(n_312)
);


endmodule