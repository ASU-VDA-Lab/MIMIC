module fake_jpeg_13593_n_177 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_177);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_33),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_8),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_13),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_31),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_44),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_24),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_4),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_2),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_4),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_2),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_42),
.Y(n_77)
);

BUFx8_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_0),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_83),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_0),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_74),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_77),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

HAxp5_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_1),
.CON(n_86),
.SN(n_86)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_86),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_1),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_56),
.Y(n_103)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_88),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_65),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_55),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_73),
.Y(n_109)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_58),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_53),
.C(n_54),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_5),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_72),
.B1(n_71),
.B2(n_69),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_69),
.B1(n_67),
.B2(n_76),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_103),
.B(n_67),
.Y(n_106)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_111),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_107),
.B(n_115),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_109),
.B(n_117),
.Y(n_128)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_76),
.B1(n_60),
.B2(n_71),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_120),
.B1(n_10),
.B2(n_11),
.Y(n_138)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_116),
.Y(n_142)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_114),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_75),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_101),
.B(n_63),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_98),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_118),
.B(n_122),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_119),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_95),
.A2(n_60),
.B1(n_64),
.B2(n_62),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_59),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_124),
.Y(n_132)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_70),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_10),
.C(n_11),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_3),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_127),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_92),
.C(n_22),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_146),
.C(n_135),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_92),
.B1(n_6),
.B2(n_7),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_131),
.A2(n_134),
.B1(n_147),
.B2(n_114),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_108),
.B(n_25),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_141),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_121),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_143),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_146),
.Y(n_155)
);

AND2x6_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_26),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_107),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_129),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_27),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_105),
.A2(n_12),
.B1(n_14),
.B2(n_16),
.Y(n_147)
);

AO22x1_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_50),
.B1(n_28),
.B2(n_17),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_SL g150 ( 
.A1(n_149),
.A2(n_12),
.B(n_14),
.C(n_18),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_157),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_152),
.A2(n_155),
.B1(n_160),
.B2(n_133),
.Y(n_163)
);

NOR2xp67_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_19),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_154),
.Y(n_167)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_128),
.B(n_140),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_158),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_132),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_139),
.A2(n_20),
.B(n_21),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_130),
.C(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_136),
.C(n_145),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_163),
.A2(n_157),
.B1(n_149),
.B2(n_150),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_168),
.C(n_161),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_166),
.A2(n_162),
.B(n_155),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_170),
.C(n_171),
.Y(n_172)
);

AO22x1_ASAP7_75t_SL g173 ( 
.A1(n_172),
.A2(n_165),
.B1(n_150),
.B2(n_141),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_151),
.B(n_167),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_174),
.A2(n_167),
.B1(n_29),
.B2(n_30),
.Y(n_175)
);

AOI21x1_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_23),
.B(n_35),
.Y(n_176)
);

A2O1A1O1Ixp25_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_41),
.B(n_43),
.C(n_45),
.D(n_48),
.Y(n_177)
);


endmodule