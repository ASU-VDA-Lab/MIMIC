module fake_jpeg_26057_n_287 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_287);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_287;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_13;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVxp67_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_19),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_29),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_19),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_18),
.Y(n_33)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_32),
.A2(n_21),
.B1(n_18),
.B2(n_23),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_21),
.B1(n_18),
.B2(n_23),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_40),
.B(n_33),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_21),
.B1(n_24),
.B2(n_22),
.Y(n_42)
);

O2A1O1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_46),
.B(n_28),
.C(n_29),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_25),
.B1(n_24),
.B2(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_50),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_43),
.B(n_28),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_31),
.C(n_44),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_31),
.C(n_35),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_57),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_62),
.B1(n_36),
.B2(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_60),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_45),
.B(n_31),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_29),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_61),
.A2(n_36),
.B1(n_47),
.B2(n_38),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_36),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_64),
.Y(n_85)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_28),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_77),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_37),
.B1(n_30),
.B2(n_40),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_84),
.B1(n_56),
.B2(n_61),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_76),
.C(n_26),
.Y(n_102)
);

OAI32xp33_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_40),
.A3(n_46),
.B1(n_31),
.B2(n_42),
.Y(n_74)
);

AOI32xp33_ASAP7_75t_L g100 ( 
.A1(n_74),
.A2(n_12),
.A3(n_14),
.B1(n_20),
.B2(n_16),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_55),
.B(n_58),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_34),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_31),
.C(n_26),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_83),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_61),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_49),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_62),
.A2(n_47),
.B1(n_39),
.B2(n_35),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_86),
.A2(n_63),
.B1(n_47),
.B2(n_65),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_70),
.B(n_50),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_88),
.B(n_90),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_89),
.A2(n_91),
.B1(n_100),
.B2(n_30),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_59),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_80),
.B(n_53),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_97),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

NOR2x1_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_62),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_96),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_63),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_99),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_65),
.Y(n_99)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_73),
.C(n_26),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_78),
.A2(n_25),
.B(n_35),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_103),
.A2(n_78),
.B(n_85),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_71),
.A2(n_63),
.B1(n_41),
.B2(n_15),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_104),
.A2(n_69),
.B1(n_72),
.B2(n_68),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_33),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_106),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_54),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_106),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_114),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_94),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_109),
.Y(n_139)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_113),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_95),
.A2(n_84),
.B1(n_74),
.B2(n_76),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_112),
.A2(n_91),
.B1(n_89),
.B2(n_100),
.Y(n_130)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_96),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_117),
.Y(n_144)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_20),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_121),
.B1(n_97),
.B2(n_105),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_127),
.C(n_128),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_91),
.A2(n_95),
.B(n_87),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_73),
.C(n_26),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_54),
.C(n_49),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_91),
.A2(n_86),
.B(n_15),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_129),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_153),
.B1(n_121),
.B2(n_119),
.Y(n_155)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_132),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_107),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_135),
.B(n_137),
.Y(n_171)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_88),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_113),
.B(n_109),
.Y(n_156)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_140),
.A2(n_149),
.B(n_151),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_141),
.A2(n_146),
.B1(n_114),
.B2(n_116),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_145),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_107),
.A2(n_103),
.B1(n_101),
.B2(n_90),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_147),
.B(n_129),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_101),
.Y(n_148)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_72),
.Y(n_152)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_112),
.A2(n_69),
.B1(n_68),
.B2(n_64),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_20),
.Y(n_154)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_155),
.A2(n_130),
.B(n_133),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_156),
.B(n_174),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_162),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_127),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_166),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_139),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_161),
.B(n_133),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_168),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_127),
.C(n_123),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_170),
.C(n_175),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_152),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_173),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_123),
.C(n_111),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_151),
.A2(n_117),
.B1(n_125),
.B2(n_121),
.Y(n_172)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_172),
.Y(n_183)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_118),
.C(n_126),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_134),
.A2(n_110),
.B1(n_69),
.B2(n_64),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_178),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_132),
.A2(n_143),
.B1(n_146),
.B2(n_153),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_170),
.Y(n_203)
);

NOR2x1_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_143),
.Y(n_181)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_186),
.B(n_188),
.Y(n_206)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_177),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_190),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_191),
.A2(n_196),
.B1(n_199),
.B2(n_176),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_194),
.A2(n_198),
.B(n_191),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_159),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_200),
.C(n_185),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_144),
.Y(n_196)
);

BUFx24_ASAP7_75t_SL g212 ( 
.A(n_197),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_144),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_140),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_160),
.B(n_137),
.C(n_135),
.Y(n_200)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_214),
.C(n_216),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_167),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_205),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_179),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_213),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_189),
.A2(n_164),
.B1(n_174),
.B2(n_131),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_208),
.A2(n_211),
.B1(n_193),
.B2(n_194),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_183),
.A2(n_33),
.B1(n_9),
.B2(n_11),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_16),
.C(n_20),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_201),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_30),
.Y(n_216)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_218),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_199),
.B(n_196),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_SL g229 ( 
.A(n_219),
.B(n_220),
.C(n_181),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_198),
.B(n_9),
.Y(n_220)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_231),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_184),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_230),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_187),
.B(n_182),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_228),
.A2(n_236),
.B(n_216),
.Y(n_238)
);

AOI322xp5_ASAP7_75t_L g247 ( 
.A1(n_229),
.A2(n_232),
.A3(n_8),
.B1(n_7),
.B2(n_13),
.C1(n_3),
.C2(n_4),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_215),
.A2(n_187),
.B1(n_184),
.B2(n_30),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_219),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_206),
.A2(n_33),
.B1(n_51),
.B2(n_17),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_210),
.A2(n_51),
.B1(n_41),
.B2(n_17),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_235),
.Y(n_240)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_220),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_214),
.A2(n_8),
.B(n_11),
.Y(n_236)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_203),
.Y(n_241)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_241),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_41),
.C(n_38),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_243),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_41),
.C(n_38),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_225),
.A2(n_7),
.B(n_9),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_245),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_230),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_38),
.C(n_17),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_246),
.B(n_38),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_247),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_260)
);

AO221x1_ASAP7_75t_L g249 ( 
.A1(n_221),
.A2(n_233),
.B1(n_228),
.B2(n_227),
.C(n_222),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_249),
.A2(n_8),
.B(n_1),
.Y(n_251)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_251),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_255),
.B(n_259),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_13),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_237),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_239),
.B(n_13),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_258),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_248),
.A2(n_0),
.B(n_1),
.Y(n_258)
);

AO22x1_ASAP7_75t_L g259 ( 
.A1(n_245),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_240),
.C(n_246),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_264),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_243),
.C(n_27),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_267),
.Y(n_275)
);

XNOR2x1_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_2),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_250),
.B(n_2),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_269),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_254),
.B(n_3),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_261),
.A2(n_256),
.B1(n_259),
.B2(n_6),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_273),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_263),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_261),
.Y(n_278)
);

NOR2x1_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_4),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_272),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_277),
.A2(n_27),
.B(n_5),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_275),
.C(n_274),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_279),
.B(n_280),
.C(n_276),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_281),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_282),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_5),
.C(n_6),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_284),
.B(n_27),
.C(n_279),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_27),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_286),
.A2(n_27),
.B(n_261),
.Y(n_287)
);


endmodule