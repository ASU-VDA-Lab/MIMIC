module fake_jpeg_19658_n_49 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_49);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_49;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_1),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_3),
.B(n_0),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_5),
.B(n_0),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g15 ( 
.A(n_4),
.B(n_0),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_12),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_17),
.A2(n_14),
.B1(n_21),
.B2(n_23),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_19),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_2),
.Y(n_19)
);

A2O1A1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_13),
.A2(n_3),
.B(n_8),
.C(n_15),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_20),
.A2(n_24),
.B(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_12),
.A2(n_16),
.B1(n_15),
.B2(n_7),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_24),
.A2(n_14),
.B1(n_25),
.B2(n_19),
.Y(n_29)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_20),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_29),
.A2(n_30),
.B1(n_37),
.B2(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_33),
.B(n_34),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_19),
.C(n_18),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_33),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_19),
.A2(n_15),
.B1(n_12),
.B2(n_16),
.Y(n_37)
);

OAI32xp33_ASAP7_75t_L g41 ( 
.A1(n_36),
.A2(n_29),
.A3(n_32),
.B1(n_35),
.B2(n_31),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_39),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_27),
.Y(n_43)
);

NAND3xp33_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_31),
.C(n_28),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_38),
.Y(n_47)
);

FAx1_ASAP7_75t_SL g45 ( 
.A(n_41),
.B(n_42),
.CI(n_40),
.CON(n_45),
.SN(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_45),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_46),
.Y(n_49)
);


endmodule