module fake_ibex_1759_n_864 (n_151, n_147, n_85, n_128, n_84, n_64, n_3, n_73, n_152, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_120, n_93, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_132, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_864);

input n_151;
input n_147;
input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_120;
input n_93;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_132;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_864;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_593;
wire n_862;
wire n_545;
wire n_583;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_608;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_375;
wire n_280;
wire n_317;
wire n_340;
wire n_708;
wire n_187;
wire n_667;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_723;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_840;
wire n_561;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_158;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_711;
wire n_228;
wire n_671;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_732;
wire n_798;
wire n_832;
wire n_673;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_155;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_758;
wire n_636;
wire n_594;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_844;
wire n_245;
wire n_648;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_589;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_704;
wire n_643;
wire n_841;
wire n_679;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_718;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_392;
wire n_206;
wire n_354;
wire n_630;
wire n_567;
wire n_548;
wire n_516;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_564;
wire n_562;
wire n_506;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_190;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_247;
wire n_288;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_741;
wire n_807;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_820;
wire n_805;
wire n_670;
wire n_728;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_266;
wire n_294;
wire n_485;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_794;
wire n_260;
wire n_620;
wire n_836;
wire n_683;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_687;
wire n_159;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_559;
wire n_425;

INVxp67_ASAP7_75t_L g155 ( 
.A(n_17),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_130),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_53),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_43),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_4),
.Y(n_160)
);

NOR2xp67_ASAP7_75t_L g161 ( 
.A(n_106),
.B(n_128),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_107),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_75),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_36),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_19),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_37),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_153),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_69),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_103),
.Y(n_169)
);

BUFx10_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_5),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_82),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_131),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_115),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_64),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_120),
.B(n_108),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_29),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_46),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_44),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_133),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_27),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_85),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_122),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_5),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_73),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_12),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_125),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_134),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_137),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_63),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_139),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_78),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_52),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_119),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_104),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_145),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_154),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_124),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_88),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_66),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_140),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_14),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_42),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_91),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_51),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_101),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_60),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_36),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_24),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_94),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_35),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_87),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_34),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_41),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_141),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_152),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_57),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_109),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_99),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_114),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_74),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_29),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_7),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_24),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_97),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_33),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_116),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_3),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_27),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_81),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_58),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_150),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_56),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_100),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_77),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_138),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_102),
.B(n_144),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_80),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_89),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_0),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_7),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_31),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_126),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_121),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_142),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_55),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_39),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_8),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_72),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_105),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_135),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_13),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_86),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_127),
.Y(n_256)
);

NOR2xp67_ASAP7_75t_L g257 ( 
.A(n_59),
.B(n_26),
.Y(n_257)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_76),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_110),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_90),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_143),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_170),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_249),
.Y(n_263)
);

AND2x4_ASAP7_75t_L g264 ( 
.A(n_165),
.B(n_1),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_1),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_258),
.Y(n_266)
);

AO22x1_ASAP7_75t_L g267 ( 
.A1(n_165),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_199),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_258),
.Y(n_269)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_199),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_175),
.B(n_2),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_199),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_249),
.Y(n_273)
);

OAI21x1_ASAP7_75t_L g274 ( 
.A1(n_171),
.A2(n_68),
.B(n_151),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_244),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_199),
.Y(n_277)
);

AND2x4_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_6),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_254),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_158),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_258),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_155),
.Y(n_283)
);

BUFx12f_ASAP7_75t_L g284 ( 
.A(n_170),
.Y(n_284)
);

AND2x6_ASAP7_75t_L g285 ( 
.A(n_159),
.B(n_45),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_157),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_162),
.Y(n_287)
);

OAI22x1_ASAP7_75t_R g288 ( 
.A1(n_167),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_186),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_160),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_163),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_203),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_216),
.A2(n_185),
.B1(n_209),
.B2(n_167),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_202),
.B(n_9),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_170),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_258),
.B(n_203),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_164),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_159),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_169),
.B(n_10),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_204),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_202),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_179),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_203),
.Y(n_303)
);

OA21x2_ASAP7_75t_L g304 ( 
.A1(n_171),
.A2(n_71),
.B(n_149),
.Y(n_304)
);

AND2x4_ASAP7_75t_L g305 ( 
.A(n_191),
.B(n_10),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_166),
.Y(n_306)
);

BUFx12f_ASAP7_75t_L g307 ( 
.A(n_245),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_203),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_258),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_220),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_172),
.B(n_11),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_185),
.Y(n_312)
);

CKINVDCx11_ASAP7_75t_R g313 ( 
.A(n_209),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_255),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_220),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_258),
.Y(n_316)
);

OAI21x1_ASAP7_75t_L g317 ( 
.A1(n_184),
.A2(n_79),
.B(n_148),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_211),
.B(n_14),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_213),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_215),
.Y(n_320)
);

INVx5_ASAP7_75t_L g321 ( 
.A(n_220),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_183),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_220),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_224),
.B(n_16),
.Y(n_324)
);

AND2x4_ASAP7_75t_L g325 ( 
.A(n_191),
.B(n_18),
.Y(n_325)
);

BUFx12f_ASAP7_75t_L g326 ( 
.A(n_245),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_177),
.Y(n_327)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_251),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_255),
.Y(n_329)
);

OAI21x1_ASAP7_75t_L g330 ( 
.A1(n_184),
.A2(n_84),
.B(n_147),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_234),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_204),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_204),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_251),
.B(n_256),
.Y(n_334)
);

OAI21x1_ASAP7_75t_L g335 ( 
.A1(n_234),
.A2(n_83),
.B(n_146),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_268),
.Y(n_336)
);

BUFx10_ASAP7_75t_L g337 ( 
.A(n_301),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_278),
.A2(n_231),
.B1(n_204),
.B2(n_225),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_268),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_266),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_278),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_301),
.B(n_248),
.Y(n_342)
);

NAND3xp33_ASAP7_75t_L g343 ( 
.A(n_281),
.B(n_193),
.C(n_190),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_262),
.B(n_248),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_266),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_286),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_278),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_268),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_290),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_286),
.B(n_188),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_295),
.B(n_210),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_269),
.Y(n_352)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_285),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_276),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_276),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_282),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_263),
.A2(n_228),
.B1(n_242),
.B2(n_250),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_282),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_309),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_262),
.B(n_168),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_309),
.Y(n_361)
);

AND2x4_ASAP7_75t_L g362 ( 
.A(n_305),
.B(n_257),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_316),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_316),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_331),
.Y(n_365)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_285),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_268),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_284),
.B(n_290),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_268),
.Y(n_369)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_264),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_334),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_272),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_294),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_289),
.B(n_201),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_302),
.B(n_322),
.Y(n_375)
);

AOI21x1_ASAP7_75t_L g376 ( 
.A1(n_296),
.A2(n_252),
.B(n_200),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_284),
.B(n_156),
.Y(n_377)
);

NOR3xp33_ASAP7_75t_L g378 ( 
.A(n_319),
.B(n_230),
.C(n_226),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_331),
.Y(n_379)
);

AND3x2_ASAP7_75t_L g380 ( 
.A(n_273),
.B(n_205),
.C(n_195),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_272),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_302),
.B(n_173),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_322),
.B(n_174),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_264),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_281),
.B(n_206),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_287),
.B(n_291),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_272),
.Y(n_387)
);

OAI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_265),
.A2(n_178),
.B1(n_247),
.B2(n_232),
.Y(n_388)
);

NAND3xp33_ASAP7_75t_L g389 ( 
.A(n_287),
.B(n_218),
.C(n_260),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_291),
.B(n_176),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_327),
.B(n_180),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g392 ( 
.A(n_283),
.B(n_256),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_300),
.Y(n_393)
);

BUFx8_ASAP7_75t_SL g394 ( 
.A(n_329),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_277),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_327),
.B(n_181),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_297),
.B(n_207),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_264),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_292),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_305),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_285),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_271),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_328),
.B(n_182),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_300),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_306),
.B(n_187),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_332),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_305),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_303),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_325),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_307),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_308),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_332),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_332),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_333),
.Y(n_414)
);

NAND3xp33_ASAP7_75t_L g415 ( 
.A(n_311),
.B(n_324),
.C(n_318),
.Y(n_415)
);

INVx2_ASAP7_75t_SL g416 ( 
.A(n_325),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_308),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_308),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_325),
.B(n_307),
.Y(n_419)
);

OAI22xp33_ASAP7_75t_L g420 ( 
.A1(n_314),
.A2(n_221),
.B1(n_229),
.B2(n_253),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_328),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_333),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_308),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_299),
.A2(n_233),
.B1(n_237),
.B2(n_240),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_308),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_326),
.Y(n_426)
);

NOR2xp67_ASAP7_75t_L g427 ( 
.A(n_410),
.B(n_326),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_402),
.B(n_298),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_371),
.B(n_298),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_371),
.B(n_320),
.Y(n_430)
);

OR2x2_ASAP7_75t_L g431 ( 
.A(n_349),
.B(n_312),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_419),
.B(n_279),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_353),
.B(n_189),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_353),
.B(n_192),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_375),
.B(n_293),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_366),
.B(n_329),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_405),
.B(n_373),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_366),
.B(n_288),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_366),
.B(n_252),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_390),
.B(n_280),
.Y(n_440)
);

NAND2xp33_ASAP7_75t_L g441 ( 
.A(n_416),
.B(n_400),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_366),
.B(n_194),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_346),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_391),
.B(n_275),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_396),
.B(n_275),
.Y(n_445)
);

AO21x2_ASAP7_75t_L g446 ( 
.A1(n_376),
.A2(n_335),
.B(n_330),
.Y(n_446)
);

NOR3xp33_ASAP7_75t_L g447 ( 
.A(n_420),
.B(n_267),
.C(n_313),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_365),
.Y(n_448)
);

NOR2xp67_ASAP7_75t_L g449 ( 
.A(n_392),
.B(n_333),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_415),
.B(n_197),
.Y(n_450)
);

OAI22xp33_ASAP7_75t_L g451 ( 
.A1(n_424),
.A2(n_267),
.B1(n_304),
.B2(n_246),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_375),
.A2(n_350),
.B1(n_415),
.B2(n_416),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_392),
.B(n_198),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_386),
.B(n_208),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_341),
.Y(n_455)
);

AND2x2_ASAP7_75t_SL g456 ( 
.A(n_346),
.B(n_304),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_350),
.B(n_313),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_351),
.B(n_196),
.Y(n_458)
);

OAI22xp33_ASAP7_75t_L g459 ( 
.A1(n_424),
.A2(n_304),
.B1(n_212),
.B2(n_222),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_401),
.B(n_214),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_401),
.B(n_217),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_401),
.A2(n_330),
.B(n_317),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_362),
.B(n_219),
.Y(n_463)
);

O2A1O1Ixp33_ASAP7_75t_L g464 ( 
.A1(n_388),
.A2(n_378),
.B(n_347),
.C(n_357),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_365),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_347),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g467 ( 
.A(n_426),
.B(n_18),
.Y(n_467)
);

A2O1A1Ixp33_ASAP7_75t_L g468 ( 
.A1(n_347),
.A2(n_335),
.B(n_274),
.C(n_317),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_362),
.B(n_223),
.Y(n_469)
);

AOI221xp5_ASAP7_75t_L g470 ( 
.A1(n_388),
.A2(n_259),
.B1(n_235),
.B2(n_238),
.C(n_241),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_379),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_382),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_421),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_362),
.B(n_383),
.Y(n_474)
);

NAND3xp33_ASAP7_75t_L g475 ( 
.A(n_338),
.B(n_227),
.C(n_239),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_360),
.B(n_344),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_337),
.B(n_161),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_370),
.B(n_270),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_370),
.A2(n_261),
.B1(n_236),
.B2(n_270),
.Y(n_479)
);

NOR3xp33_ASAP7_75t_L g480 ( 
.A(n_368),
.B(n_19),
.C(n_20),
.Y(n_480)
);

NOR3xp33_ASAP7_75t_L g481 ( 
.A(n_343),
.B(n_20),
.C(n_21),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_342),
.B(n_236),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_337),
.B(n_21),
.Y(n_483)
);

INVxp33_ASAP7_75t_L g484 ( 
.A(n_394),
.Y(n_484)
);

NAND2xp33_ASAP7_75t_L g485 ( 
.A(n_400),
.B(n_261),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_L g486 ( 
.A1(n_400),
.A2(n_261),
.B1(n_321),
.B2(n_270),
.Y(n_486)
);

INVx2_ASAP7_75t_SL g487 ( 
.A(n_380),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_384),
.B(n_398),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_374),
.B(n_261),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_407),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_407),
.B(n_409),
.Y(n_491)
);

INVx4_ASAP7_75t_L g492 ( 
.A(n_407),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_409),
.A2(n_321),
.B1(n_323),
.B2(n_315),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_385),
.A2(n_321),
.B1(n_323),
.B2(n_315),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_377),
.B(n_22),
.Y(n_495)
);

OR2x6_ASAP7_75t_L g496 ( 
.A(n_389),
.B(n_310),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_403),
.B(n_321),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_397),
.B(n_310),
.Y(n_498)
);

OAI22xp33_ASAP7_75t_L g499 ( 
.A1(n_340),
.A2(n_323),
.B1(n_315),
.B2(n_25),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_472),
.B(n_345),
.Y(n_500)
);

NAND2x1p5_ASAP7_75t_L g501 ( 
.A(n_490),
.B(n_345),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_431),
.Y(n_502)
);

A2O1A1Ixp33_ASAP7_75t_L g503 ( 
.A1(n_491),
.A2(n_352),
.B(n_354),
.C(n_355),
.Y(n_503)
);

OAI321xp33_ASAP7_75t_L g504 ( 
.A1(n_451),
.A2(n_315),
.A3(n_323),
.B1(n_376),
.B2(n_354),
.C(n_363),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_437),
.B(n_452),
.Y(n_505)
);

INVx4_ASAP7_75t_L g506 ( 
.A(n_466),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_462),
.A2(n_363),
.B(n_352),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_476),
.B(n_359),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_441),
.A2(n_361),
.B(n_359),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_443),
.Y(n_510)
);

NOR2x1p5_ASAP7_75t_SL g511 ( 
.A(n_473),
.B(n_356),
.Y(n_511)
);

O2A1O1Ixp33_ASAP7_75t_L g512 ( 
.A1(n_464),
.A2(n_361),
.B(n_364),
.C(n_356),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_476),
.B(n_428),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_468),
.A2(n_358),
.B(n_406),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_439),
.A2(n_406),
.B(n_404),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_458),
.B(n_393),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_488),
.A2(n_456),
.B(n_478),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_453),
.B(n_22),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_458),
.B(n_393),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_438),
.A2(n_404),
.B1(n_412),
.B2(n_422),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_448),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_474),
.B(n_23),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_456),
.A2(n_412),
.B(n_413),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_449),
.B(n_414),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_432),
.B(n_422),
.Y(n_525)
);

A2O1A1Ixp33_ASAP7_75t_L g526 ( 
.A1(n_491),
.A2(n_425),
.B(n_339),
.C(n_418),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_435),
.B(n_25),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_447),
.A2(n_425),
.B1(n_339),
.B2(n_418),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_465),
.Y(n_529)
);

O2A1O1Ixp33_ASAP7_75t_SL g530 ( 
.A1(n_451),
.A2(n_395),
.B(n_367),
.C(n_369),
.Y(n_530)
);

AOI21xp33_ASAP7_75t_L g531 ( 
.A1(n_450),
.A2(n_26),
.B(n_28),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_492),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_432),
.B(n_28),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_457),
.B(n_30),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_447),
.A2(n_336),
.B1(n_417),
.B2(n_411),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_430),
.B(n_30),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_440),
.B(n_31),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_463),
.B(n_32),
.Y(n_538)
);

AO21x1_ASAP7_75t_L g539 ( 
.A1(n_459),
.A2(n_336),
.B(n_348),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_429),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_444),
.B(n_32),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_436),
.B(n_423),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_445),
.B(n_33),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_470),
.B(n_34),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_427),
.B(n_35),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_471),
.B(n_37),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_495),
.B(n_38),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_455),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_496),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_454),
.B(n_40),
.Y(n_550)
);

A2O1A1Ixp33_ASAP7_75t_L g551 ( 
.A1(n_482),
.A2(n_372),
.B(n_417),
.C(n_411),
.Y(n_551)
);

A2O1A1Ixp33_ASAP7_75t_L g552 ( 
.A1(n_482),
.A2(n_372),
.B(n_411),
.C(n_408),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_469),
.B(n_40),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_483),
.B(n_47),
.Y(n_554)
);

A2O1A1Ixp33_ASAP7_75t_L g555 ( 
.A1(n_489),
.A2(n_399),
.B(n_387),
.C(n_381),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_467),
.Y(n_556)
);

A2O1A1Ixp33_ASAP7_75t_L g557 ( 
.A1(n_481),
.A2(n_497),
.B(n_475),
.C(n_480),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_477),
.B(n_48),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_480),
.B(n_49),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_487),
.B(n_50),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_498),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_481),
.A2(n_387),
.B1(n_381),
.B2(n_423),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_L g563 ( 
.A1(n_433),
.A2(n_387),
.B(n_381),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_496),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_496),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_486),
.B(n_423),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_486),
.B(n_423),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_446),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_434),
.B(n_442),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_460),
.B(n_54),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_479),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_461),
.A2(n_61),
.B1(n_62),
.B2(n_65),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_499),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_505),
.B(n_485),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_500),
.B(n_493),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_547),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_501),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_501),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_502),
.B(n_484),
.Y(n_579)
);

OAI21xp5_ASAP7_75t_L g580 ( 
.A1(n_517),
.A2(n_494),
.B(n_70),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_513),
.B(n_67),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_527),
.B(n_540),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_502),
.B(n_92),
.Y(n_583)
);

AO31x2_ASAP7_75t_L g584 ( 
.A1(n_503),
.A2(n_93),
.A3(n_95),
.B(n_98),
.Y(n_584)
);

OA22x2_ASAP7_75t_L g585 ( 
.A1(n_547),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_585)
);

OAI21xp5_ASAP7_75t_L g586 ( 
.A1(n_523),
.A2(n_117),
.B(n_118),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_510),
.B(n_123),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_525),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_537),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_549),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_544),
.B(n_522),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_545),
.Y(n_592)
);

AO21x1_ASAP7_75t_L g593 ( 
.A1(n_559),
.A2(n_566),
.B(n_567),
.Y(n_593)
);

INVx5_ASAP7_75t_L g594 ( 
.A(n_549),
.Y(n_594)
);

O2A1O1Ixp5_ASAP7_75t_L g595 ( 
.A1(n_557),
.A2(n_518),
.B(n_553),
.C(n_538),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_508),
.B(n_533),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_564),
.Y(n_597)
);

AOI221xp5_ASAP7_75t_L g598 ( 
.A1(n_556),
.A2(n_531),
.B1(n_528),
.B2(n_536),
.C(n_512),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_556),
.B(n_554),
.Y(n_599)
);

AOI221xp5_ASAP7_75t_SL g600 ( 
.A1(n_541),
.A2(n_543),
.B1(n_550),
.B2(n_571),
.C(n_546),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_L g601 ( 
.A1(n_504),
.A2(n_562),
.B(n_526),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_548),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_L g603 ( 
.A1(n_554),
.A2(n_564),
.B1(n_529),
.B2(n_521),
.Y(n_603)
);

A2O1A1Ixp33_ASAP7_75t_L g604 ( 
.A1(n_569),
.A2(n_519),
.B(n_516),
.C(n_511),
.Y(n_604)
);

AO31x2_ASAP7_75t_L g605 ( 
.A1(n_555),
.A2(n_551),
.A3(n_552),
.B(n_530),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_509),
.A2(n_515),
.B(n_563),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_521),
.B(n_529),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_L g608 ( 
.A1(n_521),
.A2(n_565),
.B1(n_558),
.B2(n_506),
.Y(n_608)
);

OAI21xp5_ASAP7_75t_SL g609 ( 
.A1(n_520),
.A2(n_572),
.B(n_524),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_532),
.B(n_561),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_SL g611 ( 
.A1(n_560),
.A2(n_570),
.B(n_535),
.Y(n_611)
);

AOI21x1_ASAP7_75t_L g612 ( 
.A1(n_539),
.A2(n_542),
.B(n_462),
.Y(n_612)
);

OAI21x1_ASAP7_75t_SL g613 ( 
.A1(n_505),
.A2(n_506),
.B(n_539),
.Y(n_613)
);

NAND3xp33_ASAP7_75t_L g614 ( 
.A(n_557),
.B(n_562),
.C(n_480),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_540),
.Y(n_615)
);

OAI21x1_ASAP7_75t_L g616 ( 
.A1(n_568),
.A2(n_514),
.B(n_507),
.Y(n_616)
);

INVx4_ASAP7_75t_L g617 ( 
.A(n_501),
.Y(n_617)
);

OAI21x1_ASAP7_75t_SL g618 ( 
.A1(n_505),
.A2(n_506),
.B(n_539),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_501),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_L g620 ( 
.A1(n_505),
.A2(n_573),
.B1(n_547),
.B2(n_554),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_540),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_500),
.B(n_513),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_500),
.B(n_513),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_505),
.A2(n_573),
.B1(n_547),
.B2(n_554),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_510),
.Y(n_625)
);

OAI21x1_ASAP7_75t_L g626 ( 
.A1(n_568),
.A2(n_514),
.B(n_507),
.Y(n_626)
);

NAND3xp33_ASAP7_75t_SL g627 ( 
.A(n_502),
.B(n_329),
.C(n_447),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_502),
.Y(n_628)
);

NAND2x1p5_ASAP7_75t_L g629 ( 
.A(n_502),
.B(n_431),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_500),
.B(n_513),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_540),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_540),
.B(n_534),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_500),
.B(n_513),
.Y(n_633)
);

OR2x6_ASAP7_75t_L g634 ( 
.A(n_547),
.B(n_457),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_547),
.A2(n_447),
.B1(n_527),
.B2(n_513),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_501),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_500),
.B(n_513),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_540),
.B(n_534),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_505),
.B(n_513),
.Y(n_639)
);

BUFx8_ASAP7_75t_L g640 ( 
.A(n_547),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_540),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_540),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_501),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_547),
.Y(n_644)
);

NAND2x1p5_ASAP7_75t_L g645 ( 
.A(n_502),
.B(n_431),
.Y(n_645)
);

INVxp67_ASAP7_75t_L g646 ( 
.A(n_502),
.Y(n_646)
);

OAI21xp33_ASAP7_75t_SL g647 ( 
.A1(n_514),
.A2(n_456),
.B(n_541),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_547),
.A2(n_447),
.B1(n_527),
.B2(n_513),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_500),
.B(n_513),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_510),
.B(n_436),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_620),
.A2(n_624),
.B1(n_635),
.B2(n_648),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_615),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_602),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_621),
.Y(n_654)
);

AOI221xp5_ASAP7_75t_L g655 ( 
.A1(n_622),
.A2(n_633),
.B1(n_637),
.B2(n_649),
.C(n_623),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_631),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_646),
.B(n_641),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_617),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_640),
.Y(n_659)
);

OAI221xp5_ASAP7_75t_L g660 ( 
.A1(n_635),
.A2(n_648),
.B1(n_630),
.B2(n_634),
.C(n_582),
.Y(n_660)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_577),
.Y(n_661)
);

A2O1A1Ixp33_ASAP7_75t_L g662 ( 
.A1(n_595),
.A2(n_639),
.B(n_620),
.C(n_624),
.Y(n_662)
);

AO31x2_ASAP7_75t_L g663 ( 
.A1(n_593),
.A2(n_606),
.A3(n_604),
.B(n_608),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_617),
.B(n_619),
.Y(n_664)
);

OAI22xp5_ASAP7_75t_L g665 ( 
.A1(n_639),
.A2(n_599),
.B1(n_577),
.B2(n_578),
.Y(n_665)
);

A2O1A1Ixp33_ASAP7_75t_L g666 ( 
.A1(n_647),
.A2(n_600),
.B(n_591),
.C(n_614),
.Y(n_666)
);

CKINVDCx6p67_ASAP7_75t_R g667 ( 
.A(n_625),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_619),
.Y(n_668)
);

AOI31xp67_ASAP7_75t_L g669 ( 
.A1(n_585),
.A2(n_607),
.A3(n_581),
.B(n_574),
.Y(n_669)
);

INVx11_ASAP7_75t_L g670 ( 
.A(n_640),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_636),
.B(n_643),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_642),
.B(n_629),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_636),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_588),
.B(n_632),
.Y(n_674)
);

BUFx2_ASAP7_75t_R g675 ( 
.A(n_628),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_594),
.Y(n_676)
);

INVxp67_ASAP7_75t_L g677 ( 
.A(n_645),
.Y(n_677)
);

OAI22xp5_ASAP7_75t_L g678 ( 
.A1(n_599),
.A2(n_578),
.B1(n_634),
.B2(n_603),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_643),
.Y(n_679)
);

AO21x2_ASAP7_75t_L g680 ( 
.A1(n_580),
.A2(n_614),
.B(n_586),
.Y(n_680)
);

OAI21xp5_ASAP7_75t_L g681 ( 
.A1(n_596),
.A2(n_647),
.B(n_575),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_632),
.B(n_638),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_594),
.Y(n_683)
);

OA21x2_ASAP7_75t_L g684 ( 
.A1(n_611),
.A2(n_609),
.B(n_598),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_627),
.A2(n_634),
.B1(n_589),
.B2(n_638),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_576),
.B(n_644),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_592),
.A2(n_650),
.B1(n_583),
.B2(n_610),
.Y(n_687)
);

BUFx2_ASAP7_75t_R g688 ( 
.A(n_587),
.Y(n_688)
);

NAND2x1p5_ASAP7_75t_L g689 ( 
.A(n_594),
.B(n_590),
.Y(n_689)
);

AO21x2_ASAP7_75t_L g690 ( 
.A1(n_605),
.A2(n_584),
.B(n_597),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_579),
.B(n_597),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_SL g692 ( 
.A1(n_584),
.A2(n_624),
.B(n_620),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_615),
.Y(n_693)
);

OAI21xp5_ASAP7_75t_L g694 ( 
.A1(n_595),
.A2(n_623),
.B(n_622),
.Y(n_694)
);

CKINVDCx11_ASAP7_75t_R g695 ( 
.A(n_634),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_640),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_617),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_646),
.B(n_502),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_640),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_620),
.A2(n_624),
.B1(n_648),
.B2(n_635),
.Y(n_700)
);

OAI21x1_ASAP7_75t_SL g701 ( 
.A1(n_620),
.A2(n_624),
.B(n_603),
.Y(n_701)
);

AO21x2_ASAP7_75t_L g702 ( 
.A1(n_613),
.A2(n_618),
.B(n_601),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_617),
.Y(n_703)
);

HB1xp67_ASAP7_75t_L g704 ( 
.A(n_577),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_640),
.Y(n_705)
);

AOI221xp5_ASAP7_75t_L g706 ( 
.A1(n_622),
.A2(n_420),
.B1(n_633),
.B2(n_630),
.C(n_623),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_640),
.Y(n_707)
);

OAI21x1_ASAP7_75t_L g708 ( 
.A1(n_612),
.A2(n_626),
.B(n_616),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_620),
.A2(n_624),
.B1(n_447),
.B2(n_591),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_620),
.A2(n_624),
.B1(n_447),
.B2(n_591),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_620),
.A2(n_624),
.B1(n_447),
.B2(n_591),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_622),
.B(n_623),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_640),
.Y(n_713)
);

OAI21xp5_ASAP7_75t_L g714 ( 
.A1(n_595),
.A2(n_623),
.B(n_622),
.Y(n_714)
);

OAI22xp5_ASAP7_75t_L g715 ( 
.A1(n_709),
.A2(n_710),
.B1(n_711),
.B2(n_660),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_SL g716 ( 
.A1(n_651),
.A2(n_700),
.B1(n_701),
.B2(n_678),
.Y(n_716)
);

INVx1_ASAP7_75t_SL g717 ( 
.A(n_667),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_709),
.A2(n_710),
.B1(n_711),
.B2(n_655),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_694),
.B(n_714),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_653),
.B(n_681),
.Y(n_720)
);

INVxp67_ASAP7_75t_SL g721 ( 
.A(n_661),
.Y(n_721)
);

HB1xp67_ASAP7_75t_L g722 ( 
.A(n_698),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_653),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_652),
.Y(n_724)
);

BUFx12f_ASAP7_75t_L g725 ( 
.A(n_659),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_654),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_706),
.B(n_712),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_656),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_693),
.Y(n_729)
);

HB1xp67_ASAP7_75t_L g730 ( 
.A(n_661),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_666),
.Y(n_731)
);

OR2x2_ASAP7_75t_L g732 ( 
.A(n_704),
.B(n_684),
.Y(n_732)
);

BUFx12f_ASAP7_75t_L g733 ( 
.A(n_659),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_672),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_662),
.Y(n_735)
);

OR2x6_ASAP7_75t_L g736 ( 
.A(n_692),
.B(n_665),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_674),
.B(n_682),
.Y(n_737)
);

OAI21xp5_ASAP7_75t_L g738 ( 
.A1(n_685),
.A2(n_669),
.B(n_687),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_657),
.B(n_691),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_702),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_687),
.A2(n_685),
.B1(n_695),
.B2(n_682),
.Y(n_741)
);

INVx3_ASAP7_75t_SL g742 ( 
.A(n_664),
.Y(n_742)
);

OAI222xp33_ASAP7_75t_L g743 ( 
.A1(n_707),
.A2(n_658),
.B1(n_703),
.B2(n_668),
.C1(n_697),
.C2(n_677),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_690),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_684),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_658),
.Y(n_746)
);

INVxp67_ASAP7_75t_L g747 ( 
.A(n_675),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_671),
.B(n_668),
.Y(n_748)
);

CKINVDCx20_ASAP7_75t_R g749 ( 
.A(n_707),
.Y(n_749)
);

CKINVDCx6p67_ASAP7_75t_R g750 ( 
.A(n_742),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_720),
.Y(n_751)
);

CKINVDCx11_ASAP7_75t_R g752 ( 
.A(n_749),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_723),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_742),
.Y(n_754)
);

BUFx3_ASAP7_75t_L g755 ( 
.A(n_742),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_732),
.B(n_663),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_727),
.B(n_737),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_745),
.B(n_663),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_745),
.B(n_663),
.Y(n_759)
);

CKINVDCx20_ASAP7_75t_R g760 ( 
.A(n_725),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_719),
.B(n_716),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_736),
.B(n_663),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_741),
.B(n_695),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_736),
.B(n_708),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_730),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_731),
.B(n_680),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_725),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_721),
.Y(n_768)
);

BUFx2_ASAP7_75t_L g769 ( 
.A(n_736),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_753),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_750),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_754),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_751),
.B(n_722),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_751),
.B(n_719),
.Y(n_774)
);

INVxp67_ASAP7_75t_L g775 ( 
.A(n_768),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_761),
.A2(n_715),
.B1(n_718),
.B2(n_736),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_750),
.Y(n_777)
);

OR2x2_ASAP7_75t_L g778 ( 
.A(n_768),
.B(n_739),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_758),
.B(n_740),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_762),
.B(n_736),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_765),
.B(n_735),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_758),
.B(n_740),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_752),
.B(n_717),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_766),
.B(n_735),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_758),
.B(n_744),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_774),
.B(n_759),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_770),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_774),
.B(n_759),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_781),
.B(n_756),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_780),
.B(n_764),
.Y(n_790)
);

INVxp67_ASAP7_75t_SL g791 ( 
.A(n_775),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_785),
.B(n_759),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_785),
.B(n_762),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_778),
.B(n_765),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_778),
.B(n_761),
.Y(n_795)
);

NOR2x1p5_ASAP7_75t_L g796 ( 
.A(n_771),
.B(n_750),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_784),
.B(n_766),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_784),
.B(n_766),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_779),
.B(n_762),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_773),
.B(n_757),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_794),
.B(n_781),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_786),
.B(n_775),
.Y(n_802)
);

OAI31xp33_ASAP7_75t_L g803 ( 
.A1(n_796),
.A2(n_743),
.A3(n_763),
.B(n_776),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_786),
.B(n_788),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_788),
.B(n_779),
.Y(n_805)
);

O2A1O1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_800),
.A2(n_747),
.B(n_763),
.C(n_738),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_792),
.B(n_782),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_787),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_792),
.B(n_782),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_790),
.B(n_780),
.Y(n_810)
);

NAND2x1_ASAP7_75t_L g811 ( 
.A(n_790),
.B(n_772),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_795),
.B(n_797),
.Y(n_812)
);

AOI222xp33_ASAP7_75t_L g813 ( 
.A1(n_802),
.A2(n_757),
.B1(n_791),
.B2(n_812),
.C1(n_783),
.C2(n_804),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_808),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_808),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_801),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_801),
.Y(n_817)
);

INVx1_ASAP7_75t_SL g818 ( 
.A(n_807),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_803),
.A2(n_780),
.B1(n_769),
.B2(n_762),
.Y(n_819)
);

AOI21xp33_ASAP7_75t_L g820 ( 
.A1(n_806),
.A2(n_726),
.B(n_724),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_804),
.B(n_789),
.Y(n_821)
);

AOI32xp33_ASAP7_75t_L g822 ( 
.A1(n_807),
.A2(n_777),
.A3(n_771),
.B1(n_793),
.B2(n_799),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_809),
.B(n_805),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_814),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_819),
.A2(n_780),
.B1(n_790),
.B2(n_769),
.Y(n_825)
);

OAI221xp5_ASAP7_75t_L g826 ( 
.A1(n_822),
.A2(n_811),
.B1(n_789),
.B2(n_797),
.C(n_798),
.Y(n_826)
);

OAI21xp33_ASAP7_75t_SL g827 ( 
.A1(n_813),
.A2(n_818),
.B(n_823),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_821),
.Y(n_828)
);

OAI32xp33_ASAP7_75t_L g829 ( 
.A1(n_820),
.A2(n_771),
.A3(n_777),
.B1(n_755),
.B2(n_754),
.Y(n_829)
);

OAI21xp33_ASAP7_75t_L g830 ( 
.A1(n_827),
.A2(n_820),
.B(n_817),
.Y(n_830)
);

AOI211x1_ASAP7_75t_L g831 ( 
.A1(n_826),
.A2(n_829),
.B(n_816),
.C(n_805),
.Y(n_831)
);

AOI21xp33_ASAP7_75t_L g832 ( 
.A1(n_824),
.A2(n_699),
.B(n_696),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_830),
.B(n_824),
.Y(n_833)
);

NOR3xp33_ASAP7_75t_L g834 ( 
.A(n_832),
.B(n_752),
.C(n_713),
.Y(n_834)
);

NOR2xp67_ASAP7_75t_L g835 ( 
.A(n_833),
.B(n_767),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_834),
.B(n_831),
.Y(n_836)
);

NOR2x1_ASAP7_75t_L g837 ( 
.A(n_835),
.B(n_760),
.Y(n_837)
);

NOR2xp67_ASAP7_75t_L g838 ( 
.A(n_836),
.B(n_733),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_837),
.B(n_760),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_838),
.Y(n_840)
);

AND2x4_ASAP7_75t_SL g841 ( 
.A(n_839),
.B(n_840),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_839),
.Y(n_842)
);

XNOR2xp5_ASAP7_75t_L g843 ( 
.A(n_839),
.B(n_705),
.Y(n_843)
);

XNOR2xp5_ASAP7_75t_L g844 ( 
.A(n_843),
.B(n_670),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_842),
.Y(n_845)
);

OAI221xp5_ASAP7_75t_L g846 ( 
.A1(n_841),
.A2(n_825),
.B1(n_733),
.B2(n_811),
.C(n_777),
.Y(n_846)
);

AOI221xp5_ASAP7_75t_L g847 ( 
.A1(n_842),
.A2(n_828),
.B1(n_724),
.B2(n_726),
.C(n_728),
.Y(n_847)
);

OAI21xp5_ASAP7_75t_L g848 ( 
.A1(n_842),
.A2(n_676),
.B(n_683),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_845),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_R g850 ( 
.A(n_844),
.B(n_686),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_847),
.B(n_815),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_848),
.B(n_728),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_846),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_844),
.A2(n_796),
.B1(n_688),
.B2(n_810),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_845),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_855),
.B(n_849),
.Y(n_856)
);

AOI21x1_ASAP7_75t_L g857 ( 
.A1(n_853),
.A2(n_734),
.B(n_729),
.Y(n_857)
);

OAI211xp5_ASAP7_75t_L g858 ( 
.A1(n_850),
.A2(n_697),
.B(n_679),
.C(n_673),
.Y(n_858)
);

OR2x6_ASAP7_75t_L g859 ( 
.A(n_854),
.B(n_689),
.Y(n_859)
);

OA21x2_ASAP7_75t_L g860 ( 
.A1(n_856),
.A2(n_851),
.B(n_852),
.Y(n_860)
);

AND3x1_ASAP7_75t_L g861 ( 
.A(n_857),
.B(n_748),
.C(n_746),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_860),
.A2(n_859),
.B(n_861),
.Y(n_862)
);

BUFx24_ASAP7_75t_SL g863 ( 
.A(n_862),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_863),
.A2(n_858),
.B1(n_810),
.B2(n_809),
.Y(n_864)
);


endmodule