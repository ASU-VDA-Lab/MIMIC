module fake_jpeg_2765_n_415 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_415);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_415;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_14),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_49),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_16),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_50),
.B(n_61),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_51),
.Y(n_136)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_54),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_18),
.B(n_14),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_83),
.Y(n_102)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_56),
.Y(n_143)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

BUFx4f_ASAP7_75t_SL g59 ( 
.A(n_23),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_59),
.Y(n_131)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_25),
.B(n_13),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

NAND2xp33_ASAP7_75t_SL g65 ( 
.A(n_29),
.B(n_0),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_79),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_72),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_75),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

AOI21xp33_ASAP7_75t_L g116 ( 
.A1(n_76),
.A2(n_87),
.B(n_47),
.Y(n_116)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_25),
.B(n_14),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_42),
.B(n_13),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_80),
.B(n_39),
.Y(n_129)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_31),
.B(n_0),
.C(n_1),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_17),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_88),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_90),
.Y(n_122)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_1),
.Y(n_145)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_93),
.Y(n_105)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_95),
.Y(n_110)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_62),
.A2(n_40),
.B1(n_19),
.B2(n_27),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_100),
.A2(n_113),
.B1(n_70),
.B2(n_64),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_94),
.A2(n_46),
.B1(n_44),
.B2(n_36),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_101),
.A2(n_138),
.B1(n_54),
.B2(n_68),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_66),
.A2(n_41),
.B1(n_37),
.B2(n_34),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_104),
.A2(n_73),
.B1(n_84),
.B2(n_86),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_71),
.A2(n_21),
.B1(n_41),
.B2(n_28),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_59),
.B(n_28),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_114),
.B(n_123),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_116),
.B(n_118),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_59),
.A2(n_34),
.B(n_37),
.C(n_21),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_51),
.B(n_39),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_129),
.B(n_133),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_91),
.B(n_27),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_85),
.A2(n_46),
.B1(n_44),
.B2(n_36),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_52),
.B(n_19),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_75),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_89),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_147),
.B(n_150),
.Y(n_215)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_146),
.Y(n_148)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_149),
.Y(n_198)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_151),
.Y(n_206)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_146),
.Y(n_152)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_152),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_74),
.B1(n_46),
.B2(n_67),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_153),
.A2(n_106),
.B1(n_130),
.B2(n_139),
.Y(n_203)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_108),
.Y(n_154)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_154),
.Y(n_197)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_155),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_102),
.B(n_78),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_159),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_157),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_158),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_118),
.B(n_72),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_107),
.Y(n_161)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_122),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_162),
.B(n_166),
.Y(n_211)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_99),
.Y(n_164)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_164),
.Y(n_209)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_122),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_108),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_167),
.B(n_171),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_168),
.A2(n_175),
.B1(n_178),
.B2(n_182),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_121),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_170),
.B(n_174),
.Y(n_200)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_172),
.Y(n_191)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_124),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_110),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_176),
.B(n_183),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_98),
.B(n_63),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_180),
.Y(n_195)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_L g179 ( 
.A1(n_100),
.A2(n_95),
.B1(n_92),
.B2(n_68),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_179),
.A2(n_187),
.B1(n_137),
.B2(n_135),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_98),
.B(n_96),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_140),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_105),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_124),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_184),
.A2(n_186),
.B1(n_188),
.B2(n_120),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_130),
.Y(n_196)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_97),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_121),
.A2(n_87),
.B1(n_22),
.B2(n_24),
.Y(n_188)
);

O2A1O1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_159),
.A2(n_131),
.B(n_140),
.C(n_109),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_193),
.A2(n_218),
.B(n_185),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_194),
.A2(n_203),
.B1(n_187),
.B2(n_182),
.Y(n_222)
);

NAND3xp33_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_158),
.C(n_160),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_96),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_152),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_213),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_176),
.A2(n_179),
.B1(n_183),
.B2(n_177),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_217),
.A2(n_182),
.B1(n_148),
.B2(n_172),
.Y(n_223)
);

AO22x1_ASAP7_75t_L g218 ( 
.A1(n_181),
.A2(n_144),
.B1(n_139),
.B2(n_143),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_173),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_221),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_189),
.A2(n_181),
.B1(n_180),
.B2(n_185),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_220),
.A2(n_237),
.B1(n_238),
.B2(n_203),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_222),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_223),
.Y(n_250)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_224),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_193),
.A2(n_181),
.B(n_189),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_225),
.A2(n_230),
.B(n_218),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_226),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_201),
.A2(n_169),
.B1(n_111),
.B2(n_115),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_227),
.A2(n_231),
.B1(n_222),
.B2(n_234),
.Y(n_252)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_232),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_195),
.B(n_211),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_212),
.C(n_216),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_193),
.A2(n_178),
.B(n_163),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_195),
.A2(n_111),
.B1(n_171),
.B2(n_165),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_127),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_235),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_208),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_239),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_204),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_161),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_191),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_194),
.A2(n_112),
.B1(n_99),
.B2(n_144),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_215),
.A2(n_112),
.B1(n_143),
.B2(n_164),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_208),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_200),
.B(n_149),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_241),
.B(n_216),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_243),
.A2(n_248),
.B(n_246),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_225),
.A2(n_215),
.B1(n_205),
.B2(n_196),
.Y(n_247)
);

AO22x1_ASAP7_75t_SL g273 ( 
.A1(n_247),
.A2(n_237),
.B1(n_238),
.B2(n_235),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_226),
.A2(n_218),
.B(n_197),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_248),
.A2(n_239),
.B(n_240),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_197),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_249),
.B(n_254),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_255),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_236),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_263),
.Y(n_275)
);

MAJx2_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_207),
.C(n_212),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_220),
.B(n_207),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_226),
.A2(n_230),
.B1(n_221),
.B2(n_227),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_256),
.A2(n_223),
.B1(n_232),
.B2(n_228),
.Y(n_266)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_257),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_259),
.B(n_219),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_191),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_262),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_241),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_262),
.Y(n_265)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_265),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_266),
.A2(n_278),
.B1(n_257),
.B2(n_260),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_259),
.Y(n_267)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_267),
.Y(n_296)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_269),
.A2(n_277),
.B(n_280),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_273),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_231),
.Y(n_272)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_272),
.Y(n_303)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_276),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_247),
.A2(n_235),
.B1(n_224),
.B2(n_199),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_253),
.B(n_244),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_281),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_243),
.A2(n_233),
.B(n_199),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_235),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_251),
.Y(n_282)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_282),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_258),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_254),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_190),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_286),
.A2(n_291),
.B1(n_206),
.B2(n_214),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_261),
.C(n_255),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_299),
.C(n_277),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_261),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_280),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_268),
.A2(n_260),
.B1(n_245),
.B2(n_246),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_290),
.A2(n_292),
.B1(n_294),
.B2(n_301),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_270),
.A2(n_244),
.B1(n_245),
.B2(n_242),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_276),
.A2(n_258),
.B1(n_250),
.B2(n_255),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_264),
.A2(n_242),
.B1(n_254),
.B2(n_249),
.Y(n_294)
);

OAI21x1_ASAP7_75t_L g326 ( 
.A1(n_295),
.A2(n_273),
.B(n_204),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_284),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_202),
.C(n_198),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_264),
.A2(n_224),
.B1(n_209),
.B2(n_198),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_284),
.A2(n_209),
.B1(n_206),
.B2(n_202),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_305),
.A2(n_266),
.B1(n_267),
.B2(n_265),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_293),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_307),
.B(n_308),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_309),
.B(n_319),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_284),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_310),
.B(n_311),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_292),
.B(n_283),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_312),
.B(n_302),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_275),
.Y(n_313)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_313),
.Y(n_332)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_314),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_287),
.B(n_279),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_315),
.B(n_297),
.Y(n_340)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_306),
.Y(n_316)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_316),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_318),
.A2(n_328),
.B1(n_303),
.B2(n_288),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_294),
.B(n_275),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_293),
.B(n_271),
.Y(n_320)
);

INVxp33_ASAP7_75t_L g330 ( 
.A(n_320),
.Y(n_330)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_306),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_321),
.B(n_323),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_299),
.B(n_269),
.C(n_282),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_322),
.B(n_325),
.Y(n_344)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_300),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_303),
.B(n_281),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_324),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_298),
.B(n_272),
.C(n_273),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_326),
.B(n_327),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_290),
.B(n_273),
.C(n_186),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_309),
.B(n_302),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_333),
.B(n_338),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_334),
.A2(n_317),
.B1(n_327),
.B2(n_313),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_318),
.A2(n_317),
.B1(n_288),
.B2(n_325),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_336),
.A2(n_337),
.B1(n_210),
.B2(n_190),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_310),
.B(n_297),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_340),
.B(n_348),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_315),
.B(n_304),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_346),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_308),
.Y(n_347)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_347),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_319),
.B(n_304),
.Y(n_348)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_351),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_331),
.A2(n_320),
.B1(n_324),
.B2(n_322),
.Y(n_352)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_356),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_330),
.A2(n_305),
.B(n_311),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_354),
.A2(n_361),
.B(n_335),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_330),
.A2(n_301),
.B1(n_206),
.B2(n_214),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_355),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_332),
.A2(n_210),
.B1(n_155),
.B2(n_157),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_357),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_329),
.B(n_344),
.C(n_346),
.Y(n_358)
);

OR2x2_ASAP7_75t_L g376 ( 
.A(n_358),
.B(n_359),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_345),
.B(n_151),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_340),
.B(n_142),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_360),
.B(n_1),
.Y(n_373)
);

A2O1A1Ixp33_ASAP7_75t_SL g361 ( 
.A1(n_339),
.A2(n_117),
.B(n_126),
.C(n_142),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_342),
.A2(n_126),
.B1(n_97),
.B2(n_117),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_362),
.B(n_341),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_329),
.B(n_106),
.C(n_120),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_363),
.B(n_333),
.C(n_338),
.Y(n_366)
);

XNOR2x1_ASAP7_75t_L g365 ( 
.A(n_358),
.B(n_343),
.Y(n_365)
);

NOR2x1_ASAP7_75t_SL g386 ( 
.A(n_365),
.B(n_361),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_366),
.B(n_369),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_367),
.A2(n_378),
.B1(n_5),
.B2(n_6),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_354),
.A2(n_343),
.B(n_347),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_368),
.A2(n_374),
.B(n_364),
.Y(n_379)
);

OAI221xp5_ASAP7_75t_L g371 ( 
.A1(n_353),
.A2(n_348),
.B1(n_120),
.B2(n_24),
.C(n_5),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_371),
.B(n_377),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_373),
.B(n_361),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_349),
.A2(n_1),
.B(n_2),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_363),
.B(n_2),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_379),
.B(n_389),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_387),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_376),
.A2(n_351),
.B(n_355),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_383),
.A2(n_386),
.B(n_5),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_372),
.A2(n_350),
.B1(n_357),
.B2(n_362),
.Y(n_384)
);

INVxp33_ASAP7_75t_L g395 ( 
.A(n_384),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_375),
.A2(n_370),
.B(n_378),
.Y(n_385)
);

NOR2xp67_ASAP7_75t_SL g391 ( 
.A(n_385),
.B(n_3),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_369),
.B(n_361),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_370),
.B(n_3),
.Y(n_388)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_388),
.Y(n_390)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_391),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_380),
.A2(n_379),
.B(n_385),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_392),
.B(n_8),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_384),
.B(n_3),
.Y(n_394)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_394),
.B(n_8),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_396),
.A2(n_382),
.B(n_7),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_389),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_397),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_399),
.B(n_403),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_395),
.B(n_6),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_400),
.A2(n_401),
.B(n_405),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_404),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_393),
.B(n_398),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_402),
.B(n_397),
.C(n_390),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_408),
.A2(n_10),
.B(n_11),
.Y(n_411)
);

NOR3xp33_ASAP7_75t_L g410 ( 
.A(n_407),
.B(n_399),
.C(n_10),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_410),
.B(n_411),
.C(n_406),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_412),
.B(n_409),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_413),
.A2(n_11),
.B(n_392),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_414),
.B(n_11),
.Y(n_415)
);


endmodule