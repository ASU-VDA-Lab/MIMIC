module fake_jpeg_22100_n_164 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_1),
.B(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_3),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_35),
.B(n_15),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_14),
.B(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_38),
.B(n_16),
.Y(n_66)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_43),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_30),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_30),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_26),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_55),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_21),
.B1(n_26),
.B2(n_19),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_47),
.A2(n_48),
.B1(n_64),
.B2(n_6),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_31),
.A2(n_18),
.B1(n_30),
.B2(n_23),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_68),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_23),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_59),
.Y(n_84)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_37),
.B(n_29),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_63),
.B(n_66),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_21),
.B1(n_19),
.B2(n_27),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_43),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_65),
.A2(n_20),
.B1(n_34),
.B2(n_22),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_28),
.Y(n_67)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_33),
.B(n_20),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_71),
.Y(n_105)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_81),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_32),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_78),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_43),
.C(n_36),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_61),
.C(n_50),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_32),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_36),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_86),
.Y(n_104)
);

AO22x1_ASAP7_75t_L g80 ( 
.A1(n_48),
.A2(n_34),
.B1(n_1),
.B2(n_2),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_80),
.A2(n_69),
.B1(n_54),
.B2(n_13),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_82),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_0),
.Y(n_83)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_1),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_2),
.Y(n_88)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_3),
.Y(n_89)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_90),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_7),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_91),
.B(n_46),
.Y(n_96)
);

AOI221xp5_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_64),
.B1(n_53),
.B2(n_46),
.C(n_52),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_103),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_100),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_73),
.A2(n_50),
.B(n_61),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_77),
.B(n_87),
.Y(n_115)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_107),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_86),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_108),
.A2(n_109),
.B1(n_85),
.B2(n_79),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_72),
.A2(n_8),
.B1(n_10),
.B2(n_13),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_8),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_111),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_121),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_115),
.B(n_93),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_92),
.Y(n_116)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_87),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_123),
.C(n_107),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_74),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_87),
.Y(n_122)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_90),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_75),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_125),
.Y(n_132)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_98),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_117),
.Y(n_137)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_131),
.Y(n_146)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_136),
.C(n_115),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_126),
.A2(n_97),
.B1(n_95),
.B2(n_100),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_135),
.A2(n_130),
.B1(n_131),
.B2(n_129),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_137),
.A2(n_76),
.B1(n_81),
.B2(n_110),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_142),
.Y(n_149)
);

XNOR2x1_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_118),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_136),
.Y(n_148)
);

AO221x1_ASAP7_75t_L g140 ( 
.A1(n_134),
.A2(n_71),
.B1(n_76),
.B2(n_108),
.C(n_123),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_140),
.B(n_141),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_129),
.A2(n_97),
.B1(n_95),
.B2(n_122),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_143),
.B(n_127),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_135),
.B(n_125),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_119),
.C(n_118),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_139),
.C(n_144),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_145),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_152),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_153),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_154),
.A2(n_157),
.B(n_147),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_146),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_155),
.A2(n_99),
.B(n_101),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_141),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_160),
.C(n_101),
.Y(n_162)
);

AOI322xp5_ASAP7_75t_L g161 ( 
.A1(n_158),
.A2(n_156),
.A3(n_155),
.B1(n_148),
.B2(n_138),
.C1(n_109),
.C2(n_99),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_162),
.C(n_120),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_163),
.B(n_84),
.Y(n_164)
);


endmodule