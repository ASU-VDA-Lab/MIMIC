module fake_jpeg_18352_n_233 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_233);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_233;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_SL g13 ( 
.A(n_11),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_36),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_22),
.Y(n_32)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_45),
.B(n_36),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_31),
.A2(n_20),
.B1(n_19),
.B2(n_23),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_34),
.B1(n_32),
.B2(n_28),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_20),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_49),
.Y(n_58)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_16),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_51),
.B(n_63),
.Y(n_80)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g77 ( 
.A(n_53),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_46),
.A2(n_19),
.B1(n_20),
.B2(n_23),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_40),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_38),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_43),
.Y(n_76)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g85 ( 
.A(n_57),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_60),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_33),
.B(n_35),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_61),
.A2(n_47),
.B(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_44),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_17),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_50),
.A2(n_19),
.B1(n_20),
.B2(n_23),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_39),
.A2(n_34),
.B1(n_28),
.B2(n_32),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_29),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_69),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_50),
.A2(n_13),
.B1(n_26),
.B2(n_21),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_14),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_72),
.A2(n_76),
.B(n_82),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_60),
.Y(n_92)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_81),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_42),
.B(n_41),
.C(n_50),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_58),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_83),
.B(n_58),
.Y(n_91)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_84),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_62),
.A2(n_26),
.B1(n_17),
.B2(n_24),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_86),
.A2(n_89),
.B1(n_32),
.B2(n_74),
.Y(n_98)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_87),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_55),
.A2(n_26),
.B1(n_17),
.B2(n_24),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_81),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_101),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_92),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_83),
.B(n_63),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_59),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_72),
.A2(n_61),
.B(n_69),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_107),
.B(n_60),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_98),
.Y(n_109)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_82),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_104),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_70),
.A2(n_56),
.B1(n_55),
.B2(n_41),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_52),
.B(n_51),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_103),
.A2(n_67),
.B(n_79),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_75),
.A2(n_70),
.B1(n_88),
.B2(n_76),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_80),
.B(n_60),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_76),
.Y(n_118)
);

XNOR2x2_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_52),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_128),
.B(n_107),
.Y(n_129)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_105),
.B(n_80),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_115),
.A2(n_119),
.B(n_121),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_75),
.C(n_65),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_126),
.C(n_104),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_118),
.B(n_120),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_59),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_102),
.Y(n_121)
);

XNOR2x1_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_13),
.Y(n_122)
);

XOR2x2_ASAP7_75t_SL g145 ( 
.A(n_122),
.B(n_124),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_85),
.Y(n_123)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

NAND3xp33_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_8),
.C(n_1),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_77),
.C(n_27),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_97),
.Y(n_127)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_128),
.B(n_122),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_116),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_134),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_116),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_97),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_139),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_125),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_136),
.B(n_94),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_125),
.Y(n_138)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_102),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_126),
.C(n_117),
.Y(n_150)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_142),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_109),
.A2(n_92),
.B1(n_108),
.B2(n_99),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_143),
.A2(n_144),
.B1(n_84),
.B2(n_87),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_109),
.A2(n_92),
.B1(n_55),
.B2(n_94),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_114),
.A2(n_64),
.B1(n_54),
.B2(n_85),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_146),
.A2(n_77),
.B1(n_71),
.B2(n_95),
.Y(n_161)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_148),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_146),
.A2(n_113),
.B1(n_119),
.B2(n_121),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_149),
.A2(n_161),
.B1(n_129),
.B2(n_141),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_158),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_152),
.B(n_130),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_132),
.A2(n_119),
.B1(n_115),
.B2(n_127),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_166),
.B1(n_78),
.B2(n_25),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_112),
.C(n_118),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_157),
.C(n_162),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_112),
.C(n_106),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_106),
.Y(n_158)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_160),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_77),
.C(n_85),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_149),
.A2(n_137),
.B1(n_144),
.B2(n_143),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_167),
.A2(n_169),
.B1(n_175),
.B2(n_176),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_177),
.Y(n_190)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_174),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_164),
.A2(n_145),
.B1(n_131),
.B2(n_147),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_152),
.A2(n_145),
.B1(n_37),
.B2(n_78),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_14),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_25),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_179),
.Y(n_191)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_181),
.B(n_16),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_180),
.A2(n_157),
.B(n_156),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_185),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_171),
.A2(n_163),
.B(n_153),
.Y(n_184)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_153),
.C(n_158),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_194),
.C(n_170),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_160),
.B1(n_37),
.B2(n_25),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_181),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_176),
.A2(n_160),
.B1(n_1),
.B2(n_2),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_18),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_16),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_177),
.C(n_172),
.Y(n_194)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_195),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_187),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_197),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_15),
.C(n_27),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_199),
.C(n_202),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_15),
.C(n_27),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_200),
.A2(n_204),
.B1(n_18),
.B2(n_1),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_15),
.C(n_27),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_201),
.A2(n_186),
.B1(n_182),
.B2(n_189),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_209),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_195),
.A2(n_185),
.B1(n_193),
.B2(n_190),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_203),
.A2(n_190),
.B1(n_24),
.B2(n_18),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_211),
.Y(n_215)
);

OAI21x1_ASAP7_75t_L g211 ( 
.A1(n_196),
.A2(n_14),
.B(n_2),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_205),
.A2(n_37),
.B(n_3),
.Y(n_213)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_213),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_205),
.A2(n_8),
.B(n_3),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_216),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_212),
.A2(n_8),
.B(n_3),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_206),
.B(n_6),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_6),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_206),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_220),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_L g225 ( 
.A1(n_223),
.A2(n_218),
.B1(n_6),
.B2(n_7),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_208),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_224),
.A2(n_12),
.B(n_7),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_225),
.A2(n_227),
.B(n_7),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_221),
.C(n_222),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_228),
.B(n_229),
.C(n_9),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_230),
.A2(n_10),
.B1(n_12),
.B2(n_0),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_10),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_10),
.Y(n_233)
);


endmodule