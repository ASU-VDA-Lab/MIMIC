module fake_jpeg_18743_n_110 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_110);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_51),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_58),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_49),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_52),
.A2(n_45),
.B1(n_41),
.B2(n_48),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_38),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_43),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_56),
.A2(n_50),
.B1(n_46),
.B2(n_49),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_65),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_70),
.Y(n_80)
);

INVx5_ASAP7_75t_SL g70 ( 
.A(n_58),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_68),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_71),
.B(n_10),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_40),
.Y(n_72)
);

XOR2x2_ASAP7_75t_SL g85 ( 
.A(n_72),
.B(n_75),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_77),
.Y(n_87)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_0),
.Y(n_75)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_60),
.B(n_1),
.C(n_3),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_78),
.A2(n_79),
.B1(n_81),
.B2(n_66),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_67),
.A2(n_18),
.B1(n_33),
.B2(n_7),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_12),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_13),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_75),
.B(n_9),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_86),
.A2(n_91),
.B1(n_72),
.B2(n_14),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_80),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_35),
.C(n_16),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_90),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_79),
.B1(n_78),
.B2(n_81),
.Y(n_92)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_85),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_94),
.A2(n_83),
.B(n_89),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_86),
.C(n_87),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

AOI322xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_97),
.A3(n_100),
.B1(n_92),
.B2(n_101),
.C1(n_95),
.C2(n_26),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_103),
.B(n_15),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_20),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_21),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_SL g107 ( 
.A1(n_106),
.A2(n_22),
.B(n_24),
.C(n_27),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_108),
.A2(n_30),
.B(n_32),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_84),
.Y(n_110)
);


endmodule