module fake_jpeg_11576_n_516 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_516);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_516;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_SL g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx8_ASAP7_75t_SL g44 ( 
.A(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_25),
.B(n_17),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_50),
.B(n_70),
.Y(n_122)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_53),
.B(n_64),
.Y(n_99)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_54),
.Y(n_136)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_57),
.Y(n_132)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_58),
.Y(n_143)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_59),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_60),
.Y(n_155)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_61),
.Y(n_151)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_63),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_44),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_65),
.B(n_66),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_18),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_18),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_69),
.B(n_74),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_0),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_25),
.B(n_16),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_72),
.B(n_82),
.Y(n_135)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_32),
.B(n_15),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

NAND2x1_ASAP7_75t_L g81 ( 
.A(n_33),
.B(n_1),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_81),
.A2(n_42),
.B(n_39),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_32),
.B(n_2),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_43),
.B(n_2),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_84),
.B(n_2),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_18),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_97),
.Y(n_129)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_41),
.Y(n_90)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_95),
.Y(n_157)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_18),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_71),
.A2(n_38),
.B1(n_24),
.B2(n_27),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_108),
.A2(n_121),
.B1(n_134),
.B2(n_140),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_55),
.A2(n_46),
.B1(n_30),
.B2(n_37),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_110),
.A2(n_120),
.B1(n_123),
.B2(n_126),
.Y(n_194)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_51),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_115),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_70),
.A2(n_46),
.B1(n_37),
.B2(n_30),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_116),
.A2(n_96),
.B1(n_49),
.B2(n_31),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_59),
.A2(n_27),
.B1(n_49),
.B2(n_31),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_60),
.A2(n_38),
.B1(n_27),
.B2(n_33),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_67),
.A2(n_28),
.B1(n_48),
.B2(n_45),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_75),
.A2(n_28),
.B1(n_48),
.B2(n_45),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_127),
.A2(n_14),
.B(n_5),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_65),
.B(n_43),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_133),
.B(n_152),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_60),
.A2(n_33),
.B1(n_29),
.B2(n_37),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_52),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_137),
.Y(n_190)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_54),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_62),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_98),
.A2(n_29),
.B1(n_46),
.B2(n_30),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_139),
.A2(n_36),
.B1(n_93),
.B2(n_76),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_78),
.A2(n_83),
.B1(n_87),
.B2(n_85),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_77),
.A2(n_29),
.B1(n_46),
.B2(n_37),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_148),
.A2(n_149),
.B1(n_90),
.B2(n_57),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_80),
.A2(n_29),
.B1(n_30),
.B2(n_39),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_65),
.B(n_35),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_156),
.B(n_19),
.Y(n_177)
);

OA22x2_ASAP7_75t_L g159 ( 
.A1(n_116),
.A2(n_81),
.B1(n_61),
.B2(n_89),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_159),
.Y(n_260)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_117),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_160),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_161),
.B(n_169),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_162),
.Y(n_233)
);

AOI21xp33_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_35),
.B(n_20),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_163),
.B(n_164),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_119),
.B(n_95),
.Y(n_164)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_167),
.Y(n_242)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_168),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_92),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_139),
.A2(n_42),
.B1(n_39),
.B2(n_36),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_171),
.A2(n_175),
.B1(n_205),
.B2(n_209),
.Y(n_253)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_106),
.Y(n_172)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_100),
.Y(n_173)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_173),
.Y(n_220)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_112),
.Y(n_174)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_174),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_117),
.A2(n_42),
.B1(n_36),
.B2(n_63),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_107),
.Y(n_176)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_176),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_177),
.B(n_179),
.Y(n_257)
);

BUFx6f_ASAP7_75t_SL g178 ( 
.A(n_124),
.Y(n_178)
);

BUFx4f_ASAP7_75t_SL g225 ( 
.A(n_178),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_99),
.B(n_58),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_101),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_180),
.Y(n_234)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_103),
.Y(n_182)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_182),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_111),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_183),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_122),
.B(n_19),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_184),
.B(n_187),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_185),
.A2(n_186),
.B1(n_199),
.B2(n_212),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_148),
.A2(n_108),
.B1(n_149),
.B2(n_134),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_104),
.B(n_20),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_102),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_188),
.B(n_202),
.Y(n_245)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_105),
.Y(n_189)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_189),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_191),
.A2(n_217),
.B1(n_145),
.B2(n_130),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_105),
.Y(n_192)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_192),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_193),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_236)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_118),
.Y(n_195)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_195),
.Y(n_268)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_114),
.Y(n_196)
);

INVx8_ASAP7_75t_L g255 ( 
.A(n_196),
.Y(n_255)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_107),
.Y(n_197)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_197),
.Y(n_235)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_136),
.Y(n_198)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_198),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_121),
.A2(n_79),
.B1(n_56),
.B2(n_86),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_125),
.B(n_18),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_200),
.A2(n_206),
.B(n_210),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_127),
.Y(n_201)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_128),
.B(n_2),
.Y(n_202)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_114),
.Y(n_203)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_203),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_136),
.B(n_3),
.Y(n_204)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_204),
.Y(n_267)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_146),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_143),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_207),
.B(n_208),
.Y(n_261)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_143),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_144),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_144),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_110),
.A2(n_3),
.B(n_5),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_216),
.C(n_157),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_142),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_150),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_158),
.Y(n_214)
);

OA22x2_ASAP7_75t_L g215 ( 
.A1(n_146),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_215)
);

NAND2x1p5_ASAP7_75t_L g216 ( 
.A(n_109),
.B(n_5),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_109),
.Y(n_217)
);

AO21x1_ASAP7_75t_L g279 ( 
.A1(n_218),
.A2(n_174),
.B(n_162),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_219),
.B(n_228),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_194),
.A2(n_142),
.B1(n_145),
.B2(n_130),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_221),
.A2(n_240),
.B1(n_244),
.B2(n_246),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_170),
.B(n_153),
.C(n_147),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_237),
.B(n_248),
.C(n_249),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_194),
.A2(n_147),
.B1(n_131),
.B2(n_113),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_211),
.A2(n_131),
.B1(n_113),
.B2(n_132),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_191),
.A2(n_132),
.B1(n_155),
.B2(n_8),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_193),
.A2(n_155),
.B1(n_7),
.B2(n_8),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_247),
.A2(n_262),
.B1(n_178),
.B2(n_192),
.Y(n_271)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_184),
.B(n_6),
.C(n_7),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_173),
.B(n_182),
.C(n_206),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_195),
.B(n_159),
.C(n_200),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_250),
.B(n_259),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_159),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_251),
.A2(n_265),
.B1(n_266),
.B2(n_190),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_165),
.B(n_9),
.Y(n_254)
);

XOR2x2_ASAP7_75t_L g285 ( 
.A(n_254),
.B(n_264),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_159),
.B(n_9),
.C(n_10),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_188),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_214),
.B(n_11),
.C(n_13),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_216),
.A2(n_14),
.B1(n_215),
.B2(n_205),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_216),
.A2(n_14),
.B1(n_215),
.B2(n_189),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_260),
.A2(n_215),
.B1(n_203),
.B2(n_196),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_269),
.A2(n_271),
.B1(n_273),
.B2(n_286),
.Y(n_340)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_261),
.Y(n_270)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_270),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_233),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_272),
.B(n_283),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_260),
.A2(n_210),
.B1(n_213),
.B2(n_212),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_275),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_331)
);

OA21x2_ASAP7_75t_L g276 ( 
.A1(n_243),
.A2(n_190),
.B(n_181),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_276),
.A2(n_295),
.B(n_226),
.Y(n_339)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_277),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_240),
.A2(n_217),
.B1(n_208),
.B2(n_207),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_250),
.A2(n_167),
.B1(n_166),
.B2(n_172),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_227),
.B(n_168),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_281),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_234),
.B(n_181),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_282),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_241),
.B(n_176),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_220),
.Y(n_284)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_284),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_263),
.A2(n_197),
.B1(n_198),
.B2(n_160),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_238),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_287),
.B(n_292),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_223),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_289),
.B(n_299),
.Y(n_321)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_268),
.Y(n_290)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_290),
.Y(n_332)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_252),
.Y(n_291)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_291),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_160),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_231),
.B(n_257),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_293),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_294),
.B(n_315),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_228),
.A2(n_219),
.B(n_253),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_262),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_296),
.B(n_300),
.Y(n_338)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_252),
.Y(n_297)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_297),
.Y(n_347)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_222),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_245),
.B(n_249),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_222),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_301),
.B(n_304),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_241),
.B(n_245),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_302),
.Y(n_334)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_242),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_303),
.Y(n_353)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_242),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_235),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_305),
.B(n_307),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_237),
.B(n_254),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_306),
.A2(n_288),
.B(n_281),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_265),
.B(n_266),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_225),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_308),
.A2(n_309),
.B1(n_314),
.B2(n_232),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_225),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_232),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_310),
.B(n_311),
.Y(n_354)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_229),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_229),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_312),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_263),
.A2(n_236),
.B1(n_259),
.B2(n_247),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_313),
.A2(n_285),
.B1(n_283),
.B2(n_296),
.Y(n_350)
);

INVxp33_ASAP7_75t_L g314 ( 
.A(n_226),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_236),
.B(n_251),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_317),
.Y(n_385)
);

AO21x2_ASAP7_75t_SL g322 ( 
.A1(n_307),
.A2(n_244),
.B(n_246),
.Y(n_322)
);

AO22x2_ASAP7_75t_L g369 ( 
.A1(n_322),
.A2(n_319),
.B1(n_323),
.B2(n_331),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_287),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_325),
.B(n_329),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_315),
.A2(n_295),
.B1(n_275),
.B2(n_274),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_326),
.B(n_333),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_294),
.B(n_248),
.C(n_239),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_328),
.B(n_337),
.C(n_343),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_305),
.Y(n_329)
);

OAI32xp33_ASAP7_75t_L g333 ( 
.A1(n_270),
.A2(n_224),
.A3(n_256),
.B1(n_255),
.B2(n_230),
.Y(n_333)
);

AO22x1_ASAP7_75t_L g336 ( 
.A1(n_277),
.A2(n_225),
.B1(n_230),
.B2(n_258),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_336),
.A2(n_339),
.B(n_341),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_298),
.B(n_258),
.C(n_264),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_313),
.A2(n_255),
.B1(n_269),
.B2(n_286),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_278),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_342),
.B(n_323),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_298),
.B(n_288),
.C(n_300),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_346),
.B(n_324),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_285),
.B(n_280),
.C(n_306),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_348),
.B(n_343),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_350),
.A2(n_304),
.B1(n_310),
.B2(n_348),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_273),
.A2(n_271),
.B1(n_279),
.B2(n_289),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_352),
.A2(n_336),
.B(n_321),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_274),
.A2(n_279),
.B1(n_285),
.B2(n_284),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_355),
.B(n_338),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_276),
.A2(n_290),
.B(n_291),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_356),
.A2(n_276),
.B(n_312),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_344),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_357),
.B(n_366),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_358),
.A2(n_360),
.B(n_370),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_322),
.A2(n_301),
.B1(n_311),
.B2(n_303),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_359),
.B(n_362),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_339),
.A2(n_297),
.B(n_299),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_361),
.B(n_364),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_322),
.A2(n_341),
.B1(n_338),
.B2(n_350),
.Y(n_362)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_345),
.Y(n_365)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_365),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_344),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_321),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_367),
.B(n_371),
.Y(n_413)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_369),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_355),
.A2(n_320),
.B(n_326),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_335),
.B(n_351),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_356),
.B(n_316),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_372),
.Y(n_407)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_327),
.Y(n_374)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_374),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_375),
.B(n_364),
.Y(n_410)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_327),
.Y(n_376)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_376),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_377),
.B(n_380),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_354),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_379),
.B(n_369),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_334),
.B(n_318),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_381),
.B(n_387),
.C(n_321),
.Y(n_400)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_332),
.Y(n_382)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_382),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_349),
.A2(n_346),
.B(n_352),
.Y(n_383)
);

AOI21xp33_ASAP7_75t_L g417 ( 
.A1(n_383),
.A2(n_389),
.B(n_390),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_334),
.B(n_318),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_384),
.B(n_391),
.Y(n_403)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_332),
.Y(n_386)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_386),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_324),
.B(n_337),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_349),
.A2(n_340),
.B(n_354),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_388),
.Y(n_393)
);

AOI322xp5_ASAP7_75t_L g389 ( 
.A1(n_319),
.A2(n_322),
.A3(n_328),
.B1(n_340),
.B2(n_333),
.C1(n_353),
.C2(n_330),
.Y(n_389)
);

NAND3xp33_ASAP7_75t_L g390 ( 
.A(n_345),
.B(n_347),
.C(n_353),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_388),
.A2(n_366),
.B1(n_357),
.B2(n_363),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_396),
.B(n_397),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_372),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_400),
.B(n_404),
.C(n_406),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_363),
.A2(n_330),
.B1(n_347),
.B2(n_336),
.Y(n_401)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_401),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_381),
.B(n_373),
.C(n_387),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_373),
.B(n_375),
.C(n_361),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_410),
.B(n_385),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_411),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_379),
.B(n_369),
.Y(n_414)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_414),
.Y(n_445)
);

XOR2x1_ASAP7_75t_L g416 ( 
.A(n_383),
.B(n_370),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_416),
.B(n_378),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_360),
.A2(n_369),
.B1(n_358),
.B2(n_362),
.Y(n_418)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_418),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_368),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_419),
.B(n_402),
.Y(n_441)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_374),
.Y(n_420)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_420),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_415),
.A2(n_378),
.B(n_391),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_421),
.A2(n_435),
.B(n_439),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_404),
.B(n_372),
.C(n_359),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_423),
.B(n_430),
.C(n_398),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_419),
.B(n_380),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_424),
.B(n_428),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_425),
.B(n_431),
.Y(n_455)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_394),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_426),
.B(n_394),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_413),
.B(n_376),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_400),
.B(n_382),
.C(n_386),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_406),
.B(n_369),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_432),
.B(n_433),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_410),
.B(n_385),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_415),
.A2(n_365),
.B(n_407),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_408),
.Y(n_436)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_436),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_396),
.Y(n_437)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_437),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_407),
.B(n_418),
.Y(n_439)
);

FAx1_ASAP7_75t_SL g440 ( 
.A(n_416),
.B(n_414),
.CI(n_411),
.CON(n_440),
.SN(n_440)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_440),
.B(n_397),
.Y(n_450)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_441),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_408),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_442),
.B(n_444),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_402),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_445),
.A2(n_403),
.B(n_392),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_448),
.A2(n_434),
.B(n_426),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_427),
.A2(n_405),
.B1(n_393),
.B2(n_401),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_449),
.B(n_458),
.Y(n_478)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_450),
.Y(n_469)
);

NOR3xp33_ASAP7_75t_SL g451 ( 
.A(n_436),
.B(n_403),
.C(n_417),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_451),
.B(n_463),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_429),
.Y(n_454)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_454),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_456),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_427),
.A2(n_405),
.B1(n_393),
.B2(n_395),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_443),
.B(n_413),
.Y(n_459)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_459),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_429),
.A2(n_395),
.B1(n_392),
.B2(n_398),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_461),
.B(n_447),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_462),
.B(n_430),
.C(n_422),
.Y(n_466)
);

NOR3xp33_ASAP7_75t_L g463 ( 
.A(n_439),
.B(n_399),
.C(n_409),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_438),
.B(n_399),
.Y(n_465)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_465),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_466),
.B(n_467),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_462),
.B(n_422),
.C(n_423),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_455),
.B(n_431),
.C(n_435),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_468),
.B(n_472),
.Y(n_492)
);

A2O1A1Ixp33_ASAP7_75t_SL g470 ( 
.A1(n_447),
.A2(n_421),
.B(n_439),
.C(n_440),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_470),
.A2(n_454),
.B1(n_465),
.B2(n_457),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_471),
.B(n_461),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_455),
.B(n_425),
.C(n_443),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_453),
.B(n_440),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_473),
.B(n_479),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_464),
.B(n_432),
.Y(n_479)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_480),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_481),
.B(n_446),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_482),
.B(n_487),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_483),
.A2(n_471),
.B(n_478),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_485),
.B(n_491),
.Y(n_497)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_480),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_469),
.A2(n_449),
.B1(n_452),
.B2(n_458),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_488),
.B(n_489),
.Y(n_502)
);

OAI211xp5_ASAP7_75t_L g489 ( 
.A1(n_476),
.A2(n_451),
.B(n_448),
.C(n_456),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_468),
.B(n_460),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_475),
.A2(n_460),
.B1(n_433),
.B2(n_426),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_493),
.A2(n_470),
.B1(n_434),
.B2(n_420),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_483),
.A2(n_467),
.B(n_466),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_494),
.B(n_498),
.Y(n_504)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_495),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_484),
.B(n_474),
.Y(n_496)
);

AOI21xp33_ASAP7_75t_L g505 ( 
.A1(n_496),
.A2(n_501),
.B(n_486),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_490),
.A2(n_472),
.B(n_477),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_492),
.B(n_478),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_500),
.B(n_485),
.C(n_491),
.Y(n_507)
);

BUFx4f_ASAP7_75t_SL g503 ( 
.A(n_496),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_503),
.B(n_499),
.Y(n_508)
);

AOI31xp33_ASAP7_75t_L g509 ( 
.A1(n_505),
.A2(n_502),
.A3(n_497),
.B(n_493),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_507),
.B(n_470),
.C(n_409),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_508),
.B(n_509),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_510),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_512),
.B(n_504),
.C(n_506),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_513),
.A2(n_511),
.B(n_503),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_514),
.A2(n_412),
.B(n_470),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_515),
.B(n_412),
.Y(n_516)
);


endmodule