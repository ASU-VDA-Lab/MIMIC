module real_aes_10983_n_16 (n_13, n_4, n_0, n_3, n_5, n_2, n_15, n_7, n_8, n_6, n_9, n_12, n_1, n_14, n_10, n_11, n_16);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_15;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_14;
input n_10;
input n_11;
output n_16;
wire n_17;
wire n_28;
wire n_22;
wire n_24;
wire n_41;
wire n_34;
wire n_19;
wire n_40;
wire n_49;
wire n_46;
wire n_53;
wire n_25;
wire n_47;
wire n_48;
wire n_43;
wire n_32;
wire n_30;
wire n_37;
wire n_51;
wire n_54;
wire n_35;
wire n_42;
wire n_45;
wire n_39;
wire n_27;
wire n_23;
wire n_38;
wire n_50;
wire n_29;
wire n_20;
wire n_52;
wire n_44;
wire n_26;
wire n_18;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
NOR2xp33_ASAP7_75t_R g23 ( .A(n_0), .B(n_5), .Y(n_23) );
NOR3xp33_ASAP7_75t_SL g21 ( .A(n_1), .B(n_8), .C(n_22), .Y(n_21) );
NOR3xp33_ASAP7_75t_SL g43 ( .A(n_1), .B(n_12), .C(n_44), .Y(n_43) );
NAND2xp33_ASAP7_75t_R g22 ( .A(n_2), .B(n_23), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g46 ( .A(n_2), .Y(n_46) );
CKINVDCx5p33_ASAP7_75t_R g24 ( .A(n_3), .Y(n_24) );
NOR4xp25_ASAP7_75t_SL g41 ( .A(n_3), .B(n_42), .C(n_45), .D(n_46), .Y(n_41) );
NOR4xp25_ASAP7_75t_SL g19 ( .A(n_4), .B(n_20), .C(n_24), .D(n_25), .Y(n_19) );
CKINVDCx5p33_ASAP7_75t_R g45 ( .A(n_4), .Y(n_45) );
CKINVDCx5p33_ASAP7_75t_R g32 ( .A(n_6), .Y(n_32) );
NOR2xp33_ASAP7_75t_R g18 ( .A(n_7), .B(n_13), .Y(n_18) );
NAND2xp33_ASAP7_75t_SL g29 ( .A(n_7), .B(n_30), .Y(n_29) );
NOR2xp33_ASAP7_75t_R g36 ( .A(n_7), .B(n_30), .Y(n_36) );
NAND2xp33_ASAP7_75t_R g38 ( .A(n_7), .B(n_13), .Y(n_38) );
CKINVDCx5p33_ASAP7_75t_R g47 ( .A(n_8), .Y(n_47) );
AOI221xp5_ASAP7_75t_R g33 ( .A1(n_9), .A2(n_14), .B1(n_34), .B2(n_37), .C(n_39), .Y(n_33) );
CKINVDCx5p33_ASAP7_75t_R g48 ( .A(n_10), .Y(n_48) );
HB1xp67_ASAP7_75t_L g54 ( .A(n_11), .Y(n_54) );
CKINVDCx5p33_ASAP7_75t_R g25 ( .A(n_12), .Y(n_25) );
CKINVDCx5p33_ASAP7_75t_R g30 ( .A(n_13), .Y(n_30) );
CKINVDCx5p33_ASAP7_75t_R g26 ( .A(n_15), .Y(n_26) );
OAI221xp5_ASAP7_75t_L g16 ( .A1(n_17), .A2(n_26), .B1(n_27), .B2(n_32), .C(n_33), .Y(n_16) );
NAND2xp33_ASAP7_75t_R g17 ( .A(n_18), .B(n_19), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g52 ( .A(n_18), .Y(n_52) );
CKINVDCx5p33_ASAP7_75t_R g31 ( .A(n_19), .Y(n_31) );
NAND2xp33_ASAP7_75t_R g35 ( .A(n_19), .B(n_36), .Y(n_35) );
CKINVDCx5p33_ASAP7_75t_R g20 ( .A(n_21), .Y(n_20) );
CKINVDCx5p33_ASAP7_75t_R g44 ( .A(n_23), .Y(n_44) );
INVxp33_ASAP7_75t_L g27 ( .A(n_28), .Y(n_27) );
NOR2xp33_ASAP7_75t_R g28 ( .A(n_29), .B(n_31), .Y(n_28) );
NOR2xp33_ASAP7_75t_R g37 ( .A(n_31), .B(n_38), .Y(n_37) );
CKINVDCx5p33_ASAP7_75t_R g34 ( .A(n_35), .Y(n_34) );
CKINVDCx5p33_ASAP7_75t_R g49 ( .A(n_36), .Y(n_49) );
OAI32xp33_ASAP7_75t_L g39 ( .A1(n_40), .A2(n_48), .A3(n_49), .B1(n_50), .B2(n_53), .Y(n_39) );
NOR2xp33_ASAP7_75t_R g51 ( .A(n_40), .B(n_52), .Y(n_51) );
NAND2xp33_ASAP7_75t_R g40 ( .A(n_41), .B(n_47), .Y(n_40) );
CKINVDCx5p33_ASAP7_75t_R g42 ( .A(n_43), .Y(n_42) );
CKINVDCx5p33_ASAP7_75t_R g50 ( .A(n_51), .Y(n_50) );
INVx1_ASAP7_75t_L g53 ( .A(n_54), .Y(n_53) );
endmodule