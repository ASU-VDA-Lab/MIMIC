module fake_netlist_6_1892_n_504 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_504);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_504;

wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_209;
wire n_367;
wire n_465;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_342;
wire n_358;
wire n_449;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_495;
wire n_350;
wire n_392;
wire n_442;
wire n_480;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_389;
wire n_415;
wire n_230;
wire n_461;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_372;
wire n_468;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_375;
wire n_338;
wire n_466;
wire n_360;
wire n_235;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_428;
wire n_432;
wire n_167;
wire n_174;
wire n_491;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_493;
wire n_397;
wire n_445;
wire n_425;
wire n_454;
wire n_218;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_172;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_185;
wire n_348;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_456;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_455;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_503;
wire n_321;
wire n_331;
wire n_227;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_357;
wire n_264;
wire n_263;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_477;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_243;
wire n_282;
wire n_436;
wire n_211;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_240;
wire n_319;
wire n_273;
wire n_311;
wire n_403;
wire n_253;
wire n_249;
wire n_201;
wire n_386;
wire n_162;
wire n_487;
wire n_241;
wire n_275;
wire n_276;
wire n_441;
wire n_221;
wire n_444;
wire n_423;
wire n_318;
wire n_303;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_277;
wire n_418;
wire n_199;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_453;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_257;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_489;
wire n_205;
wire n_251;
wire n_301;
wire n_274;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_422;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_187;
wire n_501;
wire n_361;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

INVxp67_ASAP7_75t_L g161 ( 
.A(n_40),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_154),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_1),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_81),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_2),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_97),
.Y(n_168)
);

INVxp67_ASAP7_75t_SL g169 ( 
.A(n_32),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_89),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_146),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_65),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

INVxp33_ASAP7_75t_SL g174 ( 
.A(n_117),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_16),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_4),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_28),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_100),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_83),
.Y(n_180)
);

INVxp33_ASAP7_75t_SL g181 ( 
.A(n_27),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_121),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_68),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_42),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_143),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_116),
.Y(n_186)
);

INVxp67_ASAP7_75t_SL g187 ( 
.A(n_133),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_61),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_151),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_124),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_70),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_73),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_72),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_122),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_6),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_144),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_129),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_86),
.Y(n_198)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_85),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_75),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_49),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_160),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_136),
.Y(n_203)
);

INVxp33_ASAP7_75t_SL g204 ( 
.A(n_45),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_38),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_48),
.Y(n_206)
);

INVxp33_ASAP7_75t_L g207 ( 
.A(n_141),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_113),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_130),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_74),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_54),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_59),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_29),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_60),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_147),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_15),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_3),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_79),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_80),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_35),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_20),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_135),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_138),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_9),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_50),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_125),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_18),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_87),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_123),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_67),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_64),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_39),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_71),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_155),
.Y(n_234)
);

INVxp67_ASAP7_75t_SL g235 ( 
.A(n_41),
.Y(n_235)
);

BUFx2_ASAP7_75t_SL g236 ( 
.A(n_137),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_5),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_12),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_84),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_55),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_119),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_8),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_91),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_101),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_19),
.Y(n_245)
);

INVxp67_ASAP7_75t_SL g246 ( 
.A(n_1),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_52),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_148),
.Y(n_248)
);

INVxp67_ASAP7_75t_SL g249 ( 
.A(n_26),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_90),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_109),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_24),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_134),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_31),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_10),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_76),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_47),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_110),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_145),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_150),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_158),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_30),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_157),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_82),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_153),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_102),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_77),
.Y(n_267)
);

INVxp67_ASAP7_75t_SL g268 ( 
.A(n_132),
.Y(n_268)
);

INVxp67_ASAP7_75t_SL g269 ( 
.A(n_7),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_131),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_149),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_112),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_58),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_105),
.Y(n_274)
);

INVxp67_ASAP7_75t_SL g275 ( 
.A(n_106),
.Y(n_275)
);

INVxp67_ASAP7_75t_SL g276 ( 
.A(n_95),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_69),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_152),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_11),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_13),
.Y(n_280)
);

INVxp33_ASAP7_75t_L g281 ( 
.A(n_43),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_51),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_36),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_173),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_167),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_165),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_168),
.Y(n_287)
);

NAND2xp33_ASAP7_75t_R g288 ( 
.A(n_170),
.B(n_0),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_163),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_171),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_182),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_183),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_186),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_191),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_219),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_164),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_223),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_225),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_229),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_238),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_245),
.Y(n_301)
);

AOI21x1_ASAP7_75t_L g302 ( 
.A1(n_166),
.A2(n_94),
.B(n_156),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_248),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_246),
.A2(n_0),
.B1(n_2),
.B2(n_14),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_196),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_251),
.Y(n_306)
);

NAND2xp33_ASAP7_75t_R g307 ( 
.A(n_252),
.B(n_17),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_257),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_202),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_212),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_259),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_262),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_271),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_272),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_277),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_228),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_265),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_172),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_174),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_162),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_181),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_198),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_175),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_204),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_176),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_267),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_274),
.B(n_21),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_236),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_247),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_177),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_178),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_179),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_R g333 ( 
.A(n_184),
.B(n_22),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_237),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_185),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_207),
.B(n_23),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_188),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_R g338 ( 
.A(n_190),
.B(n_192),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_R g339 ( 
.A(n_193),
.B(n_25),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_194),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_335),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_286),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_286),
.Y(n_343)
);

AND2x4_ASAP7_75t_SL g344 ( 
.A(n_320),
.B(n_180),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_284),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_322),
.B(n_169),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_284),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_326),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_289),
.Y(n_349)
);

AO22x2_ASAP7_75t_L g350 ( 
.A1(n_327),
.A2(n_240),
.B1(n_161),
.B2(n_243),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_334),
.A2(n_281),
.B1(n_243),
.B2(n_240),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_330),
.A2(n_273),
.B1(n_260),
.B2(n_241),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_296),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_323),
.Y(n_354)
);

AND2x2_ASAP7_75t_SL g355 ( 
.A(n_336),
.B(n_189),
.Y(n_355)
);

AO22x2_ASAP7_75t_L g356 ( 
.A1(n_325),
.A2(n_161),
.B1(n_200),
.B2(n_214),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_284),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_332),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_285),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_287),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_328),
.B(n_329),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_290),
.B(n_195),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_340),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_340),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_291),
.B(n_197),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_304),
.A2(n_209),
.B1(n_282),
.B2(n_280),
.Y(n_366)
);

NAND2xp33_ASAP7_75t_L g367 ( 
.A(n_318),
.B(n_283),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_319),
.A2(n_276),
.B1(n_275),
.B2(n_269),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_292),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_293),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_294),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_331),
.Y(n_372)
);

AND2x4_ASAP7_75t_L g373 ( 
.A(n_295),
.B(n_187),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_297),
.B(n_298),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_299),
.B(n_300),
.Y(n_375)
);

AO22x2_ASAP7_75t_L g376 ( 
.A1(n_288),
.A2(n_205),
.B1(n_278),
.B2(n_270),
.Y(n_376)
);

AO22x2_ASAP7_75t_L g377 ( 
.A1(n_337),
.A2(n_201),
.B1(n_266),
.B2(n_264),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_301),
.Y(n_378)
);

O2A1O1Ixp33_ASAP7_75t_L g379 ( 
.A1(n_342),
.A2(n_218),
.B(n_203),
.C(n_279),
.Y(n_379)
);

NAND2xp33_ASAP7_75t_SL g380 ( 
.A(n_366),
.B(n_321),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_345),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_361),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_347),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_343),
.A2(n_199),
.B(n_235),
.Y(n_384)
);

A2O1A1Ixp33_ASAP7_75t_L g385 ( 
.A1(n_355),
.A2(n_217),
.B(n_222),
.C(n_221),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_R g386 ( 
.A(n_378),
.B(n_316),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_359),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_369),
.B(n_303),
.Y(n_388)
);

A2O1A1Ixp33_ASAP7_75t_L g389 ( 
.A1(n_352),
.A2(n_213),
.B(n_215),
.C(n_216),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_349),
.Y(n_390)
);

A2O1A1Ixp33_ASAP7_75t_L g391 ( 
.A1(n_351),
.A2(n_211),
.B(n_210),
.C(n_208),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_372),
.B(n_306),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_353),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_376),
.A2(n_324),
.B1(n_308),
.B2(n_313),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_376),
.A2(n_350),
.B1(n_374),
.B2(n_360),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_375),
.B(n_311),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_371),
.B(n_312),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_362),
.B(n_314),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_365),
.B(n_315),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_354),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_346),
.B(n_249),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_341),
.Y(n_402)
);

OR2x6_ASAP7_75t_L g403 ( 
.A(n_348),
.B(n_206),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_357),
.Y(n_404)
);

A2O1A1Ixp33_ASAP7_75t_L g405 ( 
.A1(n_358),
.A2(n_254),
.B(n_224),
.C(n_226),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_401),
.A2(n_367),
.B(n_373),
.Y(n_406)
);

AO21x2_ASAP7_75t_L g407 ( 
.A1(n_398),
.A2(n_302),
.B(n_333),
.Y(n_407)
);

AOI221xp5_ASAP7_75t_L g408 ( 
.A1(n_391),
.A2(n_350),
.B1(n_368),
.B2(n_377),
.C(n_338),
.Y(n_408)
);

OA21x2_ASAP7_75t_L g409 ( 
.A1(n_385),
.A2(n_364),
.B(n_363),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_382),
.A2(n_370),
.B1(n_317),
.B2(n_305),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_381),
.Y(n_411)
);

AOI22xp33_ASAP7_75t_L g412 ( 
.A1(n_395),
.A2(n_356),
.B1(n_253),
.B2(n_250),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_390),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_399),
.B(n_356),
.Y(n_414)
);

OAI21x1_ASAP7_75t_L g415 ( 
.A1(n_384),
.A2(n_242),
.B(n_227),
.Y(n_415)
);

OAI21x1_ASAP7_75t_L g416 ( 
.A1(n_393),
.A2(n_244),
.B(n_230),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_387),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_390),
.Y(n_418)
);

OR2x6_ASAP7_75t_L g419 ( 
.A(n_403),
.B(n_258),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_402),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_400),
.Y(n_421)
);

NAND2x1p5_ASAP7_75t_L g422 ( 
.A(n_388),
.B(n_255),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_383),
.Y(n_423)
);

AOI21x1_ASAP7_75t_L g424 ( 
.A1(n_392),
.A2(n_256),
.B(n_231),
.Y(n_424)
);

BUFx8_ASAP7_75t_SL g425 ( 
.A(n_403),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_386),
.Y(n_426)
);

OAI21x1_ASAP7_75t_L g427 ( 
.A1(n_379),
.A2(n_239),
.B(n_232),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_397),
.A2(n_268),
.B(n_220),
.Y(n_428)
);

NOR3xp33_ASAP7_75t_SL g429 ( 
.A(n_410),
.B(n_380),
.C(n_394),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_426),
.Y(n_430)
);

OR2x2_ASAP7_75t_L g431 ( 
.A(n_414),
.B(n_396),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_L g432 ( 
.A1(n_409),
.A2(n_233),
.B1(n_234),
.B2(n_261),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_421),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_417),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_413),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_418),
.B(n_404),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_411),
.B(n_310),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_425),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_420),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_SL g440 ( 
.A1(n_422),
.A2(n_309),
.B1(n_344),
.B2(n_339),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g441 ( 
.A(n_412),
.B(n_389),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_409),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_419),
.B(n_263),
.Y(n_443)
);

OR2x6_ASAP7_75t_L g444 ( 
.A(n_419),
.B(n_405),
.Y(n_444)
);

AO31x2_ASAP7_75t_L g445 ( 
.A1(n_428),
.A2(n_307),
.A3(n_34),
.B(n_37),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_423),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_R g447 ( 
.A(n_424),
.B(n_33),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_L g448 ( 
.A1(n_408),
.A2(n_44),
.B1(n_46),
.B2(n_53),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_433),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_431),
.B(n_406),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_434),
.Y(n_451)
);

AOI22xp33_ASAP7_75t_L g452 ( 
.A1(n_448),
.A2(n_441),
.B1(n_439),
.B2(n_444),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_442),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_443),
.Y(n_454)
);

OAI22xp33_ASAP7_75t_L g455 ( 
.A1(n_435),
.A2(n_423),
.B1(n_424),
.B2(n_407),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_436),
.Y(n_456)
);

OA21x2_ASAP7_75t_L g457 ( 
.A1(n_432),
.A2(n_415),
.B(n_416),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_445),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_437),
.B(n_427),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_444),
.A2(n_56),
.B(n_57),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_445),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_446),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_454),
.B(n_429),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_462),
.B(n_440),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_453),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_449),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_451),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_456),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_459),
.B(n_430),
.Y(n_469)
);

NAND3xp33_ASAP7_75t_L g470 ( 
.A(n_452),
.B(n_438),
.C(n_447),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_450),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_455),
.B(n_159),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_461),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_460),
.B(n_62),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_463),
.B(n_464),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_471),
.B(n_458),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_466),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_465),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_468),
.B(n_457),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_467),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_475),
.B(n_469),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_480),
.B(n_470),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_477),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_478),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_476),
.A2(n_472),
.B(n_473),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_479),
.B(n_474),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_484),
.B(n_473),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_481),
.B(n_474),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_482),
.B(n_63),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_483),
.B(n_486),
.Y(n_490)
);

NAND3xp33_ASAP7_75t_SL g491 ( 
.A(n_489),
.B(n_485),
.C(n_78),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_490),
.Y(n_492)
);

OAI211xp5_ASAP7_75t_SL g493 ( 
.A1(n_487),
.A2(n_66),
.B(n_88),
.C(n_92),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_492),
.B(n_488),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_491),
.B(n_93),
.Y(n_495)
);

AOI221xp5_ASAP7_75t_SL g496 ( 
.A1(n_493),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.C(n_104),
.Y(n_496)
);

NAND2xp33_ASAP7_75t_R g497 ( 
.A(n_495),
.B(n_107),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_494),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_498),
.A2(n_496),
.B(n_497),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_498),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_SL g501 ( 
.A1(n_499),
.A2(n_457),
.B1(n_111),
.B2(n_114),
.Y(n_501)
);

OAI22xp33_ASAP7_75t_SL g502 ( 
.A1(n_501),
.A2(n_500),
.B1(n_120),
.B2(n_126),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_502),
.A2(n_108),
.B1(n_128),
.B2(n_139),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_503),
.A2(n_140),
.B(n_142),
.Y(n_504)
);


endmodule