module fake_jpeg_2804_n_154 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_154);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_154;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_24),
.B(n_10),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_SL g53 ( 
.A(n_11),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_9),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_63),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_51),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_56),
.Y(n_65)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_60),
.B(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_64),
.B(n_66),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_68),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_55),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_59),
.B1(n_46),
.B2(n_49),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_53),
.B1(n_54),
.B2(n_43),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_50),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_62),
.B(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_74),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_46),
.Y(n_74)
);

AO22x1_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_46),
.B1(n_53),
.B2(n_43),
.Y(n_76)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_86),
.B1(n_39),
.B2(n_37),
.Y(n_100)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_70),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_80),
.B(n_84),
.Y(n_103)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_70),
.A2(n_73),
.B1(n_74),
.B2(n_41),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_70),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_72),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_34),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_41),
.B1(n_73),
.B2(n_75),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_67),
.A2(n_52),
.B1(n_44),
.B2(n_45),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_45),
.B(n_1),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_76),
.A2(n_45),
.B1(n_1),
.B2(n_2),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_94),
.B1(n_96),
.B2(n_101),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_76),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_19),
.C(n_38),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_31),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_85),
.A2(n_87),
.B1(n_81),
.B2(n_79),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_102),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_82),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_4),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_6),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_105),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_109),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_6),
.B(n_7),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_7),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_8),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_115),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_28),
.B1(n_27),
.B2(n_26),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_99),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_8),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_117),
.B(n_121),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_9),
.B(n_10),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_118),
.A2(n_15),
.B(n_16),
.Y(n_131)
);

BUFx24_ASAP7_75t_SL g119 ( 
.A(n_103),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_123),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_11),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_100),
.A2(n_12),
.B(n_13),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_96),
.B(n_12),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_20),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_21),
.C(n_23),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_110),
.C(n_111),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_120),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_127),
.A2(n_131),
.B1(n_120),
.B2(n_122),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_133),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_112),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_22),
.B(n_25),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_114),
.Y(n_136)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_140),
.Y(n_142)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_134),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_138),
.A2(n_141),
.B1(n_127),
.B2(n_135),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_118),
.C(n_108),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_144),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_143),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_145),
.A2(n_139),
.B(n_130),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_139),
.B(n_146),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_146),
.Y(n_149)
);

INVxp33_ASAP7_75t_L g150 ( 
.A(n_149),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_126),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_129),
.C(n_125),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_142),
.C(n_131),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_153),
.B(n_142),
.Y(n_154)
);


endmodule