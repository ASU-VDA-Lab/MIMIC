module fake_jpeg_20822_n_153 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_153);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_153;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_14),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_6),
.Y(n_64)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_41),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_12),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx8_ASAP7_75t_SL g74 ( 
.A(n_11),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_2),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_79),
.Y(n_84)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_3),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_82),
.Y(n_86)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_78),
.A2(n_74),
.B1(n_48),
.B2(n_73),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_88),
.B1(n_90),
.B2(n_57),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_80),
.B(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_87),
.B(n_91),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_77),
.A2(n_74),
.B1(n_73),
.B2(n_49),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_61),
.B1(n_60),
.B2(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_62),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_87),
.A2(n_86),
.B(n_93),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_99),
.Y(n_110)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_89),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_102),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_59),
.B1(n_67),
.B2(n_61),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_66),
.B(n_70),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_97),
.A2(n_21),
.B1(n_43),
.B2(n_42),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_58),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_63),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_56),
.Y(n_114)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_72),
.B(n_69),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_58),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx6_ASAP7_75t_SL g105 ( 
.A(n_92),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_106),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_93),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_108),
.A2(n_120),
.B(n_109),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_98),
.B1(n_103),
.B2(n_95),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_111),
.A2(n_118),
.B1(n_121),
.B2(n_122),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_113),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_117),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_115),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_50),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_119),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_104),
.A2(n_51),
.B1(n_52),
.B2(n_71),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_98),
.B(n_65),
.Y(n_119)
);

AOI22x1_ASAP7_75t_SL g120 ( 
.A1(n_94),
.A2(n_65),
.B1(n_47),
.B2(n_25),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_94),
.A2(n_18),
.B1(n_40),
.B2(n_39),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_126),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_16),
.C(n_38),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_129),
.A2(n_132),
.B1(n_134),
.B2(n_123),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_130),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_131),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_6),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_22),
.B1(n_34),
.B2(n_33),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_134),
.C(n_125),
.Y(n_141)
);

AOI21x1_ASAP7_75t_L g143 ( 
.A1(n_141),
.A2(n_142),
.B(n_128),
.Y(n_143)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_138),
.B1(n_140),
.B2(n_137),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_127),
.C(n_139),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_133),
.C(n_116),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_137),
.B(n_27),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_147),
.A2(n_17),
.B1(n_28),
.B2(n_45),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_13),
.B(n_32),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_10),
.B(n_30),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_7),
.Y(n_153)
);


endmodule