module real_aes_8096_n_14 (n_13, n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_12, n_1, n_10, n_11, n_14);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_10;
input n_11;
output n_14;
wire n_28;
wire n_17;
wire n_22;
wire n_24;
wire n_41;
wire n_34;
wire n_19;
wire n_40;
wire n_46;
wire n_25;
wire n_47;
wire n_48;
wire n_43;
wire n_32;
wire n_30;
wire n_16;
wire n_37;
wire n_35;
wire n_42;
wire n_39;
wire n_45;
wire n_15;
wire n_27;
wire n_23;
wire n_38;
wire n_29;
wire n_20;
wire n_44;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
NOR2xp33_ASAP7_75t_R g21 ( .A(n_0), .B(n_22), .Y(n_21) );
CKINVDCx20_ASAP7_75t_R g34 ( .A(n_0), .Y(n_34) );
NAND2xp33_ASAP7_75t_SL g40 ( .A(n_0), .B(n_41), .Y(n_40) );
NOR2xp33_ASAP7_75t_R g17 ( .A(n_1), .B(n_18), .Y(n_17) );
NOR2xp33_ASAP7_75t_R g33 ( .A(n_1), .B(n_13), .Y(n_33) );
CKINVDCx20_ASAP7_75t_R g47 ( .A(n_1), .Y(n_47) );
CKINVDCx20_ASAP7_75t_R g27 ( .A(n_2), .Y(n_27) );
NOR3xp33_ASAP7_75t_SL g25 ( .A(n_3), .B(n_9), .C(n_26), .Y(n_25) );
AOI221xp5_ASAP7_75t_SL g14 ( .A1(n_4), .A2(n_6), .B1(n_15), .B2(n_28), .C(n_35), .Y(n_14) );
NOR2xp33_ASAP7_75t_R g19 ( .A(n_5), .B(n_20), .Y(n_19) );
NAND2xp33_ASAP7_75t_SL g29 ( .A(n_5), .B(n_30), .Y(n_29) );
CKINVDCx20_ASAP7_75t_R g43 ( .A(n_5), .Y(n_43) );
CKINVDCx20_ASAP7_75t_R g48 ( .A(n_7), .Y(n_48) );
CKINVDCx5p33_ASAP7_75t_R g26 ( .A(n_8), .Y(n_26) );
INVx1_ASAP7_75t_L g44 ( .A(n_10), .Y(n_44) );
CKINVDCx20_ASAP7_75t_R g23 ( .A(n_11), .Y(n_23) );
NOR4xp25_ASAP7_75t_SL g28 ( .A(n_11), .B(n_29), .C(n_32), .D(n_34), .Y(n_28) );
NOR2xp33_ASAP7_75t_R g37 ( .A(n_11), .B(n_38), .Y(n_37) );
CKINVDCx20_ASAP7_75t_R g22 ( .A(n_12), .Y(n_22) );
NAND4xp25_ASAP7_75t_SL g20 ( .A(n_13), .B(n_21), .C(n_23), .D(n_24), .Y(n_20) );
CKINVDCx20_ASAP7_75t_R g15 ( .A(n_16), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_17), .Y(n_16) );
CKINVDCx16_ASAP7_75t_R g18 ( .A(n_19), .Y(n_18) );
NOR2xp33_ASAP7_75t_R g46 ( .A(n_20), .B(n_43), .Y(n_46) );
NAND2xp33_ASAP7_75t_SL g31 ( .A(n_22), .B(n_24), .Y(n_31) );
AND2x2_ASAP7_75t_L g24 ( .A(n_25), .B(n_27), .Y(n_24) );
NAND2xp33_ASAP7_75t_SL g42 ( .A(n_30), .B(n_43), .Y(n_42) );
CKINVDCx20_ASAP7_75t_R g30 ( .A(n_31), .Y(n_30) );
CKINVDCx20_ASAP7_75t_R g32 ( .A(n_33), .Y(n_32) );
NAND2xp33_ASAP7_75t_SL g38 ( .A(n_33), .B(n_39), .Y(n_38) );
OAI22xp33_ASAP7_75t_SL g35 ( .A1(n_36), .A2(n_44), .B1(n_45), .B2(n_48), .Y(n_35) );
CKINVDCx16_ASAP7_75t_R g36 ( .A(n_37), .Y(n_36) );
CKINVDCx5p33_ASAP7_75t_R g39 ( .A(n_40), .Y(n_39) );
CKINVDCx20_ASAP7_75t_R g41 ( .A(n_42), .Y(n_41) );
NAND2xp33_ASAP7_75t_SL g45 ( .A(n_46), .B(n_47), .Y(n_45) );
endmodule