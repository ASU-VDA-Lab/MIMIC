module fake_jpeg_9984_n_48 (n_3, n_2, n_1, n_0, n_4, n_5, n_48);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_48;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_0),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_0),
.B(n_3),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_16),
.B(n_20),
.Y(n_26)
);

OAI32xp33_ASAP7_75t_L g17 ( 
.A1(n_10),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_17),
.A2(n_22),
.B1(n_23),
.B2(n_10),
.Y(n_24)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_19),
.Y(n_27)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

NAND2x1_ASAP7_75t_SL g20 ( 
.A(n_9),
.B(n_1),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_8),
.A2(n_2),
.B(n_4),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_7),
.B1(n_12),
.B2(n_14),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_13),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_16),
.A2(n_9),
.B1(n_7),
.B2(n_13),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_21),
.C(n_17),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_30),
.A2(n_31),
.B1(n_32),
.B2(n_20),
.Y(n_37)
);

MAJx2_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_20),
.C(n_25),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_35),
.B1(n_36),
.B2(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_37),
.A2(n_27),
.B1(n_23),
.B2(n_29),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_27),
.C(n_28),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_40),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_39),
.B(n_41),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_38),
.B(n_43),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_46),
.B(n_42),
.Y(n_47)
);

AOI211xp5_ASAP7_75t_SL g48 ( 
.A1(n_47),
.A2(n_45),
.B(n_11),
.C(n_18),
.Y(n_48)
);


endmodule