module fake_aes_7812_n_12 (n_3, n_1, n_2, n_0, n_12);
input n_3;
input n_1;
input n_2;
input n_0;
output n_12;
wire n_11;
wire n_6;
wire n_4;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx2_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
OAI22xp5_ASAP7_75t_L g5 ( .A1(n_0), .A2(n_2), .B1(n_1), .B2(n_3), .Y(n_5) );
INVxp67_ASAP7_75t_L g6 ( .A(n_1), .Y(n_6) );
INVx2_ASAP7_75t_L g7 ( .A(n_0), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_4), .B(n_7), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_6), .Y(n_9) );
INVxp67_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
AND2x2_ASAP7_75t_L g11 ( .A(n_10), .B(n_8), .Y(n_11) );
OR3x2_ASAP7_75t_L g12 ( .A(n_11), .B(n_5), .C(n_8), .Y(n_12) );
endmodule