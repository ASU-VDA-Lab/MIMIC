module fake_jpeg_10906_n_240 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_240);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_240;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_0),
.B(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVxp33_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_44),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_18),
.B(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_48),
.B(n_57),
.Y(n_92)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_18),
.B(n_1),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_65),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_10),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_60),
.Y(n_80)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_19),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_64),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_24),
.B(n_1),
.Y(n_65)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_41),
.A2(n_32),
.B1(n_25),
.B2(n_34),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_78),
.A2(n_83),
.B1(n_94),
.B2(n_90),
.Y(n_115)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_59),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_37),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_91),
.C(n_95),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_97),
.Y(n_116)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_36),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_40),
.A2(n_25),
.B1(n_33),
.B2(n_31),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_36),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_64),
.A2(n_30),
.B(n_28),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

INVx2_ASAP7_75t_R g102 ( 
.A(n_70),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_102),
.B(n_111),
.Y(n_137)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_99),
.A2(n_47),
.B1(n_45),
.B2(n_31),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_82),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_108),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_64),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_112),
.Y(n_150)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_72),
.A2(n_26),
.B(n_30),
.C(n_28),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_27),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_124),
.B1(n_128),
.B2(n_66),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_89),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_119),
.Y(n_133)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

INVx4_ASAP7_75t_SL g120 ( 
.A(n_66),
.Y(n_120)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_76),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_123),
.Y(n_134)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_83),
.A2(n_55),
.B1(n_27),
.B2(n_26),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_127),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_2),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_13),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_67),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_68),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_68),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_126),
.A2(n_77),
.B1(n_98),
.B2(n_69),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_141),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_116),
.A2(n_77),
.B1(n_81),
.B2(n_90),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_153),
.B1(n_118),
.B2(n_113),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_109),
.A2(n_92),
.B1(n_100),
.B2(n_74),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_121),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_74),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_147),
.B(n_152),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_120),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_148),
.B(n_154),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_106),
.B(n_100),
.C(n_74),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_118),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_103),
.B(n_14),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_104),
.A2(n_52),
.B1(n_3),
.B2(n_5),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_108),
.B(n_12),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_155),
.B(n_102),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_156),
.B(n_164),
.Y(n_186)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_110),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_160),
.B(n_171),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_143),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_170),
.Y(n_179)
);

AOI21xp33_ASAP7_75t_L g181 ( 
.A1(n_162),
.A2(n_165),
.B(n_167),
.Y(n_181)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_111),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_137),
.A2(n_121),
.B(n_107),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

XOR2x2_ASAP7_75t_SL g193 ( 
.A(n_168),
.B(n_144),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_132),
.A2(n_129),
.B(n_100),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_169),
.A2(n_176),
.B(n_153),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_134),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_101),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_142),
.A2(n_101),
.B1(n_14),
.B2(n_15),
.Y(n_172)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_149),
.Y(n_184)
);

OA22x2_ASAP7_75t_L g176 ( 
.A1(n_132),
.A2(n_13),
.B1(n_131),
.B2(n_141),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_150),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_178),
.C(n_182),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_151),
.C(n_146),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_SL g182 ( 
.A(n_164),
.B(n_155),
.C(n_136),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_183),
.A2(n_165),
.B1(n_159),
.B2(n_176),
.Y(n_198)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_159),
.A2(n_145),
.B1(n_135),
.B2(n_140),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_188),
.A2(n_166),
.B1(n_187),
.B2(n_180),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_156),
.B(n_139),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_161),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_169),
.Y(n_200)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_185),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_195),
.Y(n_210)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_190),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_197),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_198),
.B(n_203),
.Y(n_213)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_188),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_202),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_205),
.Y(n_208)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_189),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_204),
.B(n_175),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_170),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_206),
.A2(n_186),
.B(n_178),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_205),
.Y(n_220)
);

INVx11_ASAP7_75t_L g216 ( 
.A(n_209),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_193),
.C(n_191),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_212),
.C(n_200),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_182),
.C(n_183),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_213),
.A2(n_199),
.B(n_181),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_219),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_206),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_221),
.C(n_211),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_214),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_158),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_212),
.A2(n_192),
.B1(n_197),
.B2(n_194),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_217),
.B1(n_215),
.B2(n_194),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_224),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_216),
.A2(n_210),
.B1(n_196),
.B2(n_176),
.Y(n_225)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_225),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_221),
.A2(n_176),
.B(n_195),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_228),
.Y(n_232)
);

NOR3xp33_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_216),
.C(n_173),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_229),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_231),
.A2(n_222),
.B1(n_220),
.B2(n_226),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_234),
.B(n_235),
.Y(n_236)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_232),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_233),
.A2(n_230),
.B(n_223),
.Y(n_237)
);

O2A1O1Ixp33_ASAP7_75t_L g238 ( 
.A1(n_237),
.A2(n_218),
.B(n_157),
.C(n_163),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_238),
.B(n_236),
.C(n_174),
.Y(n_239)
);

AO21x1_ASAP7_75t_SL g240 ( 
.A1(n_239),
.A2(n_144),
.B(n_135),
.Y(n_240)
);


endmodule