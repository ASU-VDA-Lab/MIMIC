module fake_jpeg_10536_n_114 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_114);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_114;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

BUFx8_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx4f_ASAP7_75t_SL g20 ( 
.A(n_11),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

OR2x2_ASAP7_75t_SL g23 ( 
.A(n_6),
.B(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_29),
.Y(n_40)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_34),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_32),
.B(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_0),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_37),
.B(n_13),
.Y(n_57)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_20),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_48),
.B(n_49),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_42),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_50),
.B(n_57),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_20),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_62),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_21),
.B1(n_16),
.B2(n_34),
.Y(n_52)
);

INVxp67_ASAP7_75t_SL g70 ( 
.A(n_52),
.Y(n_70)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_56),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_21),
.B1(n_30),
.B2(n_17),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_55),
.B1(n_25),
.B2(n_24),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_35),
.A2(n_13),
.B1(n_24),
.B2(n_17),
.Y(n_55)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_59),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_18),
.Y(n_62)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_5),
.C(n_1),
.Y(n_63)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_64),
.Y(n_86)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_45),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_75),
.B(n_76),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_18),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_14),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_77),
.A2(n_53),
.B(n_25),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_74),
.A2(n_50),
.B1(n_60),
.B2(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_82),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_67),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_83),
.B(n_84),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_72),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_76),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_87),
.B(n_69),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_77),
.C(n_69),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_94),
.C(n_78),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_93),
.B(n_95),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_66),
.C(n_70),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_80),
.B(n_22),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_92),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_99),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_81),
.B(n_85),
.Y(n_98)
);

NOR2x1_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_82),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_104),
.Y(n_106)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_103),
.A2(n_102),
.B(n_101),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_105),
.A2(n_0),
.B(n_3),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_106),
.B(n_9),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_107),
.A2(n_108),
.B(n_10),
.Y(n_110)
);

OAI31xp33_ASAP7_75t_L g109 ( 
.A1(n_105),
.A2(n_4),
.A3(n_5),
.B(n_10),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_109),
.B(n_56),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

BUFx24_ASAP7_75t_SL g113 ( 
.A(n_112),
.Y(n_113)
);

NAND2xp33_ASAP7_75t_R g114 ( 
.A(n_113),
.B(n_111),
.Y(n_114)
);


endmodule