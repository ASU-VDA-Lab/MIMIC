module fake_jpeg_29537_n_469 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_469);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_469;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_7),
.B(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g111 ( 
.A(n_47),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_48),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_51),
.Y(n_138)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_14),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_54),
.B(n_59),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_55),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_25),
.B(n_31),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_57),
.B(n_91),
.Y(n_102)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_32),
.B(n_25),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_12),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_60),
.B(n_65),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_64),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_32),
.B(n_11),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_35),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_67),
.B(n_79),
.Y(n_117)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_70),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_15),
.Y(n_78)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_17),
.Y(n_79)
);

INVx11_ASAP7_75t_SL g80 ( 
.A(n_17),
.Y(n_80)
);

CKINVDCx9p33_ASAP7_75t_R g116 ( 
.A(n_80),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_21),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_82),
.Y(n_118)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_37),
.Y(n_82)
);

NAND2x1_ASAP7_75t_L g83 ( 
.A(n_21),
.B(n_1),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_83),
.B(n_2),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_88),
.Y(n_106)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_21),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_90),
.B(n_19),
.Y(n_144)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_93),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_46),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_64),
.A2(n_38),
.B1(n_44),
.B2(n_37),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_94),
.A2(n_110),
.B1(n_125),
.B2(n_129),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_61),
.A2(n_37),
.B1(n_44),
.B2(n_45),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_28),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_60),
.B(n_22),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_140),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_93),
.A2(n_46),
.B1(n_40),
.B2(n_19),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_88),
.A2(n_48),
.B1(n_78),
.B2(n_86),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_49),
.Y(n_131)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_47),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_137),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_47),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_89),
.B(n_26),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_87),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_144),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_51),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_56),
.Y(n_175)
);

OR2x2_ASAP7_75t_SL g147 ( 
.A(n_115),
.B(n_83),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_147),
.B(n_153),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_97),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_150),
.Y(n_206)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_151),
.Y(n_198)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_152),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_154),
.Y(n_210)
);

OR2x2_ASAP7_75t_SL g156 ( 
.A(n_130),
.B(n_44),
.Y(n_156)
);

NOR2x1_ASAP7_75t_L g228 ( 
.A(n_156),
.B(n_173),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_116),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_157),
.B(n_172),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_98),
.Y(n_158)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_158),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_159),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_130),
.A2(n_27),
.B1(n_22),
.B2(n_45),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_167),
.Y(n_194)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_161),
.Y(n_218)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_119),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_164),
.Y(n_214)
);

OR2x4_ASAP7_75t_L g165 ( 
.A(n_102),
.B(n_28),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g211 ( 
.A(n_165),
.B(n_189),
.Y(n_211)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_166),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_117),
.A2(n_21),
.B(n_43),
.Y(n_167)
);

AO22x1_ASAP7_75t_SL g168 ( 
.A1(n_132),
.A2(n_71),
.B1(n_63),
.B2(n_73),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_168),
.A2(n_192),
.B1(n_125),
.B2(n_55),
.Y(n_207)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_170),
.Y(n_225)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_105),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_171),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_109),
.B(n_24),
.Y(n_172)
);

AOI21xp33_ASAP7_75t_L g173 ( 
.A1(n_120),
.A2(n_24),
.B(n_20),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_118),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_174),
.B(n_178),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_175),
.Y(n_199)
);

O2A1O1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_106),
.A2(n_26),
.B(n_16),
.C(n_27),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_176),
.B(n_187),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_111),
.B(n_20),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_177),
.B(n_179),
.Y(n_229)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_114),
.B(n_33),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_136),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_180),
.B(n_181),
.Y(n_226)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_142),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_184),
.Y(n_227)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_131),
.Y(n_184)
);

CKINVDCx12_ASAP7_75t_R g186 ( 
.A(n_111),
.Y(n_186)
);

INVx11_ASAP7_75t_SL g204 ( 
.A(n_186),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_95),
.B(n_33),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_107),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_188),
.Y(n_215)
);

AND2x2_ASAP7_75t_SL g189 ( 
.A(n_121),
.B(n_53),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_107),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_190),
.A2(n_191),
.B1(n_133),
.B2(n_128),
.Y(n_212)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_142),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_94),
.A2(n_85),
.B1(n_84),
.B2(n_75),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_165),
.A2(n_129),
.B1(n_124),
.B2(n_122),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_193),
.A2(n_197),
.B1(n_200),
.B2(n_121),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_182),
.A2(n_122),
.B1(n_124),
.B2(n_103),
.Y(n_195)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_195),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_192),
.A2(n_134),
.B1(n_113),
.B2(n_104),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_156),
.A2(n_176),
.B1(n_168),
.B2(n_185),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_148),
.B(n_16),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_202),
.B(n_217),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_153),
.A2(n_103),
.B1(n_139),
.B2(n_134),
.Y(n_205)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_205),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_207),
.B(n_131),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_147),
.A2(n_139),
.B1(n_146),
.B2(n_95),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_169),
.B(n_42),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_177),
.B(n_146),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_221),
.B(n_189),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_211),
.C(n_194),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_232),
.B(n_246),
.C(n_254),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_233),
.Y(n_281)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_206),
.Y(n_235)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_235),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_236),
.B(n_202),
.Y(n_278)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_206),
.Y(n_237)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_237),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_204),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_238),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_172),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_239),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_228),
.A2(n_42),
.B(n_158),
.Y(n_240)
);

AO21x1_ASAP7_75t_L g285 ( 
.A1(n_240),
.A2(n_256),
.B(n_261),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_242),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_181),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_244),
.Y(n_263)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_210),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_245),
.A2(n_195),
.B1(n_205),
.B2(n_215),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_227),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_246),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_226),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_247),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_222),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_248),
.B(n_249),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_198),
.B(n_141),
.Y(n_249)
);

INVx4_ASAP7_75t_SL g250 ( 
.A(n_224),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_250),
.B(n_252),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_210),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_251),
.A2(n_253),
.B1(n_255),
.B2(n_258),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_213),
.Y(n_252)
);

BUFx4f_ASAP7_75t_SL g253 ( 
.A(n_222),
.Y(n_253)
);

INVx8_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_196),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_257),
.B(n_259),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_213),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_196),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_214),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_260),
.A2(n_218),
.B1(n_222),
.B2(n_215),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_198),
.B(n_171),
.Y(n_261)
);

AOI32xp33_ASAP7_75t_L g262 ( 
.A1(n_231),
.A2(n_199),
.A3(n_229),
.B1(n_228),
.B2(n_194),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_SL g294 ( 
.A(n_262),
.B(n_279),
.C(n_248),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_231),
.A2(n_193),
.B(n_219),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_265),
.A2(n_267),
.B(n_292),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_256),
.A2(n_219),
.B(n_211),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_270),
.A2(n_273),
.B(n_218),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_232),
.B(n_216),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_271),
.B(n_272),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_236),
.B(n_221),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_230),
.A2(n_207),
.B(n_199),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_211),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_275),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_203),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_276),
.A2(n_287),
.B1(n_260),
.B2(n_250),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_278),
.B(n_282),
.Y(n_306)
);

AND2x6_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_209),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_247),
.B(n_241),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_291),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_254),
.A2(n_209),
.B1(n_225),
.B2(n_161),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_234),
.B(n_214),
.C(n_225),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_230),
.A2(n_208),
.B(n_218),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_290),
.B(n_283),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_293),
.B(n_294),
.Y(n_334)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_288),
.Y(n_295)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_295),
.Y(n_332)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_281),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_297),
.Y(n_352)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_281),
.Y(n_298)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_298),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_276),
.A2(n_234),
.B1(n_259),
.B2(n_257),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_300),
.A2(n_307),
.B1(n_317),
.B2(n_277),
.Y(n_325)
);

AND2x6_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_253),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_301),
.B(n_302),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_282),
.B(n_238),
.Y(n_302)
);

OAI31xp33_ASAP7_75t_L g304 ( 
.A1(n_273),
.A2(n_288),
.A3(n_265),
.B(n_285),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_304),
.B(n_99),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_305),
.A2(n_314),
.B(n_315),
.Y(n_324)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_289),
.Y(n_308)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_308),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_280),
.B(n_253),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_309),
.B(n_311),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_244),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_316),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_284),
.B(n_255),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_277),
.B(n_201),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_312),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_264),
.A2(n_237),
.B(n_166),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_285),
.A2(n_149),
.B(n_155),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_289),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_291),
.A2(n_251),
.B1(n_235),
.B2(n_223),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_263),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_318),
.Y(n_346)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_269),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_321),
.Y(n_328)
);

AND2x6_ASAP7_75t_L g320 ( 
.A(n_286),
.B(n_101),
.Y(n_320)
);

A2O1A1Ixp33_ASAP7_75t_L g345 ( 
.A1(n_320),
.A2(n_99),
.B(n_43),
.C(n_21),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_275),
.B(n_233),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_269),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_322),
.B(n_323),
.Y(n_336)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_266),
.Y(n_323)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_325),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_294),
.A2(n_271),
.B1(n_292),
.B2(n_267),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_327),
.A2(n_331),
.B1(n_323),
.B2(n_306),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_300),
.A2(n_274),
.B1(n_272),
.B2(n_266),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_329),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_313),
.B(n_278),
.C(n_268),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_330),
.B(n_337),
.C(n_303),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_295),
.A2(n_268),
.B1(n_150),
.B2(n_159),
.Y(n_331)
);

OA21x2_ASAP7_75t_L g333 ( 
.A1(n_296),
.A2(n_170),
.B(n_163),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_333),
.B(n_351),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_299),
.B(n_99),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_335),
.B(n_303),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_313),
.B(n_184),
.C(n_155),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_310),
.B(n_316),
.Y(n_338)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_338),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_296),
.A2(n_154),
.B1(n_101),
.B2(n_127),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_339),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_304),
.A2(n_108),
.B1(n_149),
.B2(n_5),
.Y(n_341)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_341),
.Y(n_366)
);

CKINVDCx14_ASAP7_75t_R g372 ( 
.A(n_342),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_305),
.A2(n_3),
.B(n_4),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_344),
.A2(n_345),
.B(n_350),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_314),
.A2(n_3),
.B(n_5),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_315),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_352),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_353),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_330),
.B(n_299),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_355),
.B(n_356),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_337),
.B(n_306),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_334),
.A2(n_321),
.B(n_320),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_357),
.B(n_333),
.Y(n_397)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_352),
.Y(n_358)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_358),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_360),
.A2(n_371),
.B1(n_341),
.B2(n_339),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_361),
.B(n_363),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_335),
.B(n_301),
.C(n_298),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_376),
.C(n_324),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_329),
.B(n_297),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_365),
.B(n_368),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_327),
.B(n_43),
.Y(n_368)
);

MAJx2_ASAP7_75t_L g369 ( 
.A(n_340),
.B(n_43),
.C(n_21),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_369),
.B(n_370),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_328),
.B(n_43),
.Y(n_370)
);

OAI22x1_ASAP7_75t_L g371 ( 
.A1(n_333),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_371)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_336),
.Y(n_374)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_374),
.Y(n_380)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_336),
.Y(n_375)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_375),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_328),
.B(n_43),
.C(n_19),
.Y(n_376)
);

NAND3xp33_ASAP7_75t_L g379 ( 
.A(n_372),
.B(n_346),
.C(n_349),
.Y(n_379)
);

CKINVDCx14_ASAP7_75t_R g410 ( 
.A(n_379),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_359),
.A2(n_342),
.B(n_324),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_382),
.A2(n_397),
.B(n_367),
.Y(n_413)
);

BUFx24_ASAP7_75t_SL g383 ( 
.A(n_369),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_383),
.B(n_387),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_385),
.B(n_366),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_362),
.Y(n_386)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_386),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_364),
.B(n_346),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_376),
.B(n_343),
.Y(n_389)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_389),
.Y(n_405)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_370),
.Y(n_390)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_390),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_391),
.B(n_394),
.Y(n_415)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_358),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_392),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_377),
.A2(n_351),
.B1(n_325),
.B2(n_332),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_393),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_361),
.B(n_338),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_395),
.B(n_326),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_378),
.B(n_363),
.C(n_373),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_406),
.C(n_408),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_404),
.A2(n_377),
.B1(n_385),
.B2(n_371),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_378),
.B(n_391),
.C(n_395),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_381),
.B(n_373),
.C(n_354),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_393),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_409),
.B(n_386),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_411),
.B(n_415),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_397),
.B(n_394),
.C(n_388),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_412),
.B(n_344),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_413),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_382),
.A2(n_348),
.B(n_326),
.Y(n_414)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_414),
.Y(n_428)
);

INVx11_ASAP7_75t_L g416 ( 
.A(n_402),
.Y(n_416)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_416),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_403),
.A2(n_384),
.B(n_380),
.Y(n_417)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_417),
.Y(n_436)
);

OR2x2_ASAP7_75t_L g441 ( 
.A(n_418),
.B(n_420),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_419),
.Y(n_438)
);

INVx11_ASAP7_75t_L g420 ( 
.A(n_402),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_403),
.A2(n_332),
.B1(n_348),
.B2(n_345),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_421),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_422),
.A2(n_429),
.B(n_415),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_404),
.A2(n_401),
.B1(n_407),
.B2(n_410),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_424),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_408),
.A2(n_398),
.B1(n_350),
.B2(n_347),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_425),
.B(n_8),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_412),
.A2(n_398),
.B(n_347),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_405),
.B(n_353),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_430),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_399),
.B(n_396),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_431),
.B(n_427),
.Y(n_444)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_433),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_426),
.B(n_406),
.C(n_400),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_435),
.B(n_437),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_426),
.B(n_331),
.C(n_35),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_427),
.B(n_35),
.C(n_19),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_439),
.B(n_440),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_442),
.B(n_425),
.Y(n_449)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_444),
.Y(n_452)
);

OAI21xp33_ASAP7_75t_L g445 ( 
.A1(n_436),
.A2(n_423),
.B(n_428),
.Y(n_445)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_445),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_435),
.A2(n_429),
.B(n_424),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_447),
.B(n_448),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_438),
.A2(n_417),
.B(n_418),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_449),
.B(n_453),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_434),
.A2(n_438),
.B1(n_443),
.B2(n_442),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_452),
.B(n_443),
.C(n_441),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_454),
.B(n_456),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_450),
.B(n_446),
.C(n_449),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_451),
.B(n_441),
.C(n_421),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_458),
.B(n_419),
.Y(n_462)
);

AO21x1_ASAP7_75t_L g461 ( 
.A1(n_457),
.A2(n_445),
.B(n_432),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_461),
.A2(n_462),
.B(n_455),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_463),
.B(n_464),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_460),
.A2(n_459),
.B(n_416),
.Y(n_464)
);

A2O1A1Ixp33_ASAP7_75t_L g466 ( 
.A1(n_465),
.A2(n_420),
.B(n_9),
.C(n_10),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_466),
.A2(n_8),
.B(n_9),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_467),
.B(n_10),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_468),
.A2(n_35),
.B(n_293),
.Y(n_469)
);


endmodule