module fake_aes_12586_n_679 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_679);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_679;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_50), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_63), .Y(n_87) );
BUFx3_ASAP7_75t_L g88 ( .A(n_80), .Y(n_88) );
CKINVDCx20_ASAP7_75t_R g89 ( .A(n_42), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_29), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_60), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_20), .Y(n_92) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_75), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_31), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_85), .Y(n_95) );
CKINVDCx20_ASAP7_75t_R g96 ( .A(n_61), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_53), .Y(n_97) );
INVxp67_ASAP7_75t_L g98 ( .A(n_33), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_24), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_83), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_30), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_45), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_68), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_77), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_81), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_74), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_25), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_16), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_1), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_12), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_22), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_7), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_19), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_3), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_17), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_39), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_51), .Y(n_117) );
BUFx3_ASAP7_75t_L g118 ( .A(n_14), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_84), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_26), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_7), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_32), .Y(n_122) );
BUFx5_ASAP7_75t_L g123 ( .A(n_38), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_58), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_4), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_23), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_73), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_72), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_10), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_121), .Y(n_130) );
INVx4_ASAP7_75t_L g131 ( .A(n_88), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g132 ( .A(n_123), .B(n_0), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_123), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_123), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_123), .Y(n_135) );
AND2x2_ASAP7_75t_SL g136 ( .A(n_106), .B(n_82), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_114), .B(n_0), .Y(n_137) );
INVx6_ASAP7_75t_L g138 ( .A(n_123), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_121), .Y(n_139) );
BUFx2_ASAP7_75t_L g140 ( .A(n_114), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_123), .Y(n_141) );
AND2x2_ASAP7_75t_L g142 ( .A(n_118), .B(n_1), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_118), .B(n_2), .Y(n_143) );
AND2x2_ASAP7_75t_SL g144 ( .A(n_91), .B(n_21), .Y(n_144) );
AND2x4_ASAP7_75t_L g145 ( .A(n_88), .B(n_2), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_110), .B(n_3), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_123), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_91), .Y(n_148) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_92), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_138), .Y(n_150) );
OR2x2_ASAP7_75t_L g151 ( .A(n_140), .B(n_108), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_133), .Y(n_152) );
BUFx2_ASAP7_75t_L g153 ( .A(n_149), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_133), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_136), .B(n_124), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_140), .B(n_98), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_143), .Y(n_157) );
INVx4_ASAP7_75t_L g158 ( .A(n_145), .Y(n_158) );
NAND3xp33_ASAP7_75t_L g159 ( .A(n_142), .B(n_113), .C(n_112), .Y(n_159) );
INVx1_ASAP7_75t_SL g160 ( .A(n_136), .Y(n_160) );
INVx4_ASAP7_75t_SL g161 ( .A(n_138), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_134), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_131), .B(n_124), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_134), .Y(n_164) );
AND3x2_ASAP7_75t_L g165 ( .A(n_143), .B(n_129), .C(n_115), .Y(n_165) );
OR2x6_ASAP7_75t_L g166 ( .A(n_143), .B(n_125), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_131), .B(n_86), .Y(n_167) );
AND2x4_ASAP7_75t_SL g168 ( .A(n_137), .B(n_89), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_135), .Y(n_169) );
INVx5_ASAP7_75t_L g170 ( .A(n_138), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_135), .Y(n_171) );
INVx4_ASAP7_75t_L g172 ( .A(n_145), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_141), .Y(n_173) );
XNOR2xp5_ASAP7_75t_L g174 ( .A(n_136), .B(n_109), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_137), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_141), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_147), .Y(n_177) );
AOI22xp33_ASAP7_75t_L g178 ( .A1(n_144), .A2(n_128), .B1(n_127), .B2(n_95), .Y(n_178) );
AOI22xp33_ASAP7_75t_L g179 ( .A1(n_178), .A2(n_144), .B1(n_137), .B2(n_145), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_175), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_156), .B(n_146), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_158), .B(n_172), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_158), .B(n_142), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_158), .B(n_145), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_172), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_172), .B(n_144), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_153), .B(n_137), .Y(n_187) );
AO22x1_ASAP7_75t_L g188 ( .A1(n_160), .A2(n_107), .B1(n_99), .B2(n_103), .Y(n_188) );
NAND2x1p5_ASAP7_75t_L g189 ( .A(n_157), .B(n_132), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_151), .B(n_131), .Y(n_190) );
NOR2x2_ASAP7_75t_L g191 ( .A(n_174), .B(n_109), .Y(n_191) );
NAND2x1_ASAP7_75t_L g192 ( .A(n_166), .B(n_138), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_150), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_152), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_152), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_150), .Y(n_196) );
NOR2xp33_ASAP7_75t_SL g197 ( .A(n_168), .B(n_89), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_155), .A2(n_96), .B1(n_116), .B2(n_120), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_166), .A2(n_147), .B1(n_148), .B2(n_139), .Y(n_199) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_166), .A2(n_148), .B1(n_139), .B2(n_130), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_166), .A2(n_96), .B1(n_120), .B2(n_116), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_159), .B(n_87), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_163), .B(n_130), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_154), .Y(n_204) );
NOR2xp33_ASAP7_75t_SL g205 ( .A(n_153), .B(n_90), .Y(n_205) );
INVxp67_ASAP7_75t_L g206 ( .A(n_151), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_154), .Y(n_207) );
INVx3_ASAP7_75t_L g208 ( .A(n_164), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_164), .Y(n_209) );
INVxp67_ASAP7_75t_SL g210 ( .A(n_168), .Y(n_210) );
NOR3xp33_ASAP7_75t_L g211 ( .A(n_167), .B(n_119), .C(n_111), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_169), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_174), .A2(n_105), .B1(n_122), .B2(n_117), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_165), .B(n_94), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_162), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_162), .Y(n_216) );
BUFx3_ASAP7_75t_L g217 ( .A(n_150), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_181), .A2(n_173), .B(n_176), .C(n_177), .Y(n_218) );
OAI21xp5_ASAP7_75t_L g219 ( .A1(n_186), .A2(n_173), .B(n_176), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_206), .B(n_150), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_187), .B(n_169), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_185), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_215), .Y(n_223) );
OAI22xp5_ASAP7_75t_L g224 ( .A1(n_179), .A2(n_171), .B1(n_97), .B2(n_100), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_215), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_187), .A2(n_101), .B(n_102), .C(n_104), .Y(n_226) );
AO32x1_ASAP7_75t_L g227 ( .A1(n_216), .A2(n_101), .A3(n_102), .B1(n_93), .B2(n_8), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_190), .B(n_161), .Y(n_228) );
BUFx2_ASAP7_75t_L g229 ( .A(n_210), .Y(n_229) );
BUFx8_ASAP7_75t_L g230 ( .A(n_197), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_216), .Y(n_231) );
INVxp67_ASAP7_75t_SL g232 ( .A(n_201), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_201), .B(n_4), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_211), .B(n_161), .Y(n_234) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_185), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_180), .A2(n_93), .B(n_126), .C(n_150), .Y(n_236) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_185), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_183), .B(n_161), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_205), .B(n_170), .Y(n_239) );
INVxp67_ASAP7_75t_L g240 ( .A(n_197), .Y(n_240) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_200), .A2(n_93), .B1(n_170), .B2(n_8), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_185), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_213), .B(n_170), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_199), .B(n_170), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_185), .B(n_182), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_188), .B(n_170), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_SL g247 ( .A1(n_208), .A2(n_93), .B(n_48), .C(n_49), .Y(n_247) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_192), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g249 ( .A1(n_213), .A2(n_5), .B1(n_6), .B2(n_9), .Y(n_249) );
INVx4_ASAP7_75t_L g250 ( .A(n_208), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_223), .Y(n_251) );
AOI211x1_ASAP7_75t_L g252 ( .A1(n_241), .A2(n_188), .B(n_202), .C(n_203), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_238), .A2(n_184), .B(n_192), .Y(n_253) );
OAI21x1_ASAP7_75t_L g254 ( .A1(n_219), .A2(n_189), .B(n_208), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_221), .B(n_198), .Y(n_255) );
INVx3_ASAP7_75t_L g256 ( .A(n_222), .Y(n_256) );
AO21x2_ASAP7_75t_L g257 ( .A1(n_247), .A2(n_204), .B(n_194), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_232), .B(n_198), .Y(n_258) );
OAI22xp5_ASAP7_75t_L g259 ( .A1(n_225), .A2(n_204), .B1(n_194), .B2(n_212), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_231), .Y(n_260) );
OAI21x1_ASAP7_75t_L g261 ( .A1(n_219), .A2(n_189), .B(n_209), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_218), .Y(n_262) );
A2O1A1Ixp33_ASAP7_75t_L g263 ( .A1(n_226), .A2(n_209), .B(n_207), .C(n_195), .Y(n_263) );
AO221x1_ASAP7_75t_L g264 ( .A1(n_240), .A2(n_191), .B1(n_193), .B2(n_196), .C(n_195), .Y(n_264) );
INVx5_ASAP7_75t_L g265 ( .A(n_222), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_222), .Y(n_266) );
NOR2xp33_ASAP7_75t_R g267 ( .A(n_230), .B(n_214), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g268 ( .A1(n_243), .A2(n_217), .B(n_196), .C(n_193), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_235), .Y(n_269) );
AND2x4_ASAP7_75t_L g270 ( .A(n_248), .B(n_217), .Y(n_270) );
OAI21x1_ASAP7_75t_L g271 ( .A1(n_246), .A2(n_189), .B(n_196), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_248), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_245), .A2(n_196), .B(n_193), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_228), .A2(n_196), .B(n_193), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_251), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_251), .B(n_233), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_260), .Y(n_277) );
OAI21x1_ASAP7_75t_SL g278 ( .A1(n_262), .A2(n_241), .B(n_249), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_259), .Y(n_279) );
OAI21xp33_ASAP7_75t_SL g280 ( .A1(n_264), .A2(n_239), .B(n_250), .Y(n_280) );
OAI21x1_ASAP7_75t_L g281 ( .A1(n_271), .A2(n_242), .B(n_234), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_261), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_272), .Y(n_283) );
AO31x2_ASAP7_75t_L g284 ( .A1(n_262), .A2(n_236), .A3(n_227), .B(n_220), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_272), .Y(n_285) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_265), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_274), .A2(n_227), .B(n_244), .Y(n_287) );
OAI21x1_ASAP7_75t_L g288 ( .A1(n_271), .A2(n_227), .B(n_224), .Y(n_288) );
A2O1A1Ixp33_ASAP7_75t_L g289 ( .A1(n_253), .A2(n_248), .B(n_229), .C(n_237), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_265), .B(n_250), .Y(n_290) );
BUFx12f_ASAP7_75t_L g291 ( .A(n_265), .Y(n_291) );
AOI221xp5_ASAP7_75t_L g292 ( .A1(n_258), .A2(n_235), .B1(n_237), .B2(n_230), .C(n_193), .Y(n_292) );
OR2x6_ASAP7_75t_L g293 ( .A(n_252), .B(n_237), .Y(n_293) );
AO21x2_ASAP7_75t_L g294 ( .A1(n_268), .A2(n_235), .B(n_6), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_255), .B(n_5), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_275), .Y(n_296) );
AO21x2_ASAP7_75t_L g297 ( .A1(n_287), .A2(n_254), .B(n_261), .Y(n_297) );
OR2x2_ASAP7_75t_L g298 ( .A(n_275), .B(n_270), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_275), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_282), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_282), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_291), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_282), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_279), .Y(n_304) );
AO21x2_ASAP7_75t_L g305 ( .A1(n_278), .A2(n_254), .B(n_257), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_279), .Y(n_306) );
NOR2x1_ASAP7_75t_R g307 ( .A(n_291), .B(n_264), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_281), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_277), .B(n_266), .Y(n_309) );
OAI21xp5_ASAP7_75t_L g310 ( .A1(n_295), .A2(n_263), .B(n_273), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_285), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_280), .Y(n_312) );
OA21x2_ASAP7_75t_L g313 ( .A1(n_288), .A2(n_269), .B(n_266), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_281), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_285), .Y(n_315) );
BUFx3_ASAP7_75t_L g316 ( .A(n_291), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_293), .B(n_265), .Y(n_317) );
OA21x2_ASAP7_75t_L g318 ( .A1(n_288), .A2(n_269), .B(n_270), .Y(n_318) );
BUFx3_ASAP7_75t_L g319 ( .A(n_290), .Y(n_319) );
AND2x4_ASAP7_75t_L g320 ( .A(n_293), .B(n_265), .Y(n_320) );
NOR2x1_ASAP7_75t_R g321 ( .A(n_290), .B(n_256), .Y(n_321) );
INVx3_ASAP7_75t_L g322 ( .A(n_290), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_283), .Y(n_323) );
INVx3_ASAP7_75t_L g324 ( .A(n_290), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_296), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_296), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_304), .B(n_293), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_300), .Y(n_328) );
BUFx2_ASAP7_75t_L g329 ( .A(n_307), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_296), .Y(n_330) );
NOR2xp67_ASAP7_75t_L g331 ( .A(n_299), .B(n_280), .Y(n_331) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_323), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_304), .B(n_293), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_299), .Y(n_334) );
BUFx3_ASAP7_75t_L g335 ( .A(n_302), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_304), .B(n_293), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_299), .B(n_277), .Y(n_337) );
BUFx2_ASAP7_75t_L g338 ( .A(n_307), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_306), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_306), .Y(n_340) );
OAI211xp5_ASAP7_75t_L g341 ( .A1(n_302), .A2(n_276), .B(n_267), .C(n_292), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_311), .B(n_276), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_306), .B(n_294), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_302), .B(n_295), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_300), .B(n_294), .Y(n_345) );
INVx3_ASAP7_75t_L g346 ( .A(n_317), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_300), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_300), .Y(n_348) );
INVx2_ASAP7_75t_SL g349 ( .A(n_319), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_301), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_323), .A2(n_278), .B1(n_294), .B2(n_286), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_301), .B(n_294), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_311), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_301), .B(n_284), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_311), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_302), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_315), .B(n_284), .Y(n_357) );
INVx1_ASAP7_75t_SL g358 ( .A(n_319), .Y(n_358) );
INVxp67_ASAP7_75t_SL g359 ( .A(n_301), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_315), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_303), .B(n_284), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_303), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_315), .Y(n_363) );
INVxp67_ASAP7_75t_L g364 ( .A(n_307), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_316), .B(n_322), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_303), .Y(n_366) );
INVxp67_ASAP7_75t_SL g367 ( .A(n_303), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_309), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_309), .Y(n_369) );
INVx4_ASAP7_75t_L g370 ( .A(n_316), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_308), .Y(n_371) );
BUFx2_ASAP7_75t_L g372 ( .A(n_319), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_339), .Y(n_373) );
INVx1_ASAP7_75t_SL g374 ( .A(n_356), .Y(n_374) );
NAND2x1_ASAP7_75t_L g375 ( .A(n_370), .B(n_312), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_371), .Y(n_376) );
AOI221xp5_ASAP7_75t_L g377 ( .A1(n_332), .A2(n_312), .B1(n_310), .B2(n_316), .C(n_298), .Y(n_377) );
AND2x4_ASAP7_75t_L g378 ( .A(n_346), .B(n_312), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_339), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_340), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_327), .B(n_318), .Y(n_381) );
INVx1_ASAP7_75t_SL g382 ( .A(n_335), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_340), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_353), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_353), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_355), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g387 ( .A1(n_341), .A2(n_316), .B1(n_322), .B2(n_324), .Y(n_387) );
NAND4xp25_ASAP7_75t_L g388 ( .A(n_351), .B(n_310), .C(n_298), .D(n_289), .Y(n_388) );
INVxp67_ASAP7_75t_SL g389 ( .A(n_359), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_327), .B(n_318), .Y(n_390) );
BUFx2_ASAP7_75t_L g391 ( .A(n_370), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_329), .A2(n_319), .B1(n_322), .B2(n_324), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_333), .B(n_318), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_333), .B(n_318), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_333), .B(n_318), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_371), .Y(n_396) );
NAND2x1p5_ASAP7_75t_L g397 ( .A(n_370), .B(n_335), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_355), .Y(n_398) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_335), .Y(n_399) );
INVx1_ASAP7_75t_SL g400 ( .A(n_370), .Y(n_400) );
NAND2x1_ASAP7_75t_SL g401 ( .A(n_331), .B(n_317), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_328), .Y(n_402) );
AND2x4_ASAP7_75t_L g403 ( .A(n_346), .B(n_305), .Y(n_403) );
INVx4_ASAP7_75t_L g404 ( .A(n_329), .Y(n_404) );
CKINVDCx14_ASAP7_75t_R g405 ( .A(n_338), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_371), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_337), .B(n_298), .Y(n_407) );
INVx3_ASAP7_75t_L g408 ( .A(n_328), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_336), .B(n_305), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_372), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_336), .B(n_305), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_360), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_337), .B(n_322), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_343), .B(n_305), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_343), .B(n_305), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_360), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_328), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_347), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_363), .Y(n_419) );
INVx5_ASAP7_75t_L g420 ( .A(n_338), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_347), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_343), .B(n_305), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_357), .B(n_297), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_354), .B(n_297), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_357), .B(n_297), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_347), .Y(n_426) );
INVx2_ASAP7_75t_SL g427 ( .A(n_372), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_354), .B(n_297), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_354), .B(n_297), .Y(n_429) );
NAND2xp5_ASAP7_75t_SL g430 ( .A(n_364), .B(n_317), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_363), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_348), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_325), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_342), .B(n_324), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_361), .B(n_297), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_361), .B(n_308), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_361), .B(n_308), .Y(n_437) );
INVx3_ASAP7_75t_L g438 ( .A(n_348), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_346), .B(n_308), .Y(n_439) );
INVx1_ASAP7_75t_SL g440 ( .A(n_358), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_373), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_391), .B(n_349), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_373), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_424), .B(n_325), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_391), .B(n_349), .Y(n_445) );
INVx1_ASAP7_75t_SL g446 ( .A(n_400), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_379), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_413), .B(n_326), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_379), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_380), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_399), .B(n_349), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_409), .B(n_346), .Y(n_452) );
AND3x2_ASAP7_75t_L g453 ( .A(n_405), .B(n_364), .C(n_365), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_409), .B(n_358), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_407), .B(n_326), .Y(n_455) );
AND2x4_ASAP7_75t_L g456 ( .A(n_378), .B(n_345), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_408), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_433), .B(n_368), .Y(n_458) );
INVx1_ASAP7_75t_SL g459 ( .A(n_382), .Y(n_459) );
INVx2_ASAP7_75t_SL g460 ( .A(n_374), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_411), .B(n_330), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_424), .B(n_330), .Y(n_462) );
NOR2x1_ASAP7_75t_SL g463 ( .A(n_404), .B(n_341), .Y(n_463) );
NAND2x1p5_ASAP7_75t_L g464 ( .A(n_375), .B(n_322), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_383), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_428), .B(n_334), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_384), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_381), .B(n_368), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_434), .B(n_367), .Y(n_469) );
OAI21xp33_ASAP7_75t_L g470 ( .A1(n_377), .A2(n_344), .B(n_342), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_387), .A2(n_331), .B1(n_369), .B2(n_322), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_384), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_428), .B(n_369), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_381), .B(n_345), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_429), .B(n_345), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_408), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_385), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_429), .B(n_352), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_436), .B(n_367), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_387), .A2(n_324), .B1(n_366), .B2(n_320), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_408), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_385), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_435), .B(n_352), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_386), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_390), .B(n_352), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_386), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_436), .B(n_366), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_398), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_398), .Y(n_489) );
INVx3_ASAP7_75t_L g490 ( .A(n_375), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_437), .B(n_348), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_433), .B(n_350), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_412), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_390), .B(n_324), .Y(n_494) );
AND2x4_ASAP7_75t_L g495 ( .A(n_378), .B(n_317), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_412), .Y(n_496) );
OR2x2_ASAP7_75t_SL g497 ( .A(n_410), .B(n_350), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_435), .B(n_350), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_416), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_437), .B(n_362), .Y(n_500) );
AND2x4_ASAP7_75t_L g501 ( .A(n_378), .B(n_317), .Y(n_501) );
AND2x2_ASAP7_75t_SL g502 ( .A(n_404), .B(n_317), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_408), .Y(n_503) );
AND2x2_ASAP7_75t_SL g504 ( .A(n_404), .B(n_320), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_416), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_414), .B(n_362), .Y(n_506) );
NOR2xp67_ASAP7_75t_SL g507 ( .A(n_420), .B(n_321), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_393), .B(n_320), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_414), .B(n_415), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_438), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_419), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_427), .B(n_314), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_427), .B(n_314), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_415), .B(n_314), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_438), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_419), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_388), .A2(n_320), .B1(n_313), .B2(n_314), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_394), .B(n_313), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_431), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_452), .B(n_395), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_461), .B(n_422), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_441), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_443), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_447), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_460), .B(n_430), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_449), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_508), .B(n_395), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_479), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_468), .B(n_423), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_450), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_509), .B(n_425), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_444), .B(n_425), .Y(n_532) );
NAND4xp25_ASAP7_75t_L g533 ( .A(n_517), .B(n_392), .C(n_403), .D(n_440), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_444), .B(n_431), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_475), .B(n_389), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_475), .B(n_438), .Y(n_536) );
OAI21xp33_ASAP7_75t_SL g537 ( .A1(n_502), .A2(n_401), .B(n_397), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_446), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_465), .Y(n_539) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_459), .Y(n_540) );
INVxp67_ASAP7_75t_L g541 ( .A(n_446), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_467), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_462), .B(n_418), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_478), .B(n_378), .Y(n_544) );
AOI211xp5_ASAP7_75t_L g545 ( .A1(n_470), .A2(n_321), .B(n_403), .C(n_439), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_466), .B(n_439), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_512), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_472), .Y(n_548) );
AND2x2_ASAP7_75t_SL g549 ( .A(n_504), .B(n_403), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_477), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_482), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_474), .B(n_420), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_484), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_485), .B(n_420), .Y(n_554) );
OR2x6_ASAP7_75t_L g555 ( .A(n_464), .B(n_401), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_454), .B(n_420), .Y(n_556) );
INVx1_ASAP7_75t_SL g557 ( .A(n_442), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_473), .B(n_418), .Y(n_558) );
INVxp67_ASAP7_75t_L g559 ( .A(n_451), .Y(n_559) );
O2A1O1Ixp5_ASAP7_75t_R g560 ( .A1(n_473), .A2(n_420), .B(n_11), .C(n_12), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_494), .B(n_420), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_483), .B(n_418), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_483), .B(n_426), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_486), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_498), .B(n_432), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_488), .Y(n_566) );
AND2x4_ASAP7_75t_L g567 ( .A(n_495), .B(n_432), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_489), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_493), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_496), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_456), .B(n_432), .Y(n_571) );
AOI31xp33_ASAP7_75t_L g572 ( .A1(n_464), .A2(n_321), .A3(n_417), .B(n_421), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_498), .B(n_402), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_499), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_505), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_511), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_518), .B(n_417), .Y(n_577) );
NOR2xp67_ASAP7_75t_SL g578 ( .A(n_490), .B(n_256), .Y(n_578) );
INVxp67_ASAP7_75t_L g579 ( .A(n_445), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_455), .B(n_10), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_487), .B(n_421), .Y(n_581) );
INVx1_ASAP7_75t_SL g582 ( .A(n_497), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_456), .B(n_495), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_516), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_532), .B(n_506), .Y(n_585) );
AOI31xp33_ASAP7_75t_L g586 ( .A1(n_537), .A2(n_453), .A3(n_463), .B(n_480), .Y(n_586) );
INVxp67_ASAP7_75t_L g587 ( .A(n_540), .Y(n_587) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_572), .A2(n_480), .B(n_490), .Y(n_588) );
INVxp67_ASAP7_75t_SL g589 ( .A(n_541), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_522), .Y(n_590) );
INVx1_ASAP7_75t_SL g591 ( .A(n_557), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_531), .B(n_514), .Y(n_592) );
OAI32xp33_ASAP7_75t_L g593 ( .A1(n_582), .A2(n_491), .A3(n_500), .B1(n_469), .B2(n_448), .Y(n_593) );
OAI221xp5_ASAP7_75t_L g594 ( .A1(n_537), .A2(n_517), .B1(n_471), .B2(n_507), .C(n_458), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_583), .B(n_501), .Y(n_595) );
OAI21xp33_ASAP7_75t_SL g596 ( .A1(n_582), .A2(n_471), .B(n_514), .Y(n_596) );
O2A1O1Ixp33_ASAP7_75t_L g597 ( .A1(n_560), .A2(n_519), .B(n_515), .C(n_476), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_559), .B(n_501), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_580), .A2(n_510), .B1(n_503), .B2(n_481), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_549), .A2(n_513), .B1(n_492), .B2(n_457), .Y(n_600) );
INVxp67_ASAP7_75t_L g601 ( .A(n_525), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_581), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_533), .A2(n_406), .B1(n_396), .B2(n_376), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_579), .B(n_11), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_527), .B(n_406), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_523), .Y(n_606) );
AOI21xp33_ASAP7_75t_L g607 ( .A1(n_545), .A2(n_13), .B(n_15), .Y(n_607) );
AOI322xp5_ASAP7_75t_L g608 ( .A1(n_521), .A2(n_396), .A3(n_376), .B1(n_20), .B2(n_19), .C1(n_18), .C2(n_270), .Y(n_608) );
INVxp67_ASAP7_75t_SL g609 ( .A(n_538), .Y(n_609) );
O2A1O1Ixp33_ASAP7_75t_L g610 ( .A1(n_572), .A2(n_396), .B(n_18), .C(n_256), .Y(n_610) );
OAI21xp33_ASAP7_75t_L g611 ( .A1(n_533), .A2(n_284), .B(n_27), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_524), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_534), .B(n_313), .Y(n_613) );
INVx2_ASAP7_75t_SL g614 ( .A(n_557), .Y(n_614) );
O2A1O1Ixp33_ASAP7_75t_L g615 ( .A1(n_555), .A2(n_257), .B(n_284), .C(n_28), .Y(n_615) );
INVx1_ASAP7_75t_SL g616 ( .A(n_535), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_526), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_530), .Y(n_618) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_547), .Y(n_619) );
OAI222xp33_ASAP7_75t_L g620 ( .A1(n_594), .A2(n_555), .B1(n_544), .B2(n_552), .C1(n_554), .C2(n_536), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_616), .B(n_529), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_601), .A2(n_567), .B1(n_528), .B2(n_571), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_590), .Y(n_623) );
INVx2_ASAP7_75t_SL g624 ( .A(n_614), .Y(n_624) );
OAI22xp33_ASAP7_75t_L g625 ( .A1(n_586), .A2(n_555), .B1(n_546), .B2(n_563), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g626 ( .A1(n_610), .A2(n_543), .B(n_573), .Y(n_626) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_593), .A2(n_584), .B1(n_539), .B2(n_542), .C(n_576), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_594), .A2(n_567), .B1(n_562), .B2(n_577), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_588), .A2(n_520), .B1(n_565), .B2(n_561), .Y(n_629) );
OAI21xp5_ASAP7_75t_L g630 ( .A1(n_610), .A2(n_578), .B(n_573), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_606), .Y(n_631) );
AOI21xp33_ASAP7_75t_L g632 ( .A1(n_597), .A2(n_575), .B(n_574), .Y(n_632) );
OAI321xp33_ASAP7_75t_L g633 ( .A1(n_603), .A2(n_556), .A3(n_558), .B1(n_568), .B2(n_566), .C(n_564), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g634 ( .A1(n_588), .A2(n_570), .B(n_569), .Y(n_634) );
OAI21xp5_ASAP7_75t_SL g635 ( .A1(n_607), .A2(n_553), .B(n_551), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_612), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_617), .Y(n_637) );
AOI21xp33_ASAP7_75t_L g638 ( .A1(n_597), .A2(n_550), .B(n_548), .Y(n_638) );
INVxp33_ASAP7_75t_L g639 ( .A(n_604), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_591), .B(n_34), .Y(n_640) );
OAI222xp33_ASAP7_75t_L g641 ( .A1(n_600), .A2(n_35), .B1(n_36), .B2(n_37), .C1(n_40), .C2(n_41), .Y(n_641) );
OAI321xp33_ASAP7_75t_L g642 ( .A1(n_611), .A2(n_43), .A3(n_44), .B1(n_46), .B2(n_47), .C(n_52), .Y(n_642) );
OA21x2_ASAP7_75t_SL g643 ( .A1(n_596), .A2(n_54), .B(n_55), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_587), .B(n_56), .Y(n_644) );
AOI22xp5_ASAP7_75t_SL g645 ( .A1(n_589), .A2(n_57), .B1(n_59), .B2(n_62), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_585), .B(n_64), .Y(n_646) );
AO22x2_ASAP7_75t_L g647 ( .A1(n_609), .A2(n_65), .B1(n_66), .B2(n_67), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_618), .Y(n_648) );
OAI221xp5_ASAP7_75t_L g649 ( .A1(n_599), .A2(n_69), .B1(n_70), .B2(n_71), .C(n_76), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_598), .B(n_78), .Y(n_650) );
NOR2xp67_ASAP7_75t_L g651 ( .A(n_619), .B(n_79), .Y(n_651) );
OAI21xp33_ASAP7_75t_L g652 ( .A1(n_608), .A2(n_613), .B(n_592), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_595), .B(n_602), .Y(n_653) );
AOI322xp5_ASAP7_75t_L g654 ( .A1(n_605), .A2(n_596), .A3(n_582), .B1(n_603), .B2(n_560), .C1(n_604), .C2(n_616), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_615), .A2(n_586), .B(n_610), .Y(n_655) );
NOR4xp25_ASAP7_75t_L g656 ( .A(n_638), .B(n_632), .C(n_620), .D(n_625), .Y(n_656) );
NOR3xp33_ASAP7_75t_SL g657 ( .A(n_655), .B(n_635), .C(n_634), .Y(n_657) );
OAI221xp5_ASAP7_75t_L g658 ( .A1(n_654), .A2(n_628), .B1(n_634), .B2(n_627), .C(n_652), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_639), .B(n_629), .Y(n_659) );
NOR2x1_ASAP7_75t_L g660 ( .A(n_641), .B(n_651), .Y(n_660) );
NOR2x1_ASAP7_75t_L g661 ( .A(n_644), .B(n_630), .Y(n_661) );
NOR3xp33_ASAP7_75t_L g662 ( .A(n_633), .B(n_649), .C(n_642), .Y(n_662) );
NOR3xp33_ASAP7_75t_L g663 ( .A(n_658), .B(n_627), .C(n_646), .Y(n_663) );
AND2x4_ASAP7_75t_L g664 ( .A(n_657), .B(n_624), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_659), .B(n_622), .Y(n_665) );
NOR4xp75_ASAP7_75t_L g666 ( .A(n_656), .B(n_662), .C(n_661), .D(n_643), .Y(n_666) );
NOR3x2_ASAP7_75t_L g667 ( .A(n_666), .B(n_660), .C(n_647), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_663), .B(n_626), .Y(n_668) );
NOR2x1_ASAP7_75t_L g669 ( .A(n_664), .B(n_640), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_668), .Y(n_670) );
INVx3_ASAP7_75t_SL g671 ( .A(n_667), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_670), .Y(n_672) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_671), .Y(n_673) );
AO22x2_ASAP7_75t_L g674 ( .A1(n_672), .A2(n_664), .B1(n_665), .B2(n_673), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_673), .Y(n_675) );
OAI21xp5_ASAP7_75t_SL g676 ( .A1(n_675), .A2(n_669), .B(n_650), .Y(n_676) );
OAI222xp33_ASAP7_75t_L g677 ( .A1(n_676), .A2(n_674), .B1(n_645), .B2(n_636), .C1(n_623), .C2(n_631), .Y(n_677) );
AOI22x1_ASAP7_75t_L g678 ( .A1(n_677), .A2(n_647), .B1(n_648), .B2(n_637), .Y(n_678) );
AOI21xp33_ASAP7_75t_SL g679 ( .A1(n_678), .A2(n_621), .B(n_653), .Y(n_679) );
endmodule