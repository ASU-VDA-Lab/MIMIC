module real_jpeg_12085_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_416, n_6, n_415, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_416;
input n_6;
input n_415;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_0),
.Y(n_111)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_3),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_3),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_3),
.B(n_32),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_3),
.B(n_29),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_3),
.B(n_53),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_3),
.B(n_40),
.Y(n_277)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_5),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_5),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_5),
.B(n_29),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_5),
.B(n_53),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_5),
.B(n_40),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_5),
.B(n_111),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_5),
.B(n_116),
.Y(n_138)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_5),
.Y(n_346)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_6),
.Y(n_107)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_7),
.B(n_40),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_7),
.B(n_111),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_7),
.B(n_116),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_7),
.B(n_26),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_7),
.B(n_29),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_8),
.B(n_29),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_8),
.B(n_53),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_8),
.B(n_26),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_8),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_8),
.B(n_40),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_12),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_12),
.B(n_45),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_12),
.B(n_116),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_12),
.B(n_32),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_12),
.B(n_26),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_13),
.B(n_26),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_13),
.B(n_29),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_13),
.B(n_116),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_13),
.B(n_32),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_13),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_13),
.B(n_53),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_13),
.B(n_40),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_13),
.B(n_45),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_14),
.B(n_32),
.Y(n_101)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_14),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_14),
.B(n_111),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_14),
.B(n_29),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_14),
.B(n_40),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_14),
.B(n_45),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_15),
.B(n_53),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_15),
.B(n_40),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_15),
.B(n_111),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_15),
.B(n_116),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_15),
.B(n_26),
.Y(n_249)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

O2A1O1Ixp33_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_80),
.B(n_345),
.C(n_411),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_90),
.B(n_410),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_78),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_21),
.B(n_78),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_64),
.C(n_65),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_22),
.B(n_408),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_48),
.C(n_55),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_23),
.B(n_398),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_35),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_24),
.B(n_37),
.C(n_41),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.C(n_31),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_25),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_60)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_25),
.B(n_57),
.C(n_62),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_25),
.A2(n_63),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_25),
.B(n_234),
.C(n_235),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_25),
.A2(n_31),
.B1(n_63),
.B2(n_183),
.Y(n_387)
);

INVx5_ASAP7_75t_SL g125 ( 
.A(n_26),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_28),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.Y(n_275)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_28),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_28),
.B(n_274),
.C(n_277),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_28),
.A2(n_278),
.B1(n_386),
.B2(n_387),
.Y(n_385)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_30),
.B(n_38),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_31),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_31),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_31),
.B(n_179),
.C(n_181),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_31),
.A2(n_137),
.B1(n_138),
.B2(n_183),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_31),
.B(n_137),
.C(n_249),
.Y(n_390)
);

CKINVDCx14_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_33),
.B(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_33),
.B(n_51),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_33),
.B(n_43),
.Y(n_253)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_37),
.B1(n_41),
.B2(n_42),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_38),
.B(n_110),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_43),
.B(n_228),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_44),
.B(n_158),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_44),
.B(n_112),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_44),
.B(n_346),
.Y(n_345)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_48),
.A2(n_55),
.B1(n_56),
.B2(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_48),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.C(n_52),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_49),
.B(n_52),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_84),
.B1(n_85),
.B2(n_88),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_50),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_50),
.A2(n_88),
.B1(n_382),
.B2(n_383),
.Y(n_381)
);

NOR3xp33_ASAP7_75t_L g411 ( 
.A(n_50),
.B(n_69),
.C(n_86),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_53),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_57),
.A2(n_58),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_58),
.B(n_118),
.C(n_234),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_61),
.A2(n_62),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_67),
.C(n_69),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_61),
.A2(n_62),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_62),
.B(n_247),
.C(n_249),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_64),
.B(n_65),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_73),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_75),
.C(n_76),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_71),
.B2(n_72),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_67),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_67),
.A2(n_71),
.B1(n_352),
.B2(n_353),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_67),
.B(n_354),
.C(n_355),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_68),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_70),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_69),
.A2(n_70),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_70),
.B(n_288),
.C(n_290),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_89),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_86),
.A2(n_87),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_87),
.B(n_310),
.C(n_313),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_405),
.B(n_409),
.Y(n_90)
);

OAI321xp33_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_371),
.A3(n_392),
.B1(n_403),
.B2(n_404),
.C(n_415),
.Y(n_91)
);

AOI321xp33_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_299),
.A3(n_331),
.B1(n_365),
.B2(n_370),
.C(n_416),
.Y(n_92)
);

NOR3xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_238),
.C(n_294),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_206),
.B(n_237),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_173),
.B(n_205),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_142),
.B(n_172),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_119),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_98),
.B(n_119),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.C(n_113),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_122),
.B1(n_123),
.B2(n_131),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_99),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_99),
.B(n_169),
.Y(n_168)
);

FAx1_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_101),
.CI(n_102),
.CON(n_99),
.SN(n_99)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_103),
.A2(n_104),
.B1(n_113),
.B2(n_170),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_105),
.B(n_109),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.Y(n_105)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_106),
.B(n_158),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_108),
.B(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_110),
.B(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_112),
.B(n_125),
.Y(n_179)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_117),
.B2(n_118),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_114),
.B(n_118),
.Y(n_133)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_117),
.A2(n_118),
.B1(n_187),
.B2(n_188),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_117),
.A2(n_118),
.B1(n_233),
.B2(n_234),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_118),
.B(n_188),
.C(n_291),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_132),
.B2(n_141),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_122),
.B(n_131),
.C(n_141),
.Y(n_174)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_124),
.B(n_127),
.C(n_130),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_129),
.Y(n_130)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_133),
.B(n_135),
.C(n_136),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_137),
.A2(n_138),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_137),
.A2(n_138),
.B1(n_344),
.B2(n_345),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_137),
.B(n_345),
.C(n_347),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_138),
.B(n_139),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_138),
.B(n_326),
.C(n_328),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_139),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_139),
.A2(n_140),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_139),
.B(n_261),
.C(n_264),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_166),
.B(n_171),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_155),
.B(n_165),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_150),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_145),
.B(n_150),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_153),
.C(n_154),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_160),
.B(n_164),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_157),
.B(n_159),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_167),
.B(n_168),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_174),
.B(n_175),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_191),
.B2(n_192),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_193),
.C(n_204),
.Y(n_207)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_184),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_185),
.C(n_186),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_188),
.B(n_189),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_203),
.B2(n_204),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_202),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_199),
.C(n_201),
.Y(n_225)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_197),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_198),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_207),
.B(n_208),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_224),
.B2(n_236),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_223),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_211),
.B(n_223),
.C(n_236),
.Y(n_295)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_213),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_219),
.B2(n_220),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_214),
.B(n_221),
.C(n_222),
.Y(n_257)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx24_ASAP7_75t_SL g414 ( 
.A(n_215),
.Y(n_414)
);

FAx1_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_217),
.CI(n_218),
.CON(n_215),
.SN(n_215)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_216),
.B(n_217),
.C(n_218),
.Y(n_266)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_224),
.Y(n_236)
);

BUFx24_ASAP7_75t_SL g413 ( 
.A(n_224),
.Y(n_413)
);

FAx1_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_226),
.CI(n_231),
.CON(n_224),
.SN(n_224)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_225),
.B(n_226),
.C(n_231),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_229),
.B(n_230),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_229),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_230),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_265)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_230),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_235),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_233),
.Y(n_234)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

AOI21xp33_ASAP7_75t_L g366 ( 
.A1(n_239),
.A2(n_367),
.B(n_368),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_270),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_240),
.B(n_270),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_258),
.C(n_269),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_241),
.B(n_297),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_257),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_250),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_243),
.B(n_250),
.C(n_257),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_248),
.B2(n_249),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_246),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_248),
.A2(n_249),
.B1(n_360),
.B2(n_361),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_256),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_253),
.B(n_254),
.C(n_256),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_258),
.A2(n_259),
.B1(n_269),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_265),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_266),
.C(n_268),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_263),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_266),
.Y(n_267)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_269),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_293),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_282),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_272),
.B(n_282),
.C(n_293),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_279),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_273),
.B(n_280),
.C(n_281),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_283),
.B(n_285),
.C(n_286),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_290),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_288),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_295),
.B(n_296),
.Y(n_367)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_300),
.A2(n_366),
.B(n_369),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_301),
.B(n_302),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_330),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_304),
.B(n_305),
.C(n_330),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_322),
.B2(n_323),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_306),
.B(n_324),
.C(n_325),
.Y(n_364)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_314),
.B2(n_315),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_308),
.B(n_316),
.C(n_321),
.Y(n_337)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_320),
.B2(n_321),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_318),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_328),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_332),
.B(n_333),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_364),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_349),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_335),
.B(n_349),
.C(n_364),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_337),
.B1(n_338),
.B2(n_339),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_336),
.B(n_340),
.C(n_348),
.Y(n_391)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_348),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_341),
.A2(n_342),
.B1(n_343),
.B2(n_347),
.Y(n_340)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_341),
.Y(n_347)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_351),
.B1(n_356),
.B2(n_357),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_350),
.B(n_358),
.C(n_363),
.Y(n_375)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

CKINVDCx14_ASAP7_75t_R g352 ( 
.A(n_353),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_358),
.A2(n_359),
.B1(n_362),
.B2(n_363),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_363),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_372),
.B(n_373),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_391),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_375),
.B(n_376),
.C(n_391),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_384),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_378),
.A2(n_379),
.B1(n_380),
.B2(n_381),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_378),
.B(n_381),
.C(n_384),
.Y(n_402)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_382),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_385),
.B(n_388),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_385),
.B(n_389),
.C(n_390),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_387),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_390),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_394),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_393),
.B(n_394),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_402),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_397),
.B1(n_400),
.B2(n_401),
.Y(n_395)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_396),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_396),
.B(n_401),
.C(n_402),
.Y(n_406)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_397),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_406),
.B(n_407),
.Y(n_409)
);


endmodule