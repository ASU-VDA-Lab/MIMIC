module fake_jpeg_27462_n_224 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_224);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_8),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_36),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_25),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_35),
.A2(n_18),
.B1(n_27),
.B2(n_21),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_19),
.B(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_39),
.Y(n_54)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_38),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_42),
.B(n_28),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_38),
.A2(n_29),
.B1(n_25),
.B2(n_30),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_44),
.B1(n_52),
.B2(n_42),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_38),
.A2(n_29),
.B1(n_25),
.B2(n_30),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_26),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_28),
.Y(n_66)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

OA21x2_ASAP7_75t_L g86 ( 
.A1(n_48),
.A2(n_20),
.B(n_28),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_51),
.B(n_53),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_33),
.A2(n_29),
.B1(n_30),
.B2(n_26),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_33),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_56),
.A2(n_20),
.B1(n_18),
.B2(n_40),
.Y(n_78)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_58),
.Y(n_81)
);

INVxp33_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_60),
.Y(n_90)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_62),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_39),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_65),
.Y(n_103)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_57),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_66),
.B(n_80),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_67),
.B(n_75),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_35),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_69),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_71),
.B(n_74),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_40),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_82),
.Y(n_107)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_45),
.B(n_21),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_47),
.B1(n_58),
.B2(n_57),
.Y(n_89)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_50),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_50),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_28),
.Y(n_85)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_74),
.A2(n_68),
.B1(n_72),
.B2(n_77),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_88),
.A2(n_105),
.B1(n_81),
.B2(n_79),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_89),
.A2(n_23),
.B1(n_17),
.B2(n_16),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_70),
.A2(n_47),
.B1(n_52),
.B2(n_58),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_91),
.A2(n_71),
.B1(n_83),
.B2(n_60),
.Y(n_114)
);

A2O1A1O1Ixp25_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_46),
.B(n_44),
.C(n_41),
.D(n_16),
.Y(n_94)
);

AO21x1_ASAP7_75t_L g117 ( 
.A1(n_94),
.A2(n_82),
.B(n_73),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_46),
.C(n_41),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_104),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_32),
.C(n_31),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_69),
.A2(n_47),
.B1(n_32),
.B2(n_31),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_86),
.A2(n_1),
.B(n_2),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_110),
.A2(n_81),
.B(n_84),
.Y(n_116)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_76),
.Y(n_113)
);

AO22x1_ASAP7_75t_SL g112 ( 
.A1(n_88),
.A2(n_86),
.B1(n_65),
.B2(n_67),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_122),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_113),
.A2(n_116),
.B(n_119),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_123),
.B1(n_128),
.B2(n_133),
.Y(n_141)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_115),
.B(n_118),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_129),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_64),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_22),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_120),
.B(n_129),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_23),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_111),
.A2(n_61),
.B1(n_65),
.B2(n_31),
.Y(n_123)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_2),
.Y(n_124)
);

NOR4xp25_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_127),
.C(n_16),
.D(n_22),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_73),
.B(n_4),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_131),
.B(n_3),
.Y(n_156)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_126),
.B(n_132),
.Y(n_143)
);

OR2x2_ASAP7_75t_SL g127 ( 
.A(n_106),
.B(n_98),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_99),
.A2(n_32),
.B1(n_31),
.B2(n_17),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_98),
.A2(n_22),
.B1(n_17),
.B2(n_32),
.Y(n_129)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_101),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_108),
.A2(n_73),
.B(n_6),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_109),
.A2(n_87),
.B1(n_105),
.B2(n_97),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_134),
.A2(n_100),
.B1(n_109),
.B2(n_104),
.Y(n_138)
);

AOI221xp5_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_110),
.B1(n_87),
.B2(n_109),
.C(n_106),
.Y(n_135)
);

NAND3xp33_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_151),
.C(n_127),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_137),
.B(n_145),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_156),
.B1(n_118),
.B2(n_116),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_91),
.C(n_90),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_146),
.C(n_150),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_113),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_95),
.C(n_102),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_92),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_155),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_122),
.Y(n_148)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_95),
.C(n_102),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_120),
.B(n_89),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_152),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_112),
.B(n_93),
.Y(n_154)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_93),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_157),
.B(n_160),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_114),
.B1(n_119),
.B2(n_123),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_161),
.A2(n_171),
.B1(n_141),
.B2(n_144),
.Y(n_183)
);

OA21x2_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_131),
.B(n_125),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_163),
.A2(n_155),
.B(n_139),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_143),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_164),
.B(n_168),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_165),
.A2(n_173),
.B1(n_137),
.B2(n_151),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_139),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_152),
.A2(n_119),
.B1(n_128),
.B2(n_23),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_141),
.A2(n_16),
.B1(n_7),
.B2(n_8),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_6),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_147),
.Y(n_182)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_179),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_169),
.Y(n_177)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_177),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_153),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_180),
.B(n_184),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_185),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_183),
.A2(n_172),
.B1(n_162),
.B2(n_159),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_167),
.B(n_144),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_150),
.Y(n_185)
);

XOR2x2_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_163),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_158),
.B(n_140),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_166),
.C(n_174),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_191),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_166),
.C(n_158),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_196),
.C(n_175),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_194),
.A2(n_157),
.B(n_176),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_186),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_159),
.C(n_148),
.Y(n_196)
);

BUFx24_ASAP7_75t_SL g198 ( 
.A(n_190),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_199),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_200),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g210 ( 
.A1(n_201),
.A2(n_202),
.B(n_204),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_196),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_203),
.A2(n_205),
.B(n_142),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_181),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_193),
.A2(n_163),
.B(n_172),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_178),
.C(n_183),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_206),
.A2(n_194),
.B(n_192),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_208),
.B(n_212),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_7),
.Y(n_215)
);

AOI322xp5_ASAP7_75t_L g212 ( 
.A1(n_206),
.A2(n_177),
.A3(n_179),
.B1(n_171),
.B2(n_142),
.C1(n_11),
.C2(n_12),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_207),
.A2(n_199),
.B(n_201),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_213),
.A2(n_215),
.B(n_216),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_177),
.C(n_8),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_9),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_211),
.A2(n_9),
.B(n_10),
.Y(n_216)
);

A2O1A1O1Ixp25_ASAP7_75t_L g219 ( 
.A1(n_217),
.A2(n_209),
.B(n_10),
.C(n_11),
.D(n_12),
.Y(n_219)
);

AOI322xp5_ASAP7_75t_L g222 ( 
.A1(n_219),
.A2(n_220),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.C1(n_51),
.C2(n_216),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_218),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_221),
.B(n_222),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_13),
.Y(n_224)
);


endmodule