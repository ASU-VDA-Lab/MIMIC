module fake_jpeg_11025_n_239 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_239);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_239;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_0),
.B(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx5p33_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_16),
.B(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_44),
.B(n_52),
.Y(n_86)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_20),
.A2(n_23),
.B(n_36),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_49),
.B(n_26),
.C(n_30),
.Y(n_116)
);

BUFx24_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_16),
.B(n_0),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_53),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_23),
.A2(n_2),
.B(n_3),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_58),
.Y(n_98)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_2),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_60),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_68),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_33),
.B(n_5),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_67),
.B(n_70),
.Y(n_87)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_6),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_42),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_5),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_71),
.B(n_72),
.Y(n_102)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_75),
.Y(n_99)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_81),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_17),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_78),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_17),
.B(n_38),
.Y(n_78)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_79),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_18),
.B(n_6),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_80),
.B(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_18),
.B(n_6),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_43),
.A2(n_29),
.B1(n_35),
.B2(n_34),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_85),
.A2(n_93),
.B1(n_83),
.B2(n_90),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_52),
.A2(n_29),
.B1(n_35),
.B2(n_34),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_94),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_50),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_96),
.B(n_107),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_67),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_48),
.A2(n_27),
.B1(n_32),
.B2(n_22),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_109),
.A2(n_114),
.B1(n_115),
.B2(n_47),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_53),
.A2(n_32),
.B1(n_19),
.B2(n_22),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_55),
.A2(n_19),
.B1(n_26),
.B2(n_30),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_117),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_71),
.B(n_38),
.C(n_37),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_118),
.C(n_7),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_44),
.A2(n_37),
.B(n_7),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_65),
.A2(n_7),
.B1(n_70),
.B2(n_61),
.Y(n_119)
);

AO21x1_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_100),
.B(n_91),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_58),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_123),
.B(n_44),
.Y(n_158)
);

OAI32xp33_ASAP7_75t_L g125 ( 
.A1(n_98),
.A2(n_74),
.A3(n_73),
.B1(n_60),
.B2(n_54),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_128),
.Y(n_166)
);

NAND2x1_ASAP7_75t_L g183 ( 
.A(n_126),
.B(n_158),
.Y(n_183)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_86),
.B(n_82),
.Y(n_129)
);

NAND3xp33_ASAP7_75t_L g167 ( 
.A(n_129),
.B(n_152),
.C(n_156),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_82),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_136),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_85),
.A2(n_54),
.B1(n_75),
.B2(n_110),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_131),
.A2(n_141),
.B1(n_147),
.B2(n_148),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_87),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_134),
.Y(n_170)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_116),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_99),
.Y(n_135)
);

XOR2x1_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_150),
.Y(n_169)
);

OAI32xp33_ASAP7_75t_L g136 ( 
.A1(n_124),
.A2(n_101),
.A3(n_94),
.B1(n_113),
.B2(n_120),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_84),
.B(n_89),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_139),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_89),
.B(n_106),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_114),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_145),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_109),
.A2(n_119),
.B1(n_92),
.B2(n_88),
.Y(n_141)
);

AOI32xp33_ASAP7_75t_L g142 ( 
.A1(n_100),
.A2(n_92),
.A3(n_108),
.B1(n_104),
.B2(n_95),
.Y(n_142)
);

FAx1_ASAP7_75t_SL g178 ( 
.A(n_142),
.B(n_127),
.CI(n_143),
.CON(n_178),
.SN(n_178)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_104),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_100),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_149),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_122),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_83),
.B(n_90),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_88),
.B(n_121),
.C(n_95),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_157),
.C(n_160),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_155),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_107),
.B(n_123),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_107),
.B(n_117),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_107),
.B(n_98),
.Y(n_160)
);

AND2x6_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_134),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_178),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_148),
.A2(n_135),
.B1(n_132),
.B2(n_155),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_171),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_160),
.A2(n_161),
.B1(n_147),
.B2(n_128),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_161),
.A2(n_150),
.B1(n_151),
.B2(n_136),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_175),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_159),
.A2(n_126),
.B1(n_125),
.B2(n_137),
.Y(n_175)
);

AND2x6_ASAP7_75t_L g179 ( 
.A(n_133),
.B(n_152),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_175),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_144),
.B(n_126),
.C(n_134),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_182),
.Y(n_198)
);

BUFx12_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_187),
.Y(n_206)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

AO22x1_ASAP7_75t_SL g190 ( 
.A1(n_169),
.A2(n_153),
.B1(n_163),
.B2(n_174),
.Y(n_190)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_193),
.B(n_195),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_168),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_185),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_170),
.B(n_169),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_197),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_177),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_183),
.C(n_165),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_180),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_202),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_172),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_201),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_182),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_166),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_191),
.A2(n_176),
.B1(n_162),
.B2(n_181),
.Y(n_203)
);

OA21x2_ASAP7_75t_L g216 ( 
.A1(n_203),
.A2(n_208),
.B(n_214),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_194),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_213),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_191),
.A2(n_171),
.B1(n_178),
.B2(n_183),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_197),
.C(n_190),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_202),
.A2(n_178),
.B(n_173),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_215),
.B(n_198),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_219),
.C(n_222),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_201),
.Y(n_219)
);

OAI321xp33_ASAP7_75t_L g220 ( 
.A1(n_210),
.A2(n_200),
.A3(n_196),
.B1(n_188),
.B2(n_192),
.C(n_190),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_223),
.Y(n_230)
);

A2O1A1O1Ixp25_ASAP7_75t_L g221 ( 
.A1(n_213),
.A2(n_188),
.B(n_190),
.C(n_187),
.D(n_167),
.Y(n_221)
);

FAx1_ASAP7_75t_SL g227 ( 
.A(n_221),
.B(n_224),
.CI(n_173),
.CON(n_227),
.SN(n_227)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_187),
.C(n_165),
.Y(n_223)
);

FAx1_ASAP7_75t_SL g224 ( 
.A(n_212),
.B(n_208),
.CI(n_203),
.CON(n_224),
.SN(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_222),
.A2(n_209),
.B1(n_206),
.B2(n_204),
.Y(n_225)
);

AOI322xp5_ASAP7_75t_L g234 ( 
.A1(n_225),
.A2(n_227),
.A3(n_221),
.B1(n_224),
.B2(n_216),
.C1(n_214),
.C2(n_194),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_223),
.A2(n_209),
.B1(n_187),
.B2(n_207),
.Y(n_226)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_226),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_218),
.A2(n_214),
.B(n_207),
.Y(n_229)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_229),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_217),
.C(n_219),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_234),
.A2(n_230),
.B(n_226),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_235),
.A2(n_236),
.B1(n_229),
.B2(n_231),
.Y(n_237)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_233),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_225),
.C(n_230),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_238),
.B(n_232),
.Y(n_239)
);


endmodule