module fake_jpeg_32085_n_368 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_368);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_368;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_25),
.B(n_35),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_43),
.B(n_48),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_25),
.B(n_14),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_51),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_45),
.Y(n_123)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_15),
.Y(n_47)
);

INVx5_ASAP7_75t_SL g126 ( 
.A(n_47),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_14),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_17),
.B(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_50),
.B(n_17),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_26),
.B(n_13),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_52),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_26),
.B(n_12),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_58),
.Y(n_89)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_34),
.B(n_11),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_35),
.B(n_11),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_59),
.B(n_60),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_20),
.B(n_10),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_72),
.Y(n_90)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx3_ASAP7_75t_SL g108 ( 
.A(n_66),
.Y(n_108)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_70),
.Y(n_86)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_26),
.B(n_9),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

BUFx10_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_78),
.Y(n_92)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_15),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_77),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_31),
.B(n_0),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_21),
.Y(n_98)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_15),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_81),
.Y(n_93)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_41),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_82),
.B(n_21),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_82),
.A2(n_41),
.B1(n_30),
.B2(n_22),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_83),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_54),
.B(n_36),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_85),
.B(n_98),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_50),
.A2(n_28),
.B1(n_27),
.B2(n_16),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_88),
.A2(n_119),
.B1(n_75),
.B2(n_68),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_39),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_95),
.B(n_104),
.Y(n_145)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_62),
.A2(n_42),
.B1(n_19),
.B2(n_37),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g170 ( 
.A1(n_96),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_47),
.A2(n_30),
.B1(n_22),
.B2(n_28),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_100),
.A2(n_105),
.B1(n_127),
.B2(n_55),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_39),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_57),
.B1(n_49),
.B2(n_69),
.Y(n_105)
);

NOR2x1_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_19),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_109),
.B(n_113),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_22),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_116),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_65),
.A2(n_30),
.B(n_22),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_114),
.A2(n_86),
.B(n_126),
.C(n_99),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_64),
.B(n_30),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_46),
.B(n_21),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_125),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_73),
.A2(n_28),
.B1(n_27),
.B2(n_16),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_45),
.B(n_30),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_77),
.A2(n_16),
.B1(n_27),
.B2(n_42),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_128),
.Y(n_177)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_37),
.B(n_33),
.C(n_21),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_132),
.B(n_149),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_124),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_135),
.B(n_144),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_136),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_67),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_137),
.B(n_141),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_138),
.Y(n_192)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_139),
.Y(n_196)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_140),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_98),
.B(n_33),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_142),
.A2(n_170),
.B1(n_126),
.B2(n_108),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_92),
.B(n_17),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_147),
.Y(n_180)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_107),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_96),
.B(n_17),
.Y(n_147)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_148),
.B(n_151),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_84),
.A2(n_21),
.B(n_17),
.C(n_52),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_89),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_150),
.A2(n_114),
.B(n_108),
.Y(n_190)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_96),
.A2(n_74),
.B1(n_66),
.B2(n_61),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_153),
.A2(n_154),
.B1(n_157),
.B2(n_158),
.Y(n_203)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_162),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_96),
.B(n_70),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_159),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_88),
.A2(n_56),
.B1(n_1),
.B2(n_3),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_117),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_85),
.B(n_4),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_99),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_121),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_161),
.Y(n_184)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_93),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_124),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_166),
.B(n_167),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_90),
.B(n_6),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_97),
.B(n_94),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_168),
.B(n_158),
.Y(n_216)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_171),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_111),
.Y(n_171)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_111),
.Y(n_172)
);

NAND2xp33_ASAP7_75t_SL g210 ( 
.A(n_172),
.B(n_173),
.Y(n_210)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_124),
.B(n_5),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_124),
.Y(n_198)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_122),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_118),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_156),
.A2(n_102),
.B1(n_106),
.B2(n_110),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_186),
.A2(n_193),
.B1(n_194),
.B2(n_204),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_190),
.B(n_216),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_147),
.A2(n_102),
.B1(n_106),
.B2(n_129),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_142),
.A2(n_129),
.B1(n_120),
.B2(n_86),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_143),
.B(n_131),
.C(n_130),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_195),
.B(n_213),
.C(n_190),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_163),
.B(n_5),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_197),
.B(n_212),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_200),
.Y(n_223)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_130),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_137),
.B(n_118),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_209),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_176),
.A2(n_120),
.B1(n_91),
.B2(n_115),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_207),
.A2(n_215),
.B1(n_194),
.B2(n_186),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_141),
.B(n_174),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_176),
.A2(n_162),
.B(n_154),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_170),
.B(n_159),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_212),
.B(n_173),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_132),
.A2(n_103),
.B(n_115),
.Y(n_213)
);

AOI32xp33_ASAP7_75t_L g214 ( 
.A1(n_152),
.A2(n_91),
.A3(n_103),
.B1(n_146),
.B2(n_145),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_133),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_170),
.A2(n_177),
.B1(n_149),
.B2(n_172),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_202),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_217),
.B(n_226),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_170),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_218),
.B(n_245),
.Y(n_274)
);

OAI22x1_ASAP7_75t_L g219 ( 
.A1(n_211),
.A2(n_150),
.B1(n_144),
.B2(n_136),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_219),
.A2(n_221),
.B1(n_215),
.B2(n_193),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_220),
.A2(n_181),
.B(n_192),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_203),
.A2(n_171),
.B1(n_148),
.B2(n_155),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_224),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_160),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_225),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_197),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_182),
.Y(n_228)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_228),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_175),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_229),
.Y(n_263)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_196),
.Y(n_231)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_231),
.Y(n_253)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_232),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_248),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_187),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_236),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_189),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_180),
.C(n_201),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_191),
.B(n_140),
.Y(n_236)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_178),
.Y(n_238)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_185),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_239),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_207),
.A2(n_178),
.B1(n_210),
.B2(n_214),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_240),
.A2(n_244),
.B(n_195),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_241),
.A2(n_227),
.B1(n_218),
.B2(n_233),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_243),
.B(n_198),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_216),
.B(n_200),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_188),
.B(n_179),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_247),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_179),
.B(n_180),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_203),
.A2(n_201),
.B1(n_183),
.B2(n_189),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_266),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_254),
.A2(n_219),
.B1(n_222),
.B2(n_229),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_230),
.A2(n_183),
.B(n_213),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_255),
.A2(n_268),
.B(n_222),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_256),
.B(n_262),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_230),
.A2(n_210),
.B(n_185),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_258),
.Y(n_287)
);

AOI221xp5_ASAP7_75t_L g294 ( 
.A1(n_265),
.A2(n_275),
.B1(n_221),
.B2(n_229),
.C(n_232),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_237),
.B(n_185),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_224),
.Y(n_267)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_267),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_242),
.A2(n_199),
.B(n_184),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_228),
.Y(n_270)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_270),
.Y(n_296)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_231),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_271),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_237),
.B(n_199),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_223),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_244),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_276),
.B(n_278),
.C(n_281),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_235),
.C(n_272),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_297),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_223),
.C(n_248),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_239),
.Y(n_282)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_282),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_259),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_283),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_254),
.A2(n_227),
.B1(n_241),
.B2(n_218),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_284),
.A2(n_285),
.B1(n_252),
.B2(n_269),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_288),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_261),
.B(n_225),
.C(n_243),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_290),
.B(n_291),
.C(n_253),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_225),
.C(n_217),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_234),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_293),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_208),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_294),
.A2(n_268),
.B1(n_269),
.B2(n_274),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_251),
.B(n_238),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_295),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_255),
.A2(n_263),
.B(n_275),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_299),
.B(n_296),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_301),
.A2(n_312),
.B1(n_295),
.B2(n_289),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_276),
.B(n_266),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_309),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_283),
.A2(n_264),
.B1(n_265),
.B2(n_267),
.Y(n_306)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_306),
.Y(n_324)
);

XNOR2x1_ASAP7_75t_L g309 ( 
.A(n_278),
.B(n_258),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_291),
.B(n_264),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_314),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_311),
.B(n_299),
.C(n_302),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_284),
.A2(n_258),
.B1(n_271),
.B2(n_257),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_277),
.B(n_250),
.C(n_257),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_315),
.C(n_305),
.Y(n_318)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_282),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_277),
.B(n_250),
.C(n_253),
.Y(n_315)
);

AOI321xp33_ASAP7_75t_L g316 ( 
.A1(n_309),
.A2(n_288),
.A3(n_297),
.B1(n_281),
.B2(n_290),
.C(n_287),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_316),
.B(n_321),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_318),
.B(n_322),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_303),
.B(n_279),
.Y(n_319)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_319),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_312),
.A2(n_287),
.B(n_298),
.Y(n_320)
);

INVxp33_ASAP7_75t_L g337 ( 
.A(n_320),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_298),
.A2(n_285),
.B(n_279),
.Y(n_321)
);

NOR3xp33_ASAP7_75t_SL g323 ( 
.A(n_308),
.B(n_300),
.C(n_280),
.Y(n_323)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_323),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_302),
.A2(n_286),
.B(n_296),
.Y(n_326)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_326),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_305),
.B(n_315),
.C(n_313),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_330),
.C(n_311),
.Y(n_332)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_328),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_304),
.B(n_289),
.Y(n_329)
);

NAND4xp25_ASAP7_75t_SL g336 ( 
.A(n_329),
.B(n_307),
.C(n_314),
.D(n_286),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_332),
.B(n_338),
.C(n_327),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_336),
.B(n_320),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_318),
.B(n_260),
.C(n_249),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_324),
.A2(n_260),
.B1(n_249),
.B2(n_270),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_340),
.B(n_326),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_333),
.B(n_325),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_342),
.B(n_343),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_344),
.B(n_346),
.Y(n_351)
);

NAND2xp33_ASAP7_75t_SL g345 ( 
.A(n_334),
.B(n_323),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_345),
.A2(n_348),
.B1(n_332),
.B2(n_205),
.Y(n_356)
);

AOI31xp67_ASAP7_75t_SL g346 ( 
.A1(n_336),
.A2(n_316),
.A3(n_322),
.B(n_330),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_347),
.B(n_349),
.C(n_339),
.Y(n_355)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_331),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_338),
.B(n_317),
.C(n_321),
.Y(n_349)
);

AO21x1_ASAP7_75t_L g350 ( 
.A1(n_337),
.A2(n_317),
.B(n_208),
.Y(n_350)
);

AO21x1_ASAP7_75t_L g353 ( 
.A1(n_350),
.A2(n_340),
.B(n_192),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_350),
.A2(n_337),
.B1(n_335),
.B2(n_341),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_352),
.B(n_355),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_353),
.B(n_356),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_349),
.B(n_339),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_357),
.B(n_347),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_359),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_354),
.B(n_205),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_361),
.B(n_205),
.Y(n_363)
);

O2A1O1Ixp33_ASAP7_75t_L g362 ( 
.A1(n_358),
.A2(n_351),
.B(n_352),
.C(n_353),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_362),
.A2(n_357),
.B1(n_360),
.B2(n_364),
.Y(n_365)
);

INVxp33_ASAP7_75t_L g366 ( 
.A(n_363),
.Y(n_366)
);

BUFx24_ASAP7_75t_SL g367 ( 
.A(n_365),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_367),
.B(n_366),
.Y(n_368)
);


endmodule