module fake_jpeg_18599_n_201 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_201);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx8_ASAP7_75t_SL g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_21),
.Y(n_47)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

NAND2xp33_ASAP7_75t_SL g54 ( 
.A(n_39),
.B(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_40),
.B(n_29),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_29),
.C(n_22),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_36),
.C(n_41),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_29),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_47),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_19),
.B1(n_20),
.B2(n_28),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_53),
.B1(n_31),
.B2(n_27),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_17),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_33),
.A2(n_29),
.B1(n_19),
.B2(n_28),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_33),
.A2(n_19),
.B1(n_20),
.B2(n_28),
.Y(n_55)
);

AO22x2_ASAP7_75t_L g58 ( 
.A1(n_55),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_36),
.Y(n_78)
);

OR2x2_ASAP7_75t_SL g57 ( 
.A(n_55),
.B(n_15),
.Y(n_57)
);

XOR2x1_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_72),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_84),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_36),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_46),
.A2(n_34),
.B1(n_20),
.B2(n_35),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_60),
.A2(n_62),
.B1(n_63),
.B2(n_75),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_55),
.A2(n_37),
.B1(n_35),
.B2(n_41),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_15),
.B1(n_39),
.B2(n_27),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_71),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_15),
.Y(n_69)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_16),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_43),
.A2(n_16),
.B1(n_25),
.B2(n_26),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_16),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_80),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_74),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_49),
.A2(n_39),
.B1(n_25),
.B2(n_31),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_78),
.A2(n_23),
.B(n_2),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_54),
.A2(n_41),
.B1(n_26),
.B2(n_38),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_81),
.A2(n_87),
.B1(n_49),
.B2(n_30),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_82),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_83),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_44),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_42),
.A2(n_30),
.B(n_23),
.C(n_3),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_1),
.B(n_3),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_44),
.B(n_36),
.C(n_38),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_7),
.C(n_8),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_49),
.A2(n_36),
.B1(n_30),
.B2(n_23),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_90),
.A2(n_101),
.B(n_102),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_92),
.A2(n_104),
.B1(n_78),
.B2(n_58),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_82),
.A2(n_5),
.B(n_6),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_9),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_6),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_111),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_9),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_9),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_57),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_115),
.B(n_125),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_72),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_116),
.B(n_117),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_88),
.A2(n_58),
.B1(n_78),
.B2(n_59),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_119),
.B(n_123),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_88),
.A2(n_58),
.B1(n_76),
.B2(n_66),
.Y(n_120)
);

FAx1_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_90),
.CI(n_98),
.CON(n_147),
.SN(n_147)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

NOR2x1_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_85),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_122),
.B(n_124),
.Y(n_136)
);

NOR3xp33_ASAP7_75t_SL g123 ( 
.A(n_93),
.B(n_86),
.C(n_83),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_109),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_126),
.A2(n_132),
.B(n_108),
.Y(n_141)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_99),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_128),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_89),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_129),
.Y(n_140)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

A2O1A1O1Ixp25_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_80),
.B(n_70),
.C(n_64),
.D(n_65),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_77),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_110),
.C(n_90),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_107),
.B(n_92),
.C(n_97),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_139),
.B(n_141),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_106),
.B(n_102),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_121),
.A2(n_103),
.B1(n_99),
.B2(n_98),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_144),
.A2(n_131),
.B1(n_89),
.B2(n_61),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_147),
.A2(n_122),
.B1(n_132),
.B2(n_123),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_113),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_149),
.B(n_118),
.C(n_133),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_155),
.C(n_156),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_142),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_157),
.Y(n_166)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_137),
.Y(n_154)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_154),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_120),
.C(n_114),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_150),
.B(n_114),
.Y(n_157)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_117),
.C(n_124),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_136),
.C(n_139),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_142),
.Y(n_160)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_161),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_103),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_162),
.A2(n_163),
.B1(n_135),
.B2(n_134),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_165),
.A2(n_156),
.B1(n_158),
.B2(n_153),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_141),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_171),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_146),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_159),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_178),
.Y(n_185)
);

NAND3xp33_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_136),
.C(n_153),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_175),
.B(n_176),
.Y(n_188)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_148),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_170),
.C(n_171),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_166),
.A2(n_147),
.B1(n_161),
.B2(n_154),
.Y(n_180)
);

AOI322xp5_ASAP7_75t_L g183 ( 
.A1(n_180),
.A2(n_181),
.A3(n_147),
.B1(n_145),
.B2(n_163),
.C1(n_173),
.C2(n_168),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_164),
.A2(n_147),
.B(n_134),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_145),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_182),
.B(n_126),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_181),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_187),
.C(n_177),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_143),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_140),
.C(n_126),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_190),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_185),
.C(n_175),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_191),
.A2(n_13),
.B(n_14),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_192),
.A2(n_91),
.B1(n_11),
.B2(n_12),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_194),
.B(n_14),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_189),
.C(n_193),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_196),
.B(n_197),
.Y(n_198)
);

AOI21x1_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_193),
.B(n_91),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_10),
.C(n_178),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_10),
.Y(n_201)
);


endmodule