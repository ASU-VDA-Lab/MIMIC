module fake_netlist_1_5697_n_534 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_534);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_534;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_141;
wire n_119;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_295;
wire n_143;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_44), .Y(n_77) );
INVxp67_ASAP7_75t_SL g78 ( .A(n_63), .Y(n_78) );
BUFx6f_ASAP7_75t_L g79 ( .A(n_19), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_66), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_31), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_42), .Y(n_82) );
INVxp67_ASAP7_75t_SL g83 ( .A(n_46), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_68), .Y(n_84) );
BUFx10_ASAP7_75t_L g85 ( .A(n_58), .Y(n_85) );
CKINVDCx14_ASAP7_75t_R g86 ( .A(n_73), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_8), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_2), .Y(n_88) );
INVxp33_ASAP7_75t_SL g89 ( .A(n_70), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_30), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_52), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_17), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_45), .Y(n_93) );
INVxp67_ASAP7_75t_SL g94 ( .A(n_37), .Y(n_94) );
HB1xp67_ASAP7_75t_L g95 ( .A(n_23), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_39), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_17), .Y(n_97) );
INVxp67_ASAP7_75t_L g98 ( .A(n_11), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_75), .Y(n_99) );
INVx1_ASAP7_75t_SL g100 ( .A(n_16), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_6), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_43), .Y(n_102) );
BUFx5_ASAP7_75t_L g103 ( .A(n_22), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_56), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_67), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_20), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_29), .Y(n_107) );
INVxp67_ASAP7_75t_SL g108 ( .A(n_74), .Y(n_108) );
CKINVDCx14_ASAP7_75t_R g109 ( .A(n_51), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_8), .Y(n_110) );
OR2x2_ASAP7_75t_L g111 ( .A(n_9), .B(n_48), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_26), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_18), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_103), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_80), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_103), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_103), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_80), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_84), .Y(n_119) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_95), .B(n_0), .Y(n_120) );
NOR2xp33_ASAP7_75t_L g121 ( .A(n_77), .B(n_0), .Y(n_121) );
AND2x4_ASAP7_75t_L g122 ( .A(n_88), .B(n_1), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_84), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_102), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_102), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_85), .Y(n_126) );
INVx3_ASAP7_75t_L g127 ( .A(n_85), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_104), .Y(n_128) );
INVx3_ASAP7_75t_L g129 ( .A(n_85), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_104), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_113), .Y(n_131) );
BUFx2_ASAP7_75t_L g132 ( .A(n_87), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_79), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_103), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_86), .B(n_1), .Y(n_135) );
NAND3x1_ASAP7_75t_L g136 ( .A(n_135), .B(n_88), .C(n_101), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_114), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_114), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g139 ( .A(n_126), .B(n_89), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_114), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_126), .B(n_87), .Y(n_141) );
AND2x2_ASAP7_75t_L g142 ( .A(n_132), .B(n_109), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_133), .Y(n_143) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_132), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_116), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_122), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_122), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_116), .Y(n_148) );
NAND3xp33_ASAP7_75t_L g149 ( .A(n_120), .B(n_98), .C(n_92), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g150 ( .A(n_126), .B(n_89), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_116), .Y(n_151) );
INVx4_ASAP7_75t_L g152 ( .A(n_122), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_117), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_117), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_117), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_134), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_134), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_134), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_122), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_115), .Y(n_160) );
INVx3_ASAP7_75t_L g161 ( .A(n_152), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_137), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_152), .B(n_126), .Y(n_163) );
INVx5_ASAP7_75t_L g164 ( .A(n_152), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_152), .Y(n_165) );
INVx3_ASAP7_75t_L g166 ( .A(n_146), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_146), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_159), .B(n_135), .Y(n_168) );
AOI22xp33_ASAP7_75t_L g169 ( .A1(n_159), .A2(n_118), .B1(n_123), .B2(n_131), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_137), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_160), .B(n_127), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_146), .Y(n_172) );
INVx2_ASAP7_75t_SL g173 ( .A(n_160), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_141), .B(n_127), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_138), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_146), .Y(n_176) );
INVx3_ASAP7_75t_L g177 ( .A(n_147), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_147), .Y(n_178) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_151), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_144), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_151), .Y(n_181) );
INVx3_ASAP7_75t_L g182 ( .A(n_147), .Y(n_182) );
BUFx3_ASAP7_75t_L g183 ( .A(n_147), .Y(n_183) );
OAI22xp5_ASAP7_75t_L g184 ( .A1(n_136), .A2(n_119), .B1(n_115), .B2(n_131), .Y(n_184) );
INVx3_ASAP7_75t_L g185 ( .A(n_153), .Y(n_185) );
OR2x6_ASAP7_75t_L g186 ( .A(n_136), .B(n_135), .Y(n_186) );
BUFx3_ASAP7_75t_L g187 ( .A(n_138), .Y(n_187) );
INVx2_ASAP7_75t_SL g188 ( .A(n_140), .Y(n_188) );
INVx3_ASAP7_75t_L g189 ( .A(n_153), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_140), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_145), .B(n_118), .Y(n_191) );
AND2x4_ASAP7_75t_L g192 ( .A(n_142), .B(n_127), .Y(n_192) );
AOI221xp5_ASAP7_75t_L g193 ( .A1(n_184), .A2(n_149), .B1(n_142), .B2(n_123), .C(n_128), .Y(n_193) );
OR2x6_ASAP7_75t_L g194 ( .A(n_186), .B(n_127), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_162), .Y(n_195) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_180), .Y(n_196) );
INVx6_ASAP7_75t_L g197 ( .A(n_164), .Y(n_197) );
BUFx12f_ASAP7_75t_L g198 ( .A(n_180), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_162), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_192), .B(n_169), .Y(n_200) );
INVx4_ASAP7_75t_L g201 ( .A(n_164), .Y(n_201) );
INVx1_ASAP7_75t_SL g202 ( .A(n_192), .Y(n_202) );
NAND2x1p5_ASAP7_75t_L g203 ( .A(n_164), .B(n_111), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_184), .A2(n_139), .B1(n_150), .B2(n_124), .Y(n_204) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_186), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_173), .A2(n_158), .B(n_145), .Y(n_206) );
BUFx2_ASAP7_75t_L g207 ( .A(n_164), .Y(n_207) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_186), .Y(n_208) );
BUFx2_ASAP7_75t_L g209 ( .A(n_164), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_186), .B(n_129), .Y(n_210) );
BUFx3_ASAP7_75t_L g211 ( .A(n_164), .Y(n_211) );
INVx3_ASAP7_75t_L g212 ( .A(n_187), .Y(n_212) );
BUFx2_ASAP7_75t_L g213 ( .A(n_164), .Y(n_213) );
AOI21xp33_ASAP7_75t_L g214 ( .A1(n_186), .A2(n_129), .B(n_92), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_186), .B(n_129), .Y(n_215) );
INVx4_ASAP7_75t_L g216 ( .A(n_164), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_192), .B(n_129), .Y(n_217) );
BUFx12f_ASAP7_75t_L g218 ( .A(n_186), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_162), .Y(n_219) );
AND2x4_ASAP7_75t_L g220 ( .A(n_192), .B(n_119), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_162), .Y(n_221) );
BUFx2_ASAP7_75t_L g222 ( .A(n_164), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_170), .B(n_124), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_173), .A2(n_158), .B(n_148), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_195), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_195), .B(n_170), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_199), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_214), .A2(n_168), .B(n_171), .C(n_174), .Y(n_228) );
OAI211xp5_ASAP7_75t_L g229 ( .A1(n_193), .A2(n_204), .B(n_196), .C(n_210), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_218), .A2(n_192), .B1(n_183), .B2(n_163), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_199), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_219), .Y(n_232) );
INVxp67_ASAP7_75t_L g233 ( .A(n_203), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_218), .A2(n_192), .B1(n_183), .B2(n_163), .Y(n_234) );
AOI221xp5_ASAP7_75t_L g235 ( .A1(n_220), .A2(n_168), .B1(n_169), .B2(n_174), .C(n_128), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_217), .Y(n_236) );
NAND3xp33_ASAP7_75t_L g237 ( .A(n_204), .B(n_171), .C(n_121), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_220), .Y(n_238) );
BUFx2_ASAP7_75t_L g239 ( .A(n_211), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_219), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_218), .A2(n_183), .B1(n_163), .B2(n_182), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_202), .A2(n_183), .B1(n_163), .B2(n_182), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_219), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_221), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_211), .B(n_163), .Y(n_245) );
OAI22xp33_ASAP7_75t_L g246 ( .A1(n_198), .A2(n_208), .B1(n_194), .B2(n_203), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_221), .Y(n_247) );
OAI22xp5_ASAP7_75t_L g248 ( .A1(n_203), .A2(n_173), .B1(n_188), .B2(n_175), .Y(n_248) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_194), .A2(n_188), .B1(n_175), .B2(n_170), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_220), .Y(n_250) );
AOI221xp5_ASAP7_75t_L g251 ( .A1(n_237), .A2(n_220), .B1(n_200), .B2(n_125), .C(n_130), .Y(n_251) );
OR2x2_ASAP7_75t_L g252 ( .A(n_233), .B(n_221), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g253 ( .A1(n_248), .A2(n_194), .B1(n_205), .B2(n_223), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_236), .A2(n_235), .B1(n_246), .B2(n_194), .Y(n_254) );
AOI221xp5_ASAP7_75t_L g255 ( .A1(n_229), .A2(n_125), .B1(n_130), .B2(n_210), .C(n_215), .Y(n_255) );
AOI21xp33_ASAP7_75t_L g256 ( .A1(n_228), .A2(n_194), .B(n_215), .Y(n_256) );
BUFx3_ASAP7_75t_L g257 ( .A(n_239), .Y(n_257) );
OAI211xp5_ASAP7_75t_SL g258 ( .A1(n_230), .A2(n_100), .B(n_97), .C(n_110), .Y(n_258) );
AOI221xp5_ASAP7_75t_L g259 ( .A1(n_238), .A2(n_215), .B1(n_223), .B2(n_101), .C(n_163), .Y(n_259) );
INVx6_ASAP7_75t_L g260 ( .A(n_245), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_249), .A2(n_212), .B1(n_215), .B2(n_190), .Y(n_261) );
CKINVDCx6p67_ASAP7_75t_R g262 ( .A(n_245), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_250), .A2(n_198), .B1(n_190), .B2(n_170), .Y(n_263) );
INVx3_ASAP7_75t_L g264 ( .A(n_245), .Y(n_264) );
AOI22xp33_ASAP7_75t_SL g265 ( .A1(n_239), .A2(n_198), .B1(n_222), .B2(n_209), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_225), .A2(n_190), .B1(n_175), .B2(n_212), .Y(n_266) );
AOI22xp33_ASAP7_75t_SL g267 ( .A1(n_225), .A2(n_207), .B1(n_222), .B2(n_209), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g268 ( .A1(n_226), .A2(n_175), .B(n_224), .C(n_206), .Y(n_268) );
OAI321xp33_ASAP7_75t_L g269 ( .A1(n_227), .A2(n_111), .A3(n_113), .B1(n_90), .B2(n_91), .C(n_93), .Y(n_269) );
INVx1_ASAP7_75t_SL g270 ( .A(n_226), .Y(n_270) );
OAI221xp5_ASAP7_75t_L g271 ( .A1(n_234), .A2(n_213), .B1(n_207), .B2(n_172), .C(n_178), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_232), .Y(n_272) );
OAI31xp33_ASAP7_75t_SL g273 ( .A1(n_265), .A2(n_231), .A3(n_227), .B(n_243), .Y(n_273) );
AOI221xp5_ASAP7_75t_L g274 ( .A1(n_258), .A2(n_231), .B1(n_244), .B2(n_243), .C(n_247), .Y(n_274) );
OAI22xp5_ASAP7_75t_L g275 ( .A1(n_254), .A2(n_247), .B1(n_244), .B2(n_240), .Y(n_275) );
NOR2x1_ASAP7_75t_L g276 ( .A(n_257), .B(n_240), .Y(n_276) );
NAND3xp33_ASAP7_75t_L g277 ( .A(n_255), .B(n_232), .C(n_79), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_270), .Y(n_278) );
AOI22xp33_ASAP7_75t_SL g279 ( .A1(n_253), .A2(n_213), .B1(n_211), .B2(n_107), .Y(n_279) );
INVx4_ASAP7_75t_L g280 ( .A(n_262), .Y(n_280) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_251), .A2(n_242), .B1(n_241), .B2(n_212), .Y(n_281) );
OAI22xp33_ASAP7_75t_L g282 ( .A1(n_252), .A2(n_212), .B1(n_82), .B2(n_107), .Y(n_282) );
OAI221xp5_ASAP7_75t_L g283 ( .A1(n_263), .A2(n_78), .B1(n_83), .B2(n_94), .C(n_96), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_272), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_264), .Y(n_285) );
INVxp67_ASAP7_75t_SL g286 ( .A(n_261), .Y(n_286) );
OAI211xp5_ASAP7_75t_L g287 ( .A1(n_263), .A2(n_99), .B(n_108), .C(n_82), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_264), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_266), .B(n_103), .Y(n_289) );
OAI22xp5_ASAP7_75t_L g290 ( .A1(n_254), .A2(n_188), .B1(n_187), .B2(n_216), .Y(n_290) );
INVxp67_ASAP7_75t_SL g291 ( .A(n_266), .Y(n_291) );
BUFx2_ASAP7_75t_L g292 ( .A(n_268), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_260), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_267), .B(n_191), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_284), .B(n_256), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_277), .A2(n_268), .B(n_269), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_292), .B(n_103), .Y(n_297) );
OAI221xp5_ASAP7_75t_L g298 ( .A1(n_273), .A2(n_259), .B1(n_260), .B2(n_271), .C(n_105), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_278), .B(n_260), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_292), .B(n_103), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_284), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_285), .B(n_288), .Y(n_302) );
OR2x6_ASAP7_75t_L g303 ( .A(n_276), .B(n_201), .Y(n_303) );
NOR3xp33_ASAP7_75t_L g304 ( .A(n_283), .B(n_106), .C(n_81), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_276), .Y(n_305) );
AND2x2_ASAP7_75t_SL g306 ( .A(n_280), .B(n_201), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_285), .Y(n_307) );
AOI221xp5_ASAP7_75t_L g308 ( .A1(n_289), .A2(n_81), .B1(n_112), .B2(n_79), .C(n_191), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_293), .B(n_2), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_288), .B(n_103), .Y(n_310) );
OAI221xp5_ASAP7_75t_SL g311 ( .A1(n_294), .A2(n_112), .B1(n_172), .B2(n_176), .C(n_167), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_277), .A2(n_79), .B1(n_172), .B2(n_216), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_280), .Y(n_313) );
OAI221xp5_ASAP7_75t_SL g314 ( .A1(n_294), .A2(n_176), .B1(n_178), .B2(n_167), .C(n_6), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_275), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_286), .Y(n_316) );
OAI33xp33_ASAP7_75t_L g317 ( .A1(n_282), .A2(n_3), .A3(n_4), .B1(n_5), .B2(n_7), .B3(n_9), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_291), .B(n_3), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_293), .B(n_4), .Y(n_319) );
OAI22xp5_ASAP7_75t_L g320 ( .A1(n_279), .A2(n_187), .B1(n_201), .B2(n_216), .Y(n_320) );
OAI221xp5_ASAP7_75t_L g321 ( .A1(n_287), .A2(n_79), .B1(n_201), .B2(n_216), .C(n_189), .Y(n_321) );
AOI221xp5_ASAP7_75t_L g322 ( .A1(n_289), .A2(n_133), .B1(n_166), .B2(n_177), .C(n_182), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_274), .B(n_5), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_301), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_301), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_307), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_307), .Y(n_327) );
INVx3_ASAP7_75t_L g328 ( .A(n_305), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_302), .B(n_133), .Y(n_329) );
INVx2_ASAP7_75t_SL g330 ( .A(n_313), .Y(n_330) );
INVx1_ASAP7_75t_SL g331 ( .A(n_313), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_302), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_295), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_310), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_310), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_295), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_316), .B(n_280), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_299), .B(n_281), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_305), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_297), .B(n_133), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_298), .B(n_7), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_316), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_315), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_297), .B(n_133), .Y(n_344) );
NOR3xp33_ASAP7_75t_L g345 ( .A(n_317), .B(n_290), .C(n_281), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_300), .B(n_133), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_315), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_300), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_318), .B(n_10), .Y(n_349) );
OAI221xp5_ASAP7_75t_L g350 ( .A1(n_314), .A2(n_197), .B1(n_189), .B2(n_185), .C(n_187), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_318), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_303), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_303), .Y(n_353) );
INVx1_ASAP7_75t_SL g354 ( .A(n_306), .Y(n_354) );
NAND2x1p5_ASAP7_75t_L g355 ( .A(n_306), .B(n_189), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_323), .B(n_10), .Y(n_356) );
AND2x4_ASAP7_75t_L g357 ( .A(n_303), .B(n_59), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_323), .B(n_11), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_303), .B(n_12), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_303), .B(n_12), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_309), .B(n_13), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_319), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_306), .B(n_13), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_296), .B(n_14), .Y(n_364) );
INVx3_ASAP7_75t_L g365 ( .A(n_312), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_320), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_324), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_328), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_351), .B(n_304), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_351), .B(n_308), .Y(n_370) );
CKINVDCx20_ASAP7_75t_R g371 ( .A(n_331), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_332), .B(n_322), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_331), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_342), .Y(n_374) );
INVx1_ASAP7_75t_SL g375 ( .A(n_330), .Y(n_375) );
INVx1_ASAP7_75t_SL g376 ( .A(n_330), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_342), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_332), .B(n_311), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_336), .B(n_14), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_336), .B(n_15), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_333), .B(n_15), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_324), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_356), .B(n_16), .Y(n_383) );
AND5x1_ASAP7_75t_L g384 ( .A(n_341), .B(n_321), .C(n_320), .D(n_25), .E(n_27), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_325), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_358), .B(n_21), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_333), .B(n_24), .Y(n_387) );
AND2x4_ASAP7_75t_SL g388 ( .A(n_357), .B(n_189), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_354), .B(n_179), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_325), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_343), .B(n_28), .Y(n_391) );
BUFx2_ASAP7_75t_L g392 ( .A(n_337), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_326), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_343), .B(n_32), .Y(n_394) );
NOR2xp67_ASAP7_75t_L g395 ( .A(n_359), .B(n_33), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_339), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_347), .B(n_34), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_347), .B(n_35), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_348), .B(n_36), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_339), .B(n_38), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_326), .Y(n_401) );
INVx1_ASAP7_75t_SL g402 ( .A(n_337), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_348), .B(n_40), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_352), .B(n_41), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_327), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_352), .B(n_353), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_327), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_353), .B(n_47), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_334), .B(n_49), .Y(n_409) );
INVx1_ASAP7_75t_SL g410 ( .A(n_360), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_362), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_362), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_329), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_329), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_338), .B(n_364), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_328), .Y(n_416) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_340), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_328), .Y(n_418) );
O2A1O1Ixp33_ASAP7_75t_L g419 ( .A1(n_369), .A2(n_383), .B(n_349), .C(n_361), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_392), .B(n_334), .Y(n_420) );
INVxp67_ASAP7_75t_L g421 ( .A(n_373), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_411), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_412), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_371), .B(n_364), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_392), .B(n_335), .Y(n_425) );
NOR3xp33_ASAP7_75t_SL g426 ( .A(n_415), .B(n_363), .C(n_366), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_402), .B(n_366), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_374), .Y(n_428) );
INVx3_ASAP7_75t_L g429 ( .A(n_368), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_377), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_396), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_396), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_371), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_375), .B(n_340), .Y(n_434) );
INVx1_ASAP7_75t_SL g435 ( .A(n_376), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_367), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_414), .B(n_344), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_367), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_410), .B(n_359), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_382), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_382), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_405), .Y(n_442) );
NAND2xp33_ASAP7_75t_SL g443 ( .A(n_417), .B(n_360), .Y(n_443) );
INVx2_ASAP7_75t_SL g444 ( .A(n_388), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_405), .B(n_393), .Y(n_445) );
AO211x2_ASAP7_75t_L g446 ( .A1(n_416), .A2(n_345), .B(n_355), .C(n_357), .Y(n_446) );
AOI221xp5_ASAP7_75t_L g447 ( .A1(n_370), .A2(n_344), .B1(n_346), .B2(n_365), .C(n_335), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_378), .A2(n_355), .B1(n_357), .B2(n_365), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_393), .B(n_346), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_395), .B(n_357), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_406), .B(n_365), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_388), .A2(n_355), .B(n_350), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_406), .B(n_50), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_401), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_401), .B(n_53), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_413), .B(n_54), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_381), .B(n_55), .Y(n_457) );
XNOR2x1_ASAP7_75t_L g458 ( .A(n_378), .B(n_57), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_381), .B(n_60), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_385), .Y(n_460) );
AOI331xp33_ASAP7_75t_L g461 ( .A1(n_386), .A2(n_418), .A3(n_416), .B1(n_384), .B2(n_372), .B3(n_379), .C1(n_380), .Y(n_461) );
XNOR2x1_ASAP7_75t_L g462 ( .A(n_380), .B(n_61), .Y(n_462) );
AOI32xp33_ASAP7_75t_L g463 ( .A1(n_403), .A2(n_165), .A3(n_161), .B1(n_185), .B2(n_189), .Y(n_463) );
AOI221xp5_ASAP7_75t_L g464 ( .A1(n_372), .A2(n_143), .B1(n_185), .B2(n_179), .C(n_181), .Y(n_464) );
BUFx2_ASAP7_75t_L g465 ( .A(n_413), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_403), .A2(n_197), .B1(n_166), .B2(n_182), .Y(n_466) );
AOI21xp33_ASAP7_75t_L g467 ( .A1(n_379), .A2(n_62), .B(n_64), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_407), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_407), .B(n_65), .Y(n_469) );
AOI322xp5_ASAP7_75t_L g470 ( .A1(n_394), .A2(n_177), .A3(n_166), .B1(n_182), .B2(n_161), .C1(n_165), .C2(n_185), .Y(n_470) );
NAND2x1_ASAP7_75t_L g471 ( .A(n_368), .B(n_197), .Y(n_471) );
AOI31xp33_ASAP7_75t_L g472 ( .A1(n_387), .A2(n_399), .A3(n_389), .B(n_409), .Y(n_472) );
A2O1A1O1Ixp25_ASAP7_75t_L g473 ( .A1(n_418), .A2(n_69), .B(n_71), .C(n_72), .D(n_76), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g474 ( .A1(n_394), .A2(n_197), .B1(n_177), .B2(n_166), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_385), .B(n_185), .Y(n_475) );
AOI221xp5_ASAP7_75t_L g476 ( .A1(n_390), .A2(n_143), .B1(n_181), .B2(n_179), .C(n_177), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_387), .A2(n_181), .B(n_179), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_390), .Y(n_478) );
AOI21xp33_ASAP7_75t_L g479 ( .A1(n_391), .A2(n_143), .B(n_181), .Y(n_479) );
XOR2x2_ASAP7_75t_L g480 ( .A(n_384), .B(n_148), .Y(n_480) );
OAI22xp33_ASAP7_75t_SL g481 ( .A1(n_399), .A2(n_161), .B1(n_165), .B2(n_166), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_400), .Y(n_482) );
OAI22xp5_ASAP7_75t_SL g483 ( .A1(n_368), .A2(n_161), .B1(n_165), .B2(n_177), .Y(n_483) );
BUFx2_ASAP7_75t_L g484 ( .A(n_404), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_400), .Y(n_485) );
AOI32xp33_ASAP7_75t_L g486 ( .A1(n_404), .A2(n_165), .A3(n_161), .B1(n_155), .B2(n_154), .Y(n_486) );
BUFx2_ASAP7_75t_L g487 ( .A(n_408), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_409), .A2(n_179), .B(n_181), .Y(n_488) );
OAI21xp33_ASAP7_75t_L g489 ( .A1(n_408), .A2(n_143), .B(n_179), .Y(n_489) );
INVxp67_ASAP7_75t_L g490 ( .A(n_397), .Y(n_490) );
OAI22xp33_ASAP7_75t_L g491 ( .A1(n_398), .A2(n_179), .B1(n_181), .B2(n_143), .Y(n_491) );
OAI221xp5_ASAP7_75t_L g492 ( .A1(n_415), .A2(n_179), .B1(n_181), .B2(n_154), .C(n_155), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_411), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_465), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_447), .B(n_421), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_451), .B(n_427), .Y(n_496) );
AOI21xp33_ASAP7_75t_L g497 ( .A1(n_419), .A2(n_458), .B(n_446), .Y(n_497) );
INVxp67_ASAP7_75t_L g498 ( .A(n_433), .Y(n_498) );
AOI221xp5_ASAP7_75t_L g499 ( .A1(n_424), .A2(n_448), .B1(n_426), .B2(n_443), .C(n_490), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_452), .A2(n_448), .B(n_435), .C(n_463), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_420), .B(n_425), .Y(n_501) );
INVx4_ASAP7_75t_SL g502 ( .A(n_483), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_439), .A2(n_435), .B1(n_462), .B2(n_484), .Y(n_503) );
BUFx2_ASAP7_75t_L g504 ( .A(n_429), .Y(n_504) );
OAI22xp33_ASAP7_75t_L g505 ( .A1(n_472), .A2(n_487), .B1(n_444), .B2(n_450), .Y(n_505) );
AOI211xp5_ASAP7_75t_SL g506 ( .A1(n_481), .A2(n_472), .B(n_492), .C(n_467), .Y(n_506) );
AOI221xp5_ASAP7_75t_L g507 ( .A1(n_493), .A2(n_422), .B1(n_423), .B2(n_430), .C(n_428), .Y(n_507) );
XNOR2x1_ASAP7_75t_L g508 ( .A(n_480), .B(n_434), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_437), .A2(n_429), .B1(n_471), .B2(n_449), .Y(n_509) );
NOR2x1p5_ASAP7_75t_L g510 ( .A(n_482), .B(n_485), .Y(n_510) );
OAI322xp33_ASAP7_75t_L g511 ( .A1(n_505), .A2(n_449), .A3(n_459), .B1(n_457), .B2(n_445), .C1(n_432), .C2(n_431), .Y(n_511) );
OAI21xp5_ASAP7_75t_SL g512 ( .A1(n_497), .A2(n_486), .B(n_466), .Y(n_512) );
INVxp67_ASAP7_75t_L g513 ( .A(n_508), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_498), .Y(n_514) );
NAND4xp25_ASAP7_75t_L g515 ( .A(n_506), .B(n_470), .C(n_474), .D(n_464), .Y(n_515) );
AOI211xp5_ASAP7_75t_L g516 ( .A1(n_500), .A2(n_489), .B(n_453), .C(n_477), .Y(n_516) );
AOI221xp5_ASAP7_75t_L g517 ( .A1(n_499), .A2(n_442), .B1(n_441), .B2(n_436), .C(n_438), .Y(n_517) );
AOI222xp33_ASAP7_75t_L g518 ( .A1(n_502), .A2(n_440), .B1(n_445), .B2(n_468), .C1(n_454), .C2(n_478), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_495), .A2(n_461), .B(n_488), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_514), .Y(n_520) );
NOR4xp25_ASAP7_75t_L g521 ( .A(n_513), .B(n_509), .C(n_507), .D(n_494), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_515), .A2(n_502), .B1(n_503), .B2(n_510), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_518), .Y(n_523) );
NAND4xp25_ASAP7_75t_L g524 ( .A(n_517), .B(n_504), .C(n_456), .D(n_496), .Y(n_524) );
OAI221xp5_ASAP7_75t_L g525 ( .A1(n_522), .A2(n_512), .B1(n_519), .B2(n_516), .C(n_511), .Y(n_525) );
NOR2x1_ASAP7_75t_L g526 ( .A(n_520), .B(n_455), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_522), .B(n_501), .Y(n_527) );
AND3x4_ASAP7_75t_L g528 ( .A(n_525), .B(n_521), .C(n_523), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_527), .A2(n_524), .B1(n_460), .B2(n_455), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_528), .A2(n_526), .B1(n_491), .B2(n_475), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_529), .A2(n_469), .B1(n_479), .B2(n_476), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_530), .Y(n_532) );
AOI21xp33_ASAP7_75t_L g533 ( .A1(n_532), .A2(n_531), .B(n_479), .Y(n_533) );
AOI221xp5_ASAP7_75t_L g534 ( .A1(n_533), .A2(n_473), .B1(n_181), .B2(n_157), .C(n_156), .Y(n_534) );
endmodule