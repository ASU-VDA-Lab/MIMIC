module fake_jpeg_4957_n_142 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_142);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_19),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_27),
.Y(n_48)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_35),
.Y(n_40)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_31),
.Y(n_39)
);

INVx5_ASAP7_75t_SL g31 ( 
.A(n_25),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_25),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_34),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_42),
.Y(n_50)
);

NOR2x1_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_46),
.Y(n_51)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_29),
.A2(n_23),
.B1(n_20),
.B2(n_14),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_15),
.B1(n_17),
.B2(n_23),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_28),
.A2(n_32),
.B1(n_30),
.B2(n_20),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_34),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_29),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_27),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_52),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_63),
.Y(n_83)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_56),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_59),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_45),
.A2(n_15),
.B1(n_14),
.B2(n_17),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_64),
.B1(n_48),
.B2(n_22),
.Y(n_73)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_39),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_60),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_21),
.Y(n_62)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_78),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_26),
.B1(n_19),
.B2(n_57),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_46),
.C(n_38),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_76),
.A2(n_77),
.B(n_79),
.Y(n_94)
);

OAI32xp33_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_33),
.A3(n_18),
.B1(n_26),
.B2(n_22),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_59),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_24),
.B1(n_13),
.B2(n_21),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_60),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_82),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_83),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_86),
.B1(n_95),
.B2(n_70),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_54),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_89),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_76),
.A2(n_44),
.B1(n_66),
.B2(n_39),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_91),
.B1(n_92),
.B2(n_67),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_40),
.Y(n_89)
);

NOR4xp25_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_11),
.C(n_9),
.D(n_7),
.Y(n_90)
);

AOI322xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_68),
.A3(n_7),
.B1(n_9),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_69),
.A2(n_37),
.B1(n_13),
.B2(n_35),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_80),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_74),
.Y(n_99)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_67),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_84),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_98),
.B(n_108),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_101),
.C(n_86),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_87),
.A2(n_74),
.B(n_72),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_103),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_107),
.Y(n_115)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_81),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_109),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_85),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_117),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_94),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_104),
.C(n_114),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_111),
.B(n_92),
.Y(n_120)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_121),
.A2(n_122),
.B(n_112),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_118),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_116),
.A2(n_100),
.B1(n_99),
.B2(n_107),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_125),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_117),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_125),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_128),
.A2(n_123),
.B(n_24),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_132),
.C(n_133),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_129),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_130),
.B(n_110),
.Y(n_133)
);

AOI31xp67_ASAP7_75t_SL g136 ( 
.A1(n_134),
.A2(n_130),
.A3(n_13),
.B(n_6),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_SL g139 ( 
.A(n_136),
.B(n_2),
.C(n_3),
.Y(n_139)
);

AO21x1_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_0),
.B(n_1),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_0),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_139),
.C(n_2),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_135),
.B(n_80),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_21),
.Y(n_142)
);


endmodule