module fake_aes_9424_n_1214 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_345, n_236, n_340, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_331, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_54, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_344, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_346, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_343, n_127, n_291, n_170, n_281, n_341, n_58, n_122, n_187, n_138, n_323, n_347, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_332, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1214);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_236;
input n_340;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_331;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_344;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_346;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_343;
input n_127;
input n_291;
input n_170;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_347;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1214;
wire n_1173;
wire n_663;
wire n_707;
wire n_791;
wire n_513;
wire n_361;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_1024;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_1198;
wire n_484;
wire n_852;
wire n_862;
wire n_667;
wire n_496;
wire n_801;
wire n_988;
wire n_1059;
wire n_1158;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_1202;
wire n_464;
wire n_965;
wire n_448;
wire n_1196;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_1211;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_1122;
wire n_528;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_1128;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_1175;
wire n_853;
wire n_1161;
wire n_987;
wire n_1030;
wire n_765;
wire n_1177;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_545;
wire n_896;
wire n_1185;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_1197;
wire n_1163;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_1200;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_1090;
wire n_1201;
wire n_1191;
wire n_1121;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_1194;
wire n_694;
wire n_1179;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_1174;
wire n_1005;
wire n_951;
wire n_702;
wire n_1016;
wire n_1097;
wire n_1078;
wire n_572;
wire n_1017;
wire n_1125;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_1169;
wire n_1204;
wire n_652;
wire n_975;
wire n_1042;
wire n_968;
wire n_1060;
wire n_437;
wire n_512;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_955;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_1183;
wire n_567;
wire n_809;
wire n_888;
wire n_1188;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_529;
wire n_455;
wire n_1025;
wire n_1011;
wire n_1132;
wire n_1159;
wire n_1101;
wire n_1155;
wire n_630;
wire n_511;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_1180;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_624;
wire n_426;
wire n_769;
wire n_725;
wire n_818;
wire n_844;
wire n_1160;
wire n_1184;
wire n_1018;
wire n_1195;
wire n_738;
wire n_979;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1138;
wire n_1063;
wire n_506;
wire n_533;
wire n_490;
wire n_393;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_399;
wire n_892;
wire n_1171;
wire n_665;
wire n_571;
wire n_1154;
wire n_459;
wire n_863;
wire n_1062;
wire n_708;
wire n_907;
wire n_634;
wire n_610;
wire n_730;
wire n_1212;
wire n_696;
wire n_735;
wire n_771;
wire n_1091;
wire n_1203;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_935;
wire n_427;
wire n_1046;
wire n_950;
wire n_460;
wire n_910;
wire n_478;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_485;
wire n_703;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_699;
wire n_519;
wire n_729;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_1145;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_1167;
wire n_864;
wire n_1186;
wire n_810;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_1147;
wire n_1206;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_685;
wire n_362;
wire n_1178;
wire n_1209;
wire n_931;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1210;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_1176;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_649;
wire n_1047;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_446;
wire n_420;
wire n_621;
wire n_666;
wire n_423;
wire n_799;
wire n_880;
wire n_1089;
wire n_1058;
wire n_370;
wire n_1050;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_937;
wire n_874;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_970;
wire n_1181;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_806;
wire n_1066;
wire n_539;
wire n_1157;
wire n_1055;
wire n_974;
wire n_1153;
wire n_591;
wire n_933;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_1199;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_899;
wire n_654;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_1144;
wire n_677;
wire n_1023;
wire n_503;
wire n_756;
wire n_520;
wire n_1057;
wire n_1152;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_1149;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_1170;
wire n_419;
wire n_1193;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1133;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_1110;
wire n_1131;
wire n_1102;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_1208;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_1156;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_924;
wire n_912;
wire n_1043;
wire n_947;
wire n_582;
wire n_378;
wire n_1141;
wire n_1213;
wire n_359;
wire n_441;
wire n_836;
wire n_1189;
wire n_923;
wire n_1205;
wire n_561;
wire n_1096;
wire n_1172;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1142;
wire n_1109;
wire n_1008;
wire n_1026;
wire n_766;
wire n_602;
wire n_831;
wire n_1027;
wire n_1007;
wire n_859;
wire n_1117;
wire n_1040;
wire n_1165;
wire n_930;
wire n_994;
wire n_1182;
wire n_424;
wire n_714;
wire n_1143;
wire n_629;
wire n_569;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_1207;
wire n_867;
wire n_1070;
wire n_1168;
wire n_377;
wire n_510;
wire n_1112;
wire n_1075;
wire n_675;
wire n_967;
wire n_504;
wire n_581;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_1164;
wire n_1038;
wire n_1162;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_1073;
wire n_473;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_1150;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_695;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_1104;
wire n_1187;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_1190;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_1146;
wire n_606;
wire n_425;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_1192;
wire n_433;
wire n_983;
wire n_1137;
wire n_781;
wire n_916;
wire n_421;
wire n_1148;
wire n_709;
wire n_739;
wire n_1166;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_819;
wire n_405;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_992;
wire n_1127;
INVx1_ASAP7_75t_L g348 ( .A(n_15), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_135), .Y(n_349) );
INVxp67_ASAP7_75t_L g350 ( .A(n_46), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_306), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_54), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_119), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_95), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_50), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_326), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_99), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_293), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_272), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_32), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_134), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_214), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_137), .Y(n_363) );
CKINVDCx20_ASAP7_75t_R g364 ( .A(n_322), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_108), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_40), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_261), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_199), .Y(n_368) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_177), .Y(n_369) );
CKINVDCx16_ASAP7_75t_R g370 ( .A(n_88), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_328), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_28), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_173), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g374 ( .A(n_133), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_34), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_240), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_69), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_208), .Y(n_378) );
CKINVDCx16_ASAP7_75t_R g379 ( .A(n_109), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_342), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_110), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_337), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_317), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_198), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_282), .Y(n_385) );
INVx1_ASAP7_75t_SL g386 ( .A(n_329), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_193), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_21), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_225), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_38), .Y(n_390) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_78), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_139), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_229), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_18), .Y(n_394) );
INVxp67_ASAP7_75t_L g395 ( .A(n_178), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_259), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_167), .Y(n_397) );
CKINVDCx5p33_ASAP7_75t_R g398 ( .A(n_17), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_145), .Y(n_399) );
BUFx3_ASAP7_75t_L g400 ( .A(n_310), .Y(n_400) );
CKINVDCx5p33_ASAP7_75t_R g401 ( .A(n_151), .Y(n_401) );
CKINVDCx20_ASAP7_75t_R g402 ( .A(n_327), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_102), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_204), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_243), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_333), .Y(n_406) );
INVx1_ASAP7_75t_SL g407 ( .A(n_321), .Y(n_407) );
CKINVDCx5p33_ASAP7_75t_R g408 ( .A(n_44), .Y(n_408) );
BUFx3_ASAP7_75t_L g409 ( .A(n_247), .Y(n_409) );
NOR2xp67_ASAP7_75t_L g410 ( .A(n_252), .B(n_181), .Y(n_410) );
CKINVDCx5p33_ASAP7_75t_R g411 ( .A(n_280), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_324), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_55), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_65), .Y(n_414) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_315), .Y(n_415) );
CKINVDCx16_ASAP7_75t_R g416 ( .A(n_281), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_103), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_116), .Y(n_418) );
CKINVDCx20_ASAP7_75t_R g419 ( .A(n_210), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_114), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_15), .Y(n_421) );
INVx1_ASAP7_75t_SL g422 ( .A(n_74), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_279), .Y(n_423) );
INVxp67_ASAP7_75t_L g424 ( .A(n_62), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_331), .Y(n_425) );
INVxp67_ASAP7_75t_L g426 ( .A(n_227), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_98), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_262), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_148), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_169), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_97), .Y(n_431) );
CKINVDCx5p33_ASAP7_75t_R g432 ( .A(n_187), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_190), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_10), .Y(n_434) );
CKINVDCx5p33_ASAP7_75t_R g435 ( .A(n_335), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_66), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_311), .Y(n_437) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_213), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_233), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_87), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_312), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_56), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_138), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_96), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_107), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_336), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_129), .Y(n_447) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_292), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_46), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_325), .Y(n_450) );
CKINVDCx16_ASAP7_75t_R g451 ( .A(n_338), .Y(n_451) );
CKINVDCx5p33_ASAP7_75t_R g452 ( .A(n_343), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_117), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_283), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_286), .Y(n_455) );
BUFx5_ASAP7_75t_L g456 ( .A(n_23), .Y(n_456) );
BUFx3_ASAP7_75t_L g457 ( .A(n_298), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_150), .Y(n_458) );
INVxp33_ASAP7_75t_SL g459 ( .A(n_67), .Y(n_459) );
INVxp33_ASAP7_75t_L g460 ( .A(n_332), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_278), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_313), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_334), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_319), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_330), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_50), .Y(n_466) );
CKINVDCx16_ASAP7_75t_R g467 ( .A(n_236), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_308), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_16), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g470 ( .A(n_9), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_146), .Y(n_471) );
INVx1_ASAP7_75t_SL g472 ( .A(n_216), .Y(n_472) );
CKINVDCx5p33_ASAP7_75t_R g473 ( .A(n_288), .Y(n_473) );
CKINVDCx5p33_ASAP7_75t_R g474 ( .A(n_159), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g475 ( .A(n_182), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_2), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_185), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_235), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_277), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_239), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_260), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_52), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_77), .Y(n_483) );
CKINVDCx5p33_ASAP7_75t_R g484 ( .A(n_295), .Y(n_484) );
INVx2_ASAP7_75t_SL g485 ( .A(n_291), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_234), .Y(n_486) );
CKINVDCx5p33_ASAP7_75t_R g487 ( .A(n_323), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_44), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_13), .Y(n_489) );
CKINVDCx16_ASAP7_75t_R g490 ( .A(n_52), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_29), .Y(n_491) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_314), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_115), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g494 ( .A(n_194), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_320), .Y(n_495) );
INVxp67_ASAP7_75t_L g496 ( .A(n_12), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_456), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_456), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_353), .B(n_0), .Y(n_499) );
AND2x6_ASAP7_75t_L g500 ( .A(n_363), .B(n_57), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_456), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_353), .B(n_0), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_370), .Y(n_503) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_369), .Y(n_504) );
OAI22x1_ASAP7_75t_SL g505 ( .A1(n_388), .A2(n_3), .B1(n_1), .B2(n_2), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_415), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_456), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_415), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_456), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_485), .B(n_1), .Y(n_510) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_369), .Y(n_511) );
BUFx6f_ASAP7_75t_L g512 ( .A(n_369), .Y(n_512) );
AND2x4_ASAP7_75t_L g513 ( .A(n_394), .B(n_3), .Y(n_513) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_354), .A2(n_357), .B(n_356), .Y(n_514) );
INVx3_ASAP7_75t_L g515 ( .A(n_456), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_373), .Y(n_516) );
BUFx6f_ASAP7_75t_L g517 ( .A(n_391), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_437), .Y(n_518) );
BUFx12f_ASAP7_75t_L g519 ( .A(n_355), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_348), .B(n_4), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_349), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_379), .A2(n_6), .B1(n_4), .B2(n_5), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_515), .B(n_351), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_506), .B(n_416), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_513), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_513), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_508), .B(n_490), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_502), .Y(n_528) );
NAND3xp33_ASAP7_75t_L g529 ( .A(n_499), .B(n_496), .C(n_350), .Y(n_529) );
INVx2_ASAP7_75t_SL g530 ( .A(n_516), .Y(n_530) );
OAI22xp33_ASAP7_75t_L g531 ( .A1(n_522), .A2(n_489), .B1(n_496), .B2(n_350), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_515), .B(n_393), .Y(n_532) );
INVx4_ASAP7_75t_L g533 ( .A(n_500), .Y(n_533) );
AND2x2_ASAP7_75t_SL g534 ( .A(n_502), .B(n_451), .Y(n_534) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_504), .Y(n_535) );
NAND3xp33_ASAP7_75t_L g536 ( .A(n_499), .B(n_390), .C(n_360), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_497), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_510), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_510), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_518), .B(n_366), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_498), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_521), .B(n_467), .Y(n_542) );
INVx5_ASAP7_75t_L g543 ( .A(n_500), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_501), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_507), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_503), .B(n_460), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_538), .B(n_503), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_539), .B(n_528), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_537), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_542), .B(n_475), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_525), .A2(n_514), .B1(n_509), .B2(n_500), .Y(n_551) );
INVx3_ASAP7_75t_L g552 ( .A(n_533), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_530), .B(n_520), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_537), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_524), .B(n_514), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_526), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_540), .Y(n_557) );
AND2x4_ASAP7_75t_L g558 ( .A(n_536), .B(n_520), .Y(n_558) );
NOR3xp33_ASAP7_75t_L g559 ( .A(n_531), .B(n_408), .C(n_398), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_533), .A2(n_500), .B1(n_534), .B2(n_529), .Y(n_560) );
BUFx3_ASAP7_75t_L g561 ( .A(n_543), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_534), .B(n_546), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_546), .B(n_459), .Y(n_563) );
NOR2xp67_ASAP7_75t_L g564 ( .A(n_527), .B(n_519), .Y(n_564) );
BUFx2_ASAP7_75t_L g565 ( .A(n_531), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_523), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_541), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_523), .B(n_500), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_532), .B(n_395), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_532), .Y(n_570) );
NAND2x1_ASAP7_75t_L g571 ( .A(n_545), .B(n_361), .Y(n_571) );
CKINVDCx5p33_ASAP7_75t_R g572 ( .A(n_544), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_543), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_543), .A2(n_368), .B(n_365), .Y(n_574) );
NOR2xp33_ASAP7_75t_SL g575 ( .A(n_543), .B(n_362), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_535), .B(n_421), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_535), .B(n_395), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_535), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_535), .B(n_424), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_538), .B(n_424), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_538), .B(n_426), .Y(n_581) );
OAI22xp33_ASAP7_75t_L g582 ( .A1(n_528), .A2(n_374), .B1(n_402), .B2(n_364), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_538), .B(n_426), .Y(n_583) );
BUFx8_ASAP7_75t_L g584 ( .A(n_527), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_537), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_528), .Y(n_586) );
CKINVDCx5p33_ASAP7_75t_R g587 ( .A(n_534), .Y(n_587) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_568), .A2(n_376), .B(n_371), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_548), .B(n_352), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_586), .A2(n_455), .B1(n_477), .B2(n_419), .Y(n_590) );
O2A1O1Ixp33_ASAP7_75t_SL g591 ( .A1(n_555), .A2(n_381), .B(n_383), .C(n_377), .Y(n_591) );
INVx2_ASAP7_75t_SL g592 ( .A(n_584), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_562), .B(n_505), .Y(n_593) );
A2O1A1Ixp33_ASAP7_75t_L g594 ( .A1(n_553), .A2(n_375), .B(n_434), .C(n_372), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_553), .B(n_358), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_558), .B(n_470), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_558), .B(n_449), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_551), .A2(n_389), .B(n_384), .Y(n_598) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_584), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_560), .A2(n_469), .B1(n_476), .B2(n_466), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_557), .B(n_482), .Y(n_601) );
INVxp67_ASAP7_75t_SL g602 ( .A(n_582), .Y(n_602) );
BUFx4f_ASAP7_75t_L g603 ( .A(n_556), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_565), .B(n_488), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_559), .B(n_491), .Y(n_605) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_551), .A2(n_399), .B(n_392), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_549), .Y(n_607) );
O2A1O1Ixp5_ASAP7_75t_L g608 ( .A1(n_571), .A2(n_453), .B(n_458), .C(n_428), .Y(n_608) );
NAND2x1p5_ASAP7_75t_L g609 ( .A(n_561), .B(n_403), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_580), .B(n_359), .Y(n_610) );
O2A1O1Ixp33_ASAP7_75t_L g611 ( .A1(n_581), .A2(n_406), .B(n_413), .C(n_412), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_583), .B(n_367), .Y(n_612) );
AOI21xp5_ASAP7_75t_L g613 ( .A1(n_573), .A2(n_418), .B(n_417), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_547), .B(n_378), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_560), .A2(n_425), .B1(n_427), .B2(n_420), .Y(n_615) );
INVx2_ASAP7_75t_SL g616 ( .A(n_572), .Y(n_616) );
OAI22x1_ASAP7_75t_L g617 ( .A1(n_587), .A2(n_382), .B1(n_385), .B2(n_380), .Y(n_617) );
NOR3xp33_ASAP7_75t_L g618 ( .A(n_547), .B(n_407), .C(n_386), .Y(n_618) );
BUFx2_ASAP7_75t_L g619 ( .A(n_576), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_564), .A2(n_430), .B1(n_431), .B2(n_429), .Y(n_620) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_550), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_549), .Y(n_622) );
INVx1_ASAP7_75t_SL g623 ( .A(n_554), .Y(n_623) );
AND2x4_ASAP7_75t_L g624 ( .A(n_563), .B(n_433), .Y(n_624) );
O2A1O1Ixp33_ASAP7_75t_L g625 ( .A1(n_563), .A2(n_436), .B(n_440), .C(n_439), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g626 ( .A1(n_566), .A2(n_442), .B(n_441), .Y(n_626) );
INVx3_ASAP7_75t_SL g627 ( .A(n_570), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_569), .B(n_387), .Y(n_628) );
AOI33xp33_ASAP7_75t_L g629 ( .A1(n_567), .A2(n_447), .A3(n_444), .B1(n_454), .B2(n_450), .B3(n_446), .Y(n_629) );
BUFx2_ASAP7_75t_L g630 ( .A(n_585), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_569), .A2(n_461), .B1(n_465), .B2(n_464), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_554), .A2(n_471), .B(n_468), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_585), .Y(n_633) );
BUFx12f_ASAP7_75t_L g634 ( .A(n_575), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_567), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_552), .B(n_422), .Y(n_636) );
OAI21xp5_ASAP7_75t_L g637 ( .A1(n_574), .A2(n_480), .B(n_478), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_619), .Y(n_638) );
AOI21x1_ASAP7_75t_L g639 ( .A1(n_598), .A2(n_579), .B(n_577), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_621), .B(n_552), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_604), .B(n_486), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_594), .B(n_493), .Y(n_642) );
CKINVDCx8_ASAP7_75t_R g643 ( .A(n_624), .Y(n_643) );
OAI21x1_ASAP7_75t_L g644 ( .A1(n_606), .A2(n_578), .B(n_495), .Y(n_644) );
OAI21xp5_ASAP7_75t_L g645 ( .A1(n_588), .A2(n_561), .B(n_578), .Y(n_645) );
AOI21x1_ASAP7_75t_L g646 ( .A1(n_615), .A2(n_600), .B(n_632), .Y(n_646) );
BUFx6f_ASAP7_75t_L g647 ( .A(n_630), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_601), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_624), .B(n_396), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_597), .Y(n_650) );
NAND2x1p5_ASAP7_75t_L g651 ( .A(n_592), .B(n_472), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_602), .B(n_397), .Y(n_652) );
AO31x2_ASAP7_75t_L g653 ( .A1(n_600), .A2(n_631), .A3(n_607), .B(n_622), .Y(n_653) );
O2A1O1Ixp33_ASAP7_75t_L g654 ( .A1(n_625), .A2(n_479), .B(n_409), .C(n_457), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_629), .B(n_401), .Y(n_655) );
OAI21xp5_ASAP7_75t_L g656 ( .A1(n_608), .A2(n_410), .B(n_405), .Y(n_656) );
OA21x2_ASAP7_75t_L g657 ( .A1(n_637), .A2(n_411), .B(n_404), .Y(n_657) );
AOI21xp5_ASAP7_75t_SL g658 ( .A1(n_609), .A2(n_400), .B(n_391), .Y(n_658) );
CKINVDCx11_ASAP7_75t_R g659 ( .A(n_634), .Y(n_659) );
AND2x2_ASAP7_75t_SL g660 ( .A(n_603), .B(n_391), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_590), .A2(n_423), .B1(n_432), .B2(n_414), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_596), .Y(n_662) );
CKINVDCx11_ASAP7_75t_R g663 ( .A(n_627), .Y(n_663) );
INVxp67_ASAP7_75t_L g664 ( .A(n_590), .Y(n_664) );
BUFx2_ASAP7_75t_L g665 ( .A(n_616), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_605), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_635), .Y(n_667) );
AOI21xp5_ASAP7_75t_L g668 ( .A1(n_623), .A2(n_443), .B(n_435), .Y(n_668) );
BUFx4_ASAP7_75t_SL g669 ( .A(n_599), .Y(n_669) );
INVx4_ASAP7_75t_L g670 ( .A(n_603), .Y(n_670) );
AOI21xp5_ASAP7_75t_L g671 ( .A1(n_633), .A2(n_452), .B(n_445), .Y(n_671) );
AOI221xp5_ASAP7_75t_L g672 ( .A1(n_631), .A2(n_462), .B1(n_474), .B2(n_473), .C(n_463), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_609), .A2(n_483), .B1(n_484), .B2(n_481), .Y(n_673) );
OAI22xp33_ASAP7_75t_L g674 ( .A1(n_593), .A2(n_492), .B1(n_494), .B2(n_487), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_611), .Y(n_675) );
BUFx3_ASAP7_75t_L g676 ( .A(n_617), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g677 ( .A1(n_610), .A2(n_448), .B(n_438), .Y(n_677) );
AO31x2_ASAP7_75t_L g678 ( .A1(n_626), .A2(n_511), .A3(n_512), .B(n_504), .Y(n_678) );
INVxp67_ASAP7_75t_L g679 ( .A(n_589), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_614), .B(n_620), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_618), .B(n_5), .Y(n_681) );
OR2x2_ASAP7_75t_L g682 ( .A(n_612), .B(n_6), .Y(n_682) );
AO32x2_ASAP7_75t_L g683 ( .A1(n_591), .A2(n_504), .A3(n_517), .B1(n_512), .B2(n_511), .Y(n_683) );
OAI21xp5_ASAP7_75t_L g684 ( .A1(n_637), .A2(n_448), .B(n_438), .Y(n_684) );
OAI21x1_ASAP7_75t_L g685 ( .A1(n_613), .A2(n_448), .B(n_438), .Y(n_685) );
OAI21x1_ASAP7_75t_L g686 ( .A1(n_595), .A2(n_59), .B(n_58), .Y(n_686) );
AND2x2_ASAP7_75t_SL g687 ( .A(n_636), .B(n_7), .Y(n_687) );
BUFx3_ASAP7_75t_L g688 ( .A(n_628), .Y(n_688) );
AOI21x1_ASAP7_75t_L g689 ( .A1(n_598), .A2(n_511), .B(n_504), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_619), .Y(n_690) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_590), .Y(n_691) );
BUFx2_ASAP7_75t_L g692 ( .A(n_616), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_621), .B(n_7), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_590), .A2(n_512), .B1(n_517), .B2(n_511), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_684), .A2(n_517), .B(n_512), .Y(n_695) );
AND2x4_ASAP7_75t_L g696 ( .A(n_670), .B(n_8), .Y(n_696) );
OAI21x1_ASAP7_75t_L g697 ( .A1(n_689), .A2(n_517), .B(n_61), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_667), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_648), .B(n_8), .Y(n_699) );
OAI21x1_ASAP7_75t_L g700 ( .A1(n_644), .A2(n_63), .B(n_60), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_638), .Y(n_701) );
AND2x4_ASAP7_75t_L g702 ( .A(n_670), .B(n_10), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_653), .Y(n_703) );
CKINVDCx11_ASAP7_75t_R g704 ( .A(n_659), .Y(n_704) );
BUFx6f_ASAP7_75t_L g705 ( .A(n_647), .Y(n_705) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_647), .Y(n_706) );
OAI21x1_ASAP7_75t_L g707 ( .A1(n_639), .A2(n_68), .B(n_64), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_677), .A2(n_71), .B(n_70), .Y(n_708) );
INVx2_ASAP7_75t_SL g709 ( .A(n_669), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g710 ( .A1(n_645), .A2(n_73), .B(n_72), .Y(n_710) );
CKINVDCx6p67_ASAP7_75t_R g711 ( .A(n_665), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_690), .Y(n_712) );
OA21x2_ASAP7_75t_L g713 ( .A1(n_656), .A2(n_76), .B(n_75), .Y(n_713) );
OR2x6_ASAP7_75t_L g714 ( .A(n_651), .B(n_11), .Y(n_714) );
OA21x2_ASAP7_75t_L g715 ( .A1(n_685), .A2(n_80), .B(n_79), .Y(n_715) );
AND2x4_ASAP7_75t_L g716 ( .A(n_688), .B(n_11), .Y(n_716) );
OAI21xp5_ASAP7_75t_L g717 ( .A1(n_662), .A2(n_12), .B(n_13), .Y(n_717) );
A2O1A1Ixp33_ASAP7_75t_L g718 ( .A1(n_654), .A2(n_17), .B(n_14), .C(n_16), .Y(n_718) );
AND2x4_ASAP7_75t_L g719 ( .A(n_650), .B(n_14), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_666), .B(n_18), .Y(n_720) );
AOI21x1_ASAP7_75t_L g721 ( .A1(n_646), .A2(n_82), .B(n_81), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_653), .Y(n_722) );
BUFx4f_ASAP7_75t_SL g723 ( .A(n_692), .Y(n_723) );
NAND2xp5_ASAP7_75t_SL g724 ( .A(n_660), .B(n_19), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g725 ( .A1(n_675), .A2(n_84), .B(n_83), .Y(n_725) );
AO21x2_ASAP7_75t_L g726 ( .A1(n_642), .A2(n_86), .B(n_85), .Y(n_726) );
AND2x2_ASAP7_75t_L g727 ( .A(n_664), .B(n_19), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g728 ( .A1(n_657), .A2(n_90), .B(n_89), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_653), .Y(n_729) );
AO21x2_ASAP7_75t_L g730 ( .A1(n_686), .A2(n_694), .B(n_655), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_641), .B(n_20), .Y(n_731) );
OAI21x1_ASAP7_75t_L g732 ( .A1(n_658), .A2(n_92), .B(n_91), .Y(n_732) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_647), .Y(n_733) );
BUFx6f_ASAP7_75t_L g734 ( .A(n_683), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_693), .B(n_20), .Y(n_735) );
OA21x2_ASAP7_75t_L g736 ( .A1(n_681), .A2(n_94), .B(n_93), .Y(n_736) );
NOR2x1_ASAP7_75t_R g737 ( .A(n_676), .B(n_21), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_682), .Y(n_738) );
BUFx2_ASAP7_75t_L g739 ( .A(n_687), .Y(n_739) );
AOI21x1_ASAP7_75t_L g740 ( .A1(n_657), .A2(n_101), .B(n_100), .Y(n_740) );
OAI21x1_ASAP7_75t_L g741 ( .A1(n_668), .A2(n_105), .B(n_104), .Y(n_741) );
OAI21x1_ASAP7_75t_L g742 ( .A1(n_671), .A2(n_640), .B(n_683), .Y(n_742) );
AOI21xp5_ASAP7_75t_L g743 ( .A1(n_652), .A2(n_679), .B(n_649), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_678), .Y(n_744) );
AO31x2_ASAP7_75t_L g745 ( .A1(n_683), .A2(n_24), .A3(n_22), .B(n_23), .Y(n_745) );
OAI21x1_ASAP7_75t_L g746 ( .A1(n_673), .A2(n_111), .B(n_106), .Y(n_746) );
OA21x2_ASAP7_75t_L g747 ( .A1(n_678), .A2(n_113), .B(n_112), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_643), .Y(n_748) );
CKINVDCx16_ASAP7_75t_R g749 ( .A(n_661), .Y(n_749) );
AOI21xp5_ASAP7_75t_L g750 ( .A1(n_672), .A2(n_120), .B(n_118), .Y(n_750) );
CKINVDCx5p33_ASAP7_75t_R g751 ( .A(n_674), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_678), .A2(n_25), .B1(n_22), .B2(n_24), .Y(n_752) );
INVx2_ASAP7_75t_L g753 ( .A(n_667), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_648), .Y(n_754) );
OAI21x1_ASAP7_75t_L g755 ( .A1(n_689), .A2(n_122), .B(n_121), .Y(n_755) );
CKINVDCx6p67_ASAP7_75t_R g756 ( .A(n_663), .Y(n_756) );
OA21x2_ASAP7_75t_L g757 ( .A1(n_684), .A2(n_124), .B(n_123), .Y(n_757) );
OAI21xp5_ASAP7_75t_L g758 ( .A1(n_680), .A2(n_25), .B(n_26), .Y(n_758) );
OAI21x1_ASAP7_75t_L g759 ( .A1(n_689), .A2(n_126), .B(n_125), .Y(n_759) );
AND2x4_ASAP7_75t_L g760 ( .A(n_670), .B(n_26), .Y(n_760) );
AOI21xp5_ASAP7_75t_L g761 ( .A1(n_684), .A2(n_128), .B(n_127), .Y(n_761) );
AND2x2_ASAP7_75t_L g762 ( .A(n_691), .B(n_27), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_716), .B(n_27), .Y(n_763) );
AND2x2_ASAP7_75t_L g764 ( .A(n_716), .B(n_28), .Y(n_764) );
INVx2_ASAP7_75t_L g765 ( .A(n_698), .Y(n_765) );
INVx3_ASAP7_75t_L g766 ( .A(n_705), .Y(n_766) );
AND2x2_ASAP7_75t_L g767 ( .A(n_719), .B(n_29), .Y(n_767) );
INVx3_ASAP7_75t_L g768 ( .A(n_705), .Y(n_768) );
INVx2_ASAP7_75t_L g769 ( .A(n_753), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_754), .Y(n_770) );
BUFx2_ASAP7_75t_L g771 ( .A(n_723), .Y(n_771) );
INVx2_ASAP7_75t_SL g772 ( .A(n_709), .Y(n_772) );
INVx2_ASAP7_75t_L g773 ( .A(n_701), .Y(n_773) );
AND2x2_ASAP7_75t_L g774 ( .A(n_719), .B(n_30), .Y(n_774) );
AND2x2_ASAP7_75t_L g775 ( .A(n_739), .B(n_30), .Y(n_775) );
INVx2_ASAP7_75t_SL g776 ( .A(n_705), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_712), .Y(n_777) );
AND2x4_ASAP7_75t_L g778 ( .A(n_706), .B(n_31), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_749), .B(n_31), .Y(n_779) );
NOR2xp33_ASAP7_75t_SL g780 ( .A(n_756), .B(n_32), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_703), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_720), .Y(n_782) );
HB1xp67_ASAP7_75t_L g783 ( .A(n_722), .Y(n_783) );
AND2x2_ASAP7_75t_L g784 ( .A(n_714), .B(n_33), .Y(n_784) );
AO21x2_ASAP7_75t_L g785 ( .A1(n_744), .A2(n_33), .B(n_34), .Y(n_785) );
OR2x2_ASAP7_75t_L g786 ( .A(n_733), .B(n_35), .Y(n_786) );
BUFx3_ASAP7_75t_L g787 ( .A(n_711), .Y(n_787) );
BUFx2_ASAP7_75t_L g788 ( .A(n_748), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_729), .B(n_35), .Y(n_789) );
BUFx6f_ASAP7_75t_L g790 ( .A(n_734), .Y(n_790) );
OAI21x1_ASAP7_75t_SL g791 ( .A1(n_758), .A2(n_36), .B(n_37), .Y(n_791) );
INVx2_ASAP7_75t_L g792 ( .A(n_729), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_699), .Y(n_793) );
OR2x2_ASAP7_75t_L g794 ( .A(n_738), .B(n_36), .Y(n_794) );
AOI21x1_ASAP7_75t_L g795 ( .A1(n_721), .A2(n_740), .B(n_695), .Y(n_795) );
BUFx2_ASAP7_75t_L g796 ( .A(n_714), .Y(n_796) );
NAND2x1p5_ASAP7_75t_L g797 ( .A(n_696), .B(n_37), .Y(n_797) );
CKINVDCx14_ASAP7_75t_R g798 ( .A(n_704), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_696), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_762), .B(n_38), .Y(n_800) );
INVx2_ASAP7_75t_L g801 ( .A(n_745), .Y(n_801) );
AND2x2_ASAP7_75t_L g802 ( .A(n_727), .B(n_39), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_702), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_702), .Y(n_804) );
INVx2_ASAP7_75t_L g805 ( .A(n_734), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_760), .B(n_39), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_760), .Y(n_807) );
AND2x2_ASAP7_75t_L g808 ( .A(n_751), .B(n_40), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_717), .A2(n_43), .B1(n_41), .B2(n_42), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_730), .B(n_743), .Y(n_810) );
AND2x2_ASAP7_75t_L g811 ( .A(n_731), .B(n_41), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_735), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_745), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_745), .Y(n_814) );
AND2x2_ASAP7_75t_L g815 ( .A(n_724), .B(n_43), .Y(n_815) );
OR2x2_ASAP7_75t_L g816 ( .A(n_718), .B(n_45), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_752), .Y(n_817) );
AND2x4_ASAP7_75t_L g818 ( .A(n_732), .B(n_45), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_742), .B(n_47), .Y(n_819) );
BUFx3_ASAP7_75t_L g820 ( .A(n_746), .Y(n_820) );
AND2x2_ASAP7_75t_L g821 ( .A(n_736), .B(n_47), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_713), .B(n_48), .Y(n_822) );
INVx2_ASAP7_75t_L g823 ( .A(n_734), .Y(n_823) );
AO21x2_ASAP7_75t_L g824 ( .A1(n_707), .A2(n_728), .B(n_697), .Y(n_824) );
OR2x2_ASAP7_75t_L g825 ( .A(n_736), .B(n_48), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_737), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_747), .Y(n_827) );
INVx2_ASAP7_75t_L g828 ( .A(n_747), .Y(n_828) );
BUFx3_ASAP7_75t_L g829 ( .A(n_741), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_700), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_726), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_713), .A2(n_53), .B1(n_49), .B2(n_51), .Y(n_832) );
INVx2_ASAP7_75t_L g833 ( .A(n_715), .Y(n_833) );
AOI222xp33_ASAP7_75t_L g834 ( .A1(n_755), .A2(n_53), .B1(n_130), .B2(n_131), .C1(n_132), .C2(n_136), .Y(n_834) );
OA21x2_ASAP7_75t_L g835 ( .A1(n_759), .A2(n_140), .B(n_141), .Y(n_835) );
HB1xp67_ASAP7_75t_L g836 ( .A(n_757), .Y(n_836) );
AND2x2_ASAP7_75t_L g837 ( .A(n_757), .B(n_142), .Y(n_837) );
AO21x2_ASAP7_75t_L g838 ( .A1(n_710), .A2(n_143), .B(n_144), .Y(n_838) );
INVx2_ASAP7_75t_L g839 ( .A(n_715), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_750), .B(n_147), .Y(n_840) );
INVx2_ASAP7_75t_L g841 ( .A(n_761), .Y(n_841) );
BUFx2_ASAP7_75t_L g842 ( .A(n_708), .Y(n_842) );
AND2x2_ASAP7_75t_L g843 ( .A(n_725), .B(n_149), .Y(n_843) );
AOI221xp5_ASAP7_75t_L g844 ( .A1(n_739), .A2(n_152), .B1(n_153), .B2(n_154), .C(n_155), .Y(n_844) );
AO21x2_ASAP7_75t_L g845 ( .A1(n_744), .A2(n_156), .B(n_157), .Y(n_845) );
INVx2_ASAP7_75t_L g846 ( .A(n_703), .Y(n_846) );
INVx2_ASAP7_75t_L g847 ( .A(n_703), .Y(n_847) );
BUFx6f_ASAP7_75t_L g848 ( .A(n_705), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_754), .B(n_158), .Y(n_849) );
OA21x2_ASAP7_75t_L g850 ( .A1(n_744), .A2(n_160), .B(n_161), .Y(n_850) );
NOR2xp33_ASAP7_75t_L g851 ( .A(n_749), .B(n_162), .Y(n_851) );
AOI21xp5_ASAP7_75t_L g852 ( .A1(n_695), .A2(n_347), .B(n_163), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_754), .Y(n_853) );
INVx2_ASAP7_75t_L g854 ( .A(n_698), .Y(n_854) );
AOI21x1_ASAP7_75t_L g855 ( .A1(n_721), .A2(n_346), .B(n_164), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_754), .Y(n_856) );
INVx2_ASAP7_75t_L g857 ( .A(n_703), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_777), .Y(n_858) );
AND2x4_ASAP7_75t_L g859 ( .A(n_766), .B(n_165), .Y(n_859) );
INVx2_ASAP7_75t_L g860 ( .A(n_765), .Y(n_860) );
NOR2x1_ASAP7_75t_L g861 ( .A(n_796), .B(n_166), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_817), .B(n_168), .Y(n_862) );
BUFx2_ASAP7_75t_L g863 ( .A(n_787), .Y(n_863) );
INVx2_ASAP7_75t_L g864 ( .A(n_769), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_770), .Y(n_865) );
INVx2_ASAP7_75t_L g866 ( .A(n_854), .Y(n_866) );
AND2x2_ASAP7_75t_L g867 ( .A(n_806), .B(n_763), .Y(n_867) );
AND2x2_ASAP7_75t_L g868 ( .A(n_764), .B(n_170), .Y(n_868) );
OR2x2_ASAP7_75t_L g869 ( .A(n_773), .B(n_171), .Y(n_869) );
AND2x2_ASAP7_75t_L g870 ( .A(n_767), .B(n_172), .Y(n_870) );
AND2x4_ASAP7_75t_L g871 ( .A(n_766), .B(n_174), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_853), .Y(n_872) );
AND2x2_ASAP7_75t_L g873 ( .A(n_774), .B(n_175), .Y(n_873) );
AOI22xp5_ASAP7_75t_L g874 ( .A1(n_779), .A2(n_176), .B1(n_179), .B2(n_180), .Y(n_874) );
BUFx6f_ASAP7_75t_L g875 ( .A(n_848), .Y(n_875) );
INVxp67_ASAP7_75t_SL g876 ( .A(n_783), .Y(n_876) );
INVx2_ASAP7_75t_L g877 ( .A(n_856), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_789), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_789), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_794), .Y(n_880) );
AND2x2_ASAP7_75t_L g881 ( .A(n_808), .B(n_183), .Y(n_881) );
INVx3_ASAP7_75t_L g882 ( .A(n_848), .Y(n_882) );
AND2x2_ASAP7_75t_L g883 ( .A(n_775), .B(n_184), .Y(n_883) );
HB1xp67_ASAP7_75t_L g884 ( .A(n_781), .Y(n_884) );
OR2x2_ASAP7_75t_L g885 ( .A(n_786), .B(n_186), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_792), .B(n_188), .Y(n_886) );
AND2x2_ASAP7_75t_L g887 ( .A(n_784), .B(n_189), .Y(n_887) );
OR2x2_ASAP7_75t_L g888 ( .A(n_800), .B(n_345), .Y(n_888) );
INVx4_ASAP7_75t_L g889 ( .A(n_771), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_802), .B(n_191), .Y(n_890) );
HB1xp67_ASAP7_75t_L g891 ( .A(n_781), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_799), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_803), .Y(n_893) );
AND2x2_ASAP7_75t_L g894 ( .A(n_778), .B(n_192), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_804), .Y(n_895) );
HB1xp67_ASAP7_75t_L g896 ( .A(n_846), .Y(n_896) );
INVx3_ASAP7_75t_L g897 ( .A(n_848), .Y(n_897) );
AND2x2_ASAP7_75t_L g898 ( .A(n_797), .B(n_195), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_779), .A2(n_196), .B1(n_197), .B2(n_200), .Y(n_899) );
AND2x2_ASAP7_75t_L g900 ( .A(n_797), .B(n_201), .Y(n_900) );
INVx3_ASAP7_75t_L g901 ( .A(n_848), .Y(n_901) );
HB1xp67_ASAP7_75t_L g902 ( .A(n_846), .Y(n_902) );
INVx2_ASAP7_75t_L g903 ( .A(n_792), .Y(n_903) );
OR2x2_ASAP7_75t_L g904 ( .A(n_800), .B(n_202), .Y(n_904) );
AND2x2_ASAP7_75t_L g905 ( .A(n_811), .B(n_203), .Y(n_905) );
AND2x2_ASAP7_75t_L g906 ( .A(n_851), .B(n_205), .Y(n_906) );
OR2x2_ASAP7_75t_L g907 ( .A(n_807), .B(n_344), .Y(n_907) );
INVx2_ASAP7_75t_L g908 ( .A(n_847), .Y(n_908) );
AND2x2_ASAP7_75t_L g909 ( .A(n_851), .B(n_206), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_793), .B(n_207), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_785), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_812), .B(n_209), .Y(n_912) );
INVx2_ASAP7_75t_L g913 ( .A(n_847), .Y(n_913) );
AND2x4_ASAP7_75t_L g914 ( .A(n_768), .B(n_211), .Y(n_914) );
INVx1_ASAP7_75t_SL g915 ( .A(n_768), .Y(n_915) );
INVx2_ASAP7_75t_L g916 ( .A(n_857), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g917 ( .A(n_782), .B(n_212), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_785), .Y(n_918) );
INVx2_ASAP7_75t_SL g919 ( .A(n_787), .Y(n_919) );
OR2x2_ASAP7_75t_L g920 ( .A(n_776), .B(n_341), .Y(n_920) );
AND2x4_ASAP7_75t_SL g921 ( .A(n_772), .B(n_215), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_849), .Y(n_922) );
AND2x2_ASAP7_75t_L g923 ( .A(n_815), .B(n_217), .Y(n_923) );
BUFx4f_ASAP7_75t_L g924 ( .A(n_826), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_849), .Y(n_925) );
INVx2_ASAP7_75t_SL g926 ( .A(n_788), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_819), .Y(n_927) );
NOR2xp33_ASAP7_75t_L g928 ( .A(n_816), .B(n_218), .Y(n_928) );
AO21x2_ASAP7_75t_L g929 ( .A1(n_819), .A2(n_219), .B(n_220), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_818), .Y(n_930) );
NOR2x1_ASAP7_75t_R g931 ( .A(n_798), .B(n_221), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_818), .Y(n_932) );
INVx2_ASAP7_75t_L g933 ( .A(n_825), .Y(n_933) );
AO21x2_ASAP7_75t_L g934 ( .A1(n_795), .A2(n_222), .B(n_223), .Y(n_934) );
AND2x2_ASAP7_75t_L g935 ( .A(n_780), .B(n_809), .Y(n_935) );
HB1xp67_ASAP7_75t_L g936 ( .A(n_805), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_791), .Y(n_937) );
INVx2_ASAP7_75t_L g938 ( .A(n_813), .Y(n_938) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_814), .B(n_224), .Y(n_939) );
HB1xp67_ASAP7_75t_L g940 ( .A(n_823), .Y(n_940) );
HB1xp67_ASAP7_75t_L g941 ( .A(n_823), .Y(n_941) );
OR2x2_ASAP7_75t_L g942 ( .A(n_809), .B(n_340), .Y(n_942) );
AND2x2_ASAP7_75t_L g943 ( .A(n_821), .B(n_226), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_822), .Y(n_944) );
AND2x2_ASAP7_75t_L g945 ( .A(n_832), .B(n_228), .Y(n_945) );
AND2x2_ASAP7_75t_L g946 ( .A(n_832), .B(n_230), .Y(n_946) );
AND2x2_ASAP7_75t_L g947 ( .A(n_844), .B(n_231), .Y(n_947) );
BUFx2_ASAP7_75t_L g948 ( .A(n_798), .Y(n_948) );
INVx2_ASAP7_75t_L g949 ( .A(n_801), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_844), .B(n_232), .Y(n_950) );
AND2x2_ASAP7_75t_L g951 ( .A(n_834), .B(n_237), .Y(n_951) );
BUFx2_ASAP7_75t_L g952 ( .A(n_845), .Y(n_952) );
AND2x2_ASAP7_75t_L g953 ( .A(n_822), .B(n_238), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_810), .B(n_842), .Y(n_954) );
HB1xp67_ASAP7_75t_L g955 ( .A(n_790), .Y(n_955) );
INVx2_ASAP7_75t_L g956 ( .A(n_790), .Y(n_956) );
AND2x2_ASAP7_75t_L g957 ( .A(n_843), .B(n_241), .Y(n_957) );
INVx1_ASAP7_75t_L g958 ( .A(n_810), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_845), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_830), .Y(n_960) );
INVx2_ASAP7_75t_L g961 ( .A(n_790), .Y(n_961) );
OR2x2_ASAP7_75t_L g962 ( .A(n_790), .B(n_339), .Y(n_962) );
INVx1_ASAP7_75t_L g963 ( .A(n_850), .Y(n_963) );
BUFx2_ASAP7_75t_L g964 ( .A(n_820), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_820), .B(n_242), .Y(n_965) );
BUFx6f_ASAP7_75t_L g966 ( .A(n_829), .Y(n_966) );
NAND2xp5_ASAP7_75t_L g967 ( .A(n_831), .B(n_244), .Y(n_967) );
AND2x2_ASAP7_75t_L g968 ( .A(n_837), .B(n_245), .Y(n_968) );
HB1xp67_ASAP7_75t_L g969 ( .A(n_833), .Y(n_969) );
INVx3_ASAP7_75t_L g970 ( .A(n_850), .Y(n_970) );
HB1xp67_ASAP7_75t_L g971 ( .A(n_833), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_838), .B(n_246), .Y(n_972) );
AND2x2_ASAP7_75t_L g973 ( .A(n_838), .B(n_248), .Y(n_973) );
INVx2_ASAP7_75t_SL g974 ( .A(n_829), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_858), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_867), .B(n_836), .Y(n_976) );
NAND2xp5_ASAP7_75t_L g977 ( .A(n_878), .B(n_836), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_865), .Y(n_978) );
INVx2_ASAP7_75t_L g979 ( .A(n_860), .Y(n_979) );
AND2x2_ASAP7_75t_L g980 ( .A(n_877), .B(n_827), .Y(n_980) );
AND2x4_ASAP7_75t_L g981 ( .A(n_930), .B(n_827), .Y(n_981) );
INVxp67_ASAP7_75t_SL g982 ( .A(n_884), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_872), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_880), .B(n_828), .Y(n_984) );
AOI33xp33_ASAP7_75t_L g985 ( .A1(n_935), .A2(n_839), .A3(n_841), .B1(n_250), .B2(n_251), .B3(n_253), .Y(n_985) );
AND2x2_ASAP7_75t_L g986 ( .A(n_864), .B(n_841), .Y(n_986) );
INVx2_ASAP7_75t_L g987 ( .A(n_866), .Y(n_987) );
AND2x2_ASAP7_75t_L g988 ( .A(n_932), .B(n_824), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_892), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_893), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g991 ( .A(n_879), .B(n_824), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_895), .Y(n_992) );
INVx2_ASAP7_75t_L g993 ( .A(n_884), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_876), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_889), .B(n_835), .Y(n_995) );
INVx2_ASAP7_75t_L g996 ( .A(n_891), .Y(n_996) );
AND2x2_ASAP7_75t_L g997 ( .A(n_889), .B(n_835), .Y(n_997) );
INVxp67_ASAP7_75t_L g998 ( .A(n_876), .Y(n_998) );
INVx2_ASAP7_75t_L g999 ( .A(n_891), .Y(n_999) );
HB1xp67_ASAP7_75t_L g1000 ( .A(n_896), .Y(n_1000) );
INVx2_ASAP7_75t_L g1001 ( .A(n_896), .Y(n_1001) );
NAND2x1p5_ASAP7_75t_L g1002 ( .A(n_863), .B(n_835), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_926), .B(n_840), .Y(n_1003) );
AND2x2_ASAP7_75t_SL g1004 ( .A(n_964), .B(n_852), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_903), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_902), .Y(n_1006) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_927), .B(n_852), .Y(n_1007) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_944), .B(n_855), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_938), .Y(n_1009) );
AND2x2_ASAP7_75t_L g1010 ( .A(n_933), .B(n_249), .Y(n_1010) );
INVx2_ASAP7_75t_L g1011 ( .A(n_908), .Y(n_1011) );
INVx1_ASAP7_75t_L g1012 ( .A(n_913), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_916), .Y(n_1013) );
NAND2xp5_ASAP7_75t_SL g1014 ( .A(n_974), .B(n_254), .Y(n_1014) );
AND2x2_ASAP7_75t_L g1015 ( .A(n_887), .B(n_255), .Y(n_1015) );
INVx1_ASAP7_75t_L g1016 ( .A(n_960), .Y(n_1016) );
NOR2xp33_ASAP7_75t_L g1017 ( .A(n_888), .B(n_256), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_881), .B(n_257), .Y(n_1018) );
NOR2xp67_ASAP7_75t_L g1019 ( .A(n_919), .B(n_258), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_915), .B(n_263), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_911), .Y(n_1021) );
AND2x2_ASAP7_75t_L g1022 ( .A(n_915), .B(n_264), .Y(n_1022) );
HB1xp67_ASAP7_75t_L g1023 ( .A(n_936), .Y(n_1023) );
OR2x2_ASAP7_75t_L g1024 ( .A(n_954), .B(n_265), .Y(n_1024) );
INVx2_ASAP7_75t_SL g1025 ( .A(n_948), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_918), .Y(n_1026) );
BUFx2_ASAP7_75t_L g1027 ( .A(n_882), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_868), .B(n_266), .Y(n_1028) );
INVx1_ASAP7_75t_SL g1029 ( .A(n_955), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_958), .Y(n_1030) );
OR2x2_ASAP7_75t_L g1031 ( .A(n_954), .B(n_267), .Y(n_1031) );
AND2x4_ASAP7_75t_L g1032 ( .A(n_955), .B(n_268), .Y(n_1032) );
AND2x4_ASAP7_75t_L g1033 ( .A(n_936), .B(n_269), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_870), .B(n_270), .Y(n_1034) );
INVx1_ASAP7_75t_L g1035 ( .A(n_886), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_873), .B(n_271), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_886), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_890), .B(n_273), .Y(n_1038) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_937), .B(n_274), .Y(n_1039) );
INVx1_ASAP7_75t_L g1040 ( .A(n_922), .Y(n_1040) );
NAND3xp33_ASAP7_75t_L g1041 ( .A(n_874), .B(n_275), .C(n_276), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_925), .Y(n_1042) );
NAND2x1_ASAP7_75t_L g1043 ( .A(n_861), .B(n_284), .Y(n_1043) );
INVx4_ASAP7_75t_L g1044 ( .A(n_859), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_940), .B(n_285), .Y(n_1045) );
AND2x4_ASAP7_75t_SL g1046 ( .A(n_859), .B(n_287), .Y(n_1046) );
INVxp67_ASAP7_75t_SL g1047 ( .A(n_969), .Y(n_1047) );
NAND2xp5_ASAP7_75t_L g1048 ( .A(n_940), .B(n_289), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_939), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_939), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g1051 ( .A(n_941), .B(n_290), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1052 ( .A(n_883), .B(n_294), .Y(n_1052) );
AND2x2_ASAP7_75t_SL g1053 ( .A(n_921), .B(n_296), .Y(n_1053) );
INVx1_ASAP7_75t_L g1054 ( .A(n_967), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_941), .B(n_297), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_943), .B(n_299), .Y(n_1056) );
INVx2_ASAP7_75t_L g1057 ( .A(n_969), .Y(n_1057) );
INVx1_ASAP7_75t_L g1058 ( .A(n_967), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g1059 ( .A1(n_951), .A2(n_300), .B1(n_301), .B2(n_302), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g1060 ( .A(n_949), .B(n_303), .Y(n_1060) );
AND2x2_ASAP7_75t_L g1061 ( .A(n_894), .B(n_304), .Y(n_1061) );
INVx2_ASAP7_75t_L g1062 ( .A(n_971), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_953), .B(n_305), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_869), .Y(n_1064) );
INVx2_ASAP7_75t_L g1065 ( .A(n_882), .Y(n_1065) );
AND2x2_ASAP7_75t_L g1066 ( .A(n_976), .B(n_956), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_975), .B(n_978), .Y(n_1067) );
OR2x2_ASAP7_75t_L g1068 ( .A(n_1000), .B(n_961), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_983), .B(n_897), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_1030), .B(n_959), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_984), .B(n_897), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_1040), .B(n_952), .Y(n_1072) );
INVx2_ASAP7_75t_SL g1073 ( .A(n_1025), .Y(n_1073) );
OR2x2_ASAP7_75t_SL g1074 ( .A(n_1041), .B(n_931), .Y(n_1074) );
NAND2xp5_ASAP7_75t_L g1075 ( .A(n_1042), .B(n_963), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1003), .B(n_901), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_989), .B(n_901), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g1078 ( .A(n_990), .B(n_928), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_992), .B(n_966), .Y(n_1079) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1016), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_979), .B(n_966), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_987), .B(n_924), .Y(n_1082) );
HB1xp67_ASAP7_75t_L g1083 ( .A(n_1023), .Y(n_1083) );
OR2x2_ASAP7_75t_L g1084 ( .A(n_1000), .B(n_965), .Y(n_1084) );
NAND2xp5_ASAP7_75t_L g1085 ( .A(n_977), .B(n_970), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_977), .B(n_970), .Y(n_1086) );
AND2x2_ASAP7_75t_L g1087 ( .A(n_1029), .B(n_898), .Y(n_1087) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_994), .B(n_965), .Y(n_1088) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1009), .Y(n_1089) );
AND2x4_ASAP7_75t_L g1090 ( .A(n_988), .B(n_875), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_1027), .B(n_900), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1006), .Y(n_1092) );
INVx2_ASAP7_75t_L g1093 ( .A(n_1057), .Y(n_1093) );
NOR2xp67_ASAP7_75t_L g1094 ( .A(n_1044), .B(n_874), .Y(n_1094) );
INVx2_ASAP7_75t_L g1095 ( .A(n_1062), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1096 ( .A(n_1023), .B(n_923), .Y(n_1096) );
NOR2xp33_ASAP7_75t_L g1097 ( .A(n_1053), .B(n_906), .Y(n_1097) );
NAND2xp5_ASAP7_75t_L g1098 ( .A(n_991), .B(n_928), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_998), .B(n_968), .Y(n_1099) );
OAI211xp5_ASAP7_75t_SL g1100 ( .A1(n_1059), .A2(n_899), .B(n_904), .C(n_912), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_998), .B(n_875), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_1005), .B(n_905), .Y(n_1102) );
CKINVDCx16_ASAP7_75t_R g1103 ( .A(n_1015), .Y(n_1103) );
NAND2xp5_ASAP7_75t_L g1104 ( .A(n_1054), .B(n_862), .Y(n_1104) );
INVx2_ASAP7_75t_SL g1105 ( .A(n_1053), .Y(n_1105) );
INVx1_ASAP7_75t_SL g1106 ( .A(n_993), .Y(n_1106) );
INVx1_ASAP7_75t_L g1107 ( .A(n_982), .Y(n_1107) );
OR2x2_ASAP7_75t_L g1108 ( .A(n_982), .B(n_885), .Y(n_1108) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_991), .B(n_945), .Y(n_1109) );
INVxp67_ASAP7_75t_SL g1110 ( .A(n_1047), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1012), .Y(n_1111) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1013), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_996), .B(n_972), .Y(n_1113) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_1021), .B(n_946), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1047), .Y(n_1115) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_1026), .B(n_973), .Y(n_1116) );
INVx1_ASAP7_75t_SL g1117 ( .A(n_999), .Y(n_1117) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1001), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_980), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_1058), .B(n_862), .Y(n_1120) );
AND2x4_ASAP7_75t_L g1121 ( .A(n_981), .B(n_921), .Y(n_1121) );
AND2x4_ASAP7_75t_L g1122 ( .A(n_1079), .B(n_981), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1080), .Y(n_1123) );
NAND4xp25_ASAP7_75t_L g1124 ( .A(n_1094), .B(n_1059), .C(n_899), .D(n_1017), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1067), .Y(n_1125) );
AND2x4_ASAP7_75t_L g1126 ( .A(n_1101), .B(n_1090), .Y(n_1126) );
INVxp67_ASAP7_75t_L g1127 ( .A(n_1073), .Y(n_1127) );
NAND2x1p5_ASAP7_75t_L g1128 ( .A(n_1121), .B(n_1019), .Y(n_1128) );
HB1xp67_ASAP7_75t_L g1129 ( .A(n_1083), .Y(n_1129) );
NOR2xp33_ASAP7_75t_L g1130 ( .A(n_1103), .B(n_1064), .Y(n_1130) );
OR4x1_ASAP7_75t_L g1131 ( .A(n_1105), .B(n_1043), .C(n_1050), .D(n_1049), .Y(n_1131) );
NOR2xp33_ASAP7_75t_L g1132 ( .A(n_1097), .B(n_909), .Y(n_1132) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1089), .Y(n_1133) );
AND2x2_ASAP7_75t_L g1134 ( .A(n_1076), .B(n_995), .Y(n_1134) );
INVx1_ASAP7_75t_SL g1135 ( .A(n_1066), .Y(n_1135) );
INVxp67_ASAP7_75t_SL g1136 ( .A(n_1110), .Y(n_1136) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1092), .Y(n_1137) );
INVx2_ASAP7_75t_L g1138 ( .A(n_1068), .Y(n_1138) );
OAI21xp33_ASAP7_75t_SL g1139 ( .A1(n_1091), .A2(n_1004), .B(n_997), .Y(n_1139) );
NAND2xp5_ASAP7_75t_SL g1140 ( .A(n_1082), .B(n_1004), .Y(n_1140) );
NAND2xp5_ASAP7_75t_L g1141 ( .A(n_1119), .B(n_1098), .Y(n_1141) );
HB1xp67_ASAP7_75t_L g1142 ( .A(n_1106), .Y(n_1142) );
NAND3xp33_ASAP7_75t_L g1143 ( .A(n_1107), .B(n_985), .C(n_1007), .Y(n_1143) );
AOI32xp33_ASAP7_75t_L g1144 ( .A1(n_1100), .A2(n_1046), .A3(n_947), .B1(n_950), .B2(n_1017), .Y(n_1144) );
CKINVDCx20_ASAP7_75t_R g1145 ( .A(n_1071), .Y(n_1145) );
INVxp67_ASAP7_75t_SL g1146 ( .A(n_1115), .Y(n_1146) );
NAND2x1_ASAP7_75t_L g1147 ( .A(n_1111), .B(n_1033), .Y(n_1147) );
NAND2xp5_ASAP7_75t_L g1148 ( .A(n_1098), .B(n_1035), .Y(n_1148) );
BUFx2_ASAP7_75t_L g1149 ( .A(n_1117), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1150 ( .A(n_1087), .B(n_1011), .Y(n_1150) );
NAND4xp25_ASAP7_75t_L g1151 ( .A(n_1078), .B(n_985), .C(n_1018), .D(n_1061), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1152 ( .A(n_1126), .B(n_1096), .Y(n_1152) );
INVx3_ASAP7_75t_SL g1153 ( .A(n_1145), .Y(n_1153) );
INVx5_ASAP7_75t_L g1154 ( .A(n_1149), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1129), .Y(n_1155) );
AOI22xp33_ASAP7_75t_L g1156 ( .A1(n_1124), .A2(n_1099), .B1(n_1109), .B2(n_1116), .Y(n_1156) );
AOI221xp5_ASAP7_75t_L g1157 ( .A1(n_1139), .A2(n_1144), .B1(n_1148), .B2(n_1141), .C(n_1130), .Y(n_1157) );
INVx2_ASAP7_75t_L g1158 ( .A(n_1142), .Y(n_1158) );
OR2x2_ASAP7_75t_L g1159 ( .A(n_1135), .B(n_1085), .Y(n_1159) );
NOR2xp33_ASAP7_75t_L g1160 ( .A(n_1127), .B(n_1074), .Y(n_1160) );
AND2x2_ASAP7_75t_SL g1161 ( .A(n_1122), .B(n_1108), .Y(n_1161) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1146), .Y(n_1162) );
OAI21xp5_ASAP7_75t_L g1163 ( .A1(n_1136), .A2(n_1014), .B(n_1033), .Y(n_1163) );
AOI33xp33_ASAP7_75t_L g1164 ( .A1(n_1125), .A2(n_1102), .A3(n_1069), .B1(n_1077), .B2(n_1112), .B3(n_1113), .Y(n_1164) );
O2A1O1Ixp33_ASAP7_75t_L g1165 ( .A1(n_1140), .A2(n_1120), .B(n_1104), .C(n_1088), .Y(n_1165) );
OAI22xp33_ASAP7_75t_L g1166 ( .A1(n_1147), .A2(n_1084), .B1(n_1114), .B2(n_1109), .Y(n_1166) );
A2O1A1Ixp33_ASAP7_75t_L g1167 ( .A1(n_1144), .A2(n_1038), .B(n_1034), .C(n_1028), .Y(n_1167) );
OR2x2_ASAP7_75t_L g1168 ( .A(n_1138), .B(n_1085), .Y(n_1168) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1123), .Y(n_1169) );
AOI21xp33_ASAP7_75t_L g1170 ( .A1(n_1143), .A2(n_1120), .B(n_1024), .Y(n_1170) );
OAI31xp33_ASAP7_75t_L g1171 ( .A1(n_1167), .A2(n_1151), .A3(n_1128), .B(n_1132), .Y(n_1171) );
NAND2xp5_ASAP7_75t_L g1172 ( .A(n_1156), .B(n_1133), .Y(n_1172) );
AOI21xp5_ASAP7_75t_L g1173 ( .A1(n_1157), .A2(n_1072), .B(n_1086), .Y(n_1173) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1162), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1161), .B(n_1134), .Y(n_1175) );
AOI21xp33_ASAP7_75t_L g1176 ( .A1(n_1160), .A2(n_1072), .B(n_1137), .Y(n_1176) );
XNOR2x1_ASAP7_75t_L g1177 ( .A(n_1152), .B(n_1150), .Y(n_1177) );
AOI22xp5_ASAP7_75t_L g1178 ( .A1(n_1166), .A2(n_1114), .B1(n_1090), .B2(n_1118), .Y(n_1178) );
AOI21xp5_ASAP7_75t_R g1179 ( .A1(n_1153), .A2(n_1131), .B(n_1032), .Y(n_1179) );
OAI21xp5_ASAP7_75t_SL g1180 ( .A1(n_1163), .A2(n_1052), .B(n_1036), .Y(n_1180) );
OAI21xp5_ASAP7_75t_L g1181 ( .A1(n_1163), .A2(n_1088), .B(n_1056), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1169), .Y(n_1182) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1165), .B(n_1093), .Y(n_1183) );
OAI22xp5_ASAP7_75t_L g1184 ( .A1(n_1154), .A2(n_1031), .B1(n_1002), .B2(n_1095), .Y(n_1184) );
AOI221xp5_ASAP7_75t_L g1185 ( .A1(n_1170), .A2(n_1070), .B1(n_1075), .B2(n_1037), .C(n_1007), .Y(n_1185) );
NOR3xp33_ASAP7_75t_L g1186 ( .A(n_1170), .B(n_1063), .C(n_1039), .Y(n_1186) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1159), .Y(n_1187) );
NOR2xp33_ASAP7_75t_L g1188 ( .A(n_1155), .B(n_1075), .Y(n_1188) );
AOI221xp5_ASAP7_75t_L g1189 ( .A1(n_1158), .A2(n_912), .B1(n_917), .B2(n_910), .C(n_1081), .Y(n_1189) );
OAI22xp33_ASAP7_75t_L g1190 ( .A1(n_1154), .A2(n_1002), .B1(n_1048), .B2(n_1045), .Y(n_1190) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1164), .B(n_986), .Y(n_1191) );
AOI311xp33_ASAP7_75t_L g1192 ( .A1(n_1168), .A2(n_1008), .A3(n_1051), .B(n_1060), .C(n_942), .Y(n_1192) );
NOR2xp33_ASAP7_75t_L g1193 ( .A(n_1172), .B(n_1176), .Y(n_1193) );
NOR2xp33_ASAP7_75t_L g1194 ( .A(n_1183), .B(n_1191), .Y(n_1194) );
NAND2xp5_ASAP7_75t_L g1195 ( .A(n_1173), .B(n_1185), .Y(n_1195) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1182), .Y(n_1196) );
NOR2xp33_ASAP7_75t_L g1197 ( .A(n_1174), .B(n_1187), .Y(n_1197) );
OAI221xp5_ASAP7_75t_L g1198 ( .A1(n_1171), .A2(n_1180), .B1(n_1181), .B2(n_1192), .C(n_1178), .Y(n_1198) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1194), .B(n_1188), .Y(n_1199) );
NAND3xp33_ASAP7_75t_SL g1200 ( .A(n_1198), .B(n_1179), .C(n_1186), .Y(n_1200) );
NOR3xp33_ASAP7_75t_L g1201 ( .A(n_1195), .B(n_1189), .C(n_1190), .Y(n_1201) );
INVxp67_ASAP7_75t_SL g1202 ( .A(n_1197), .Y(n_1202) );
NOR2xp33_ASAP7_75t_L g1203 ( .A(n_1200), .B(n_1193), .Y(n_1203) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1202), .Y(n_1204) );
NAND4xp75_ASAP7_75t_L g1205 ( .A(n_1199), .B(n_1196), .C(n_1175), .D(n_957), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1204), .Y(n_1206) );
AOI22x1_ASAP7_75t_L g1207 ( .A1(n_1203), .A2(n_1201), .B1(n_871), .B2(n_914), .Y(n_1207) );
OAI22xp5_ASAP7_75t_L g1208 ( .A1(n_1207), .A2(n_1205), .B1(n_1177), .B2(n_1184), .Y(n_1208) );
AND5x1_ASAP7_75t_L g1209 ( .A(n_1206), .B(n_1010), .C(n_1022), .D(n_1020), .E(n_1055), .Y(n_1209) );
OAI22xp5_ASAP7_75t_L g1210 ( .A1(n_1208), .A2(n_907), .B1(n_1065), .B2(n_1008), .Y(n_1210) );
OAI22xp5_ASAP7_75t_SL g1211 ( .A1(n_1210), .A2(n_1209), .B1(n_920), .B2(n_962), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1212 ( .A(n_1211), .B(n_929), .Y(n_1212) );
OAI21xp33_ASAP7_75t_L g1213 ( .A1(n_1212), .A2(n_307), .B(n_309), .Y(n_1213) );
AOI22xp5_ASAP7_75t_L g1214 ( .A1(n_1213), .A2(n_934), .B1(n_316), .B2(n_318), .Y(n_1214) );
endmodule