module real_aes_7523_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_721, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_721;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_449;
wire n_182;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g175 ( .A1(n_0), .A2(n_176), .B(n_177), .C(n_181), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_1), .B(n_170), .Y(n_183) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_2), .B(n_93), .C(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g427 ( .A(n_2), .Y(n_427) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_3), .B(n_155), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_4), .A2(n_144), .B(n_161), .C(n_469), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_5), .A2(n_164), .B(n_490), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_6), .A2(n_164), .B(n_266), .Y(n_265) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_7), .A2(n_38), .B1(n_123), .B2(n_124), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_7), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_7), .B(n_170), .Y(n_496) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_8), .A2(n_136), .B(n_223), .Y(n_222) );
AND2x6_ASAP7_75t_L g161 ( .A(n_9), .B(n_162), .Y(n_161) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_10), .A2(n_144), .B(n_161), .C(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g461 ( .A(n_11), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_12), .B(n_43), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_13), .B(n_180), .Y(n_471) );
INVx1_ASAP7_75t_L g141 ( .A(n_14), .Y(n_141) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_15), .A2(n_105), .B1(n_114), .B2(n_719), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_16), .B(n_155), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g428 ( .A(n_17), .B(n_429), .Y(n_428) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_18), .A2(n_156), .B(n_480), .C(n_482), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_19), .B(n_170), .Y(n_483) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_20), .A2(n_68), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_20), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_21), .B(n_213), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_22), .A2(n_144), .B(n_207), .C(n_212), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g450 ( .A1(n_23), .A2(n_179), .B(n_231), .C(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_24), .B(n_180), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_25), .B(n_180), .Y(n_512) );
CKINVDCx16_ASAP7_75t_R g499 ( .A(n_26), .Y(n_499) );
INVx1_ASAP7_75t_L g511 ( .A(n_27), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_28), .A2(n_144), .B(n_212), .C(n_226), .Y(n_225) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_29), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_30), .Y(n_467) );
AOI222xp33_ASAP7_75t_L g431 ( .A1(n_31), .A2(n_432), .B1(n_701), .B2(n_702), .C1(n_711), .C2(n_714), .Y(n_431) );
INVx1_ASAP7_75t_L g528 ( .A(n_32), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_33), .A2(n_164), .B(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g146 ( .A(n_34), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_35), .A2(n_159), .B(n_191), .C(n_192), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_36), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g492 ( .A1(n_37), .A2(n_179), .B(n_493), .C(n_495), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_38), .Y(n_124) );
INVxp67_ASAP7_75t_L g529 ( .A(n_39), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_40), .B(n_228), .Y(n_227) );
CKINVDCx14_ASAP7_75t_R g491 ( .A(n_41), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_42), .A2(n_144), .B(n_212), .C(n_510), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_L g458 ( .A1(n_44), .A2(n_181), .B(n_459), .C(n_460), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_45), .B(n_205), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g245 ( .A(n_46), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_47), .B(n_155), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_48), .B(n_164), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_49), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_50), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_51), .A2(n_159), .B(n_191), .C(n_252), .Y(n_251) );
OAI22xp5_ASAP7_75t_SL g702 ( .A1(n_52), .A2(n_703), .B1(n_704), .B2(n_710), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_52), .Y(n_710) );
INVx1_ASAP7_75t_L g178 ( .A(n_53), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_54), .A2(n_705), .B1(n_706), .B2(n_707), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_54), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_55), .A2(n_85), .B1(n_708), .B2(n_709), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_55), .Y(n_709) );
INVx1_ASAP7_75t_L g253 ( .A(n_56), .Y(n_253) );
INVx1_ASAP7_75t_L g449 ( .A(n_57), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_58), .B(n_164), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_59), .Y(n_216) );
CKINVDCx14_ASAP7_75t_R g457 ( .A(n_60), .Y(n_457) );
INVx1_ASAP7_75t_L g162 ( .A(n_61), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_62), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_63), .B(n_170), .Y(n_271) );
A2O1A1Ixp33_ASAP7_75t_L g268 ( .A1(n_64), .A2(n_151), .B(n_211), .C(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g140 ( .A(n_65), .Y(n_140) );
INVx1_ASAP7_75t_SL g494 ( .A(n_66), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_67), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_68), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_69), .B(n_155), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_70), .B(n_170), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_71), .B(n_156), .Y(n_242) );
INVx1_ASAP7_75t_L g502 ( .A(n_72), .Y(n_502) );
CKINVDCx16_ASAP7_75t_R g173 ( .A(n_73), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_74), .B(n_195), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g143 ( .A1(n_75), .A2(n_144), .B(n_149), .C(n_159), .Y(n_143) );
CKINVDCx16_ASAP7_75t_R g267 ( .A(n_76), .Y(n_267) );
INVx1_ASAP7_75t_L g113 ( .A(n_77), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_78), .A2(n_164), .B(n_456), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_79), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_80), .A2(n_164), .B(n_477), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_81), .A2(n_205), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g478 ( .A(n_82), .Y(n_478) );
CKINVDCx16_ASAP7_75t_R g508 ( .A(n_83), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_84), .B(n_194), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_85), .Y(n_708) );
CKINVDCx20_ASAP7_75t_R g200 ( .A(n_86), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g447 ( .A1(n_87), .A2(n_164), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g481 ( .A(n_88), .Y(n_481) );
INVx2_ASAP7_75t_L g138 ( .A(n_89), .Y(n_138) );
INVx1_ASAP7_75t_L g470 ( .A(n_90), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_91), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_92), .B(n_180), .Y(n_243) );
OR2x2_ASAP7_75t_L g424 ( .A(n_93), .B(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g435 ( .A(n_93), .B(n_426), .Y(n_435) );
INVx2_ASAP7_75t_L g439 ( .A(n_93), .Y(n_439) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_94), .A2(n_144), .B(n_159), .C(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_95), .B(n_164), .Y(n_189) );
INVx1_ASAP7_75t_L g193 ( .A(n_96), .Y(n_193) );
INVxp67_ASAP7_75t_L g270 ( .A(n_97), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_98), .B(n_136), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_99), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g150 ( .A(n_100), .Y(n_150) );
INVx1_ASAP7_75t_L g238 ( .A(n_101), .Y(n_238) );
INVx2_ASAP7_75t_L g452 ( .A(n_102), .Y(n_452) );
AND2x2_ASAP7_75t_L g255 ( .A(n_103), .B(n_198), .Y(n_255) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx12_ASAP7_75t_R g719 ( .A(n_107), .Y(n_719) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
AND2x2_ASAP7_75t_L g426 ( .A(n_108), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
AO21x1_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_120), .B(n_430), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_SL g718 ( .A(n_117), .Y(n_718) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI21xp5_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_422), .B(n_428), .Y(n_120) );
AOI22xp33_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_125), .B1(n_420), .B2(n_421), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_122), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_125), .Y(n_421) );
XNOR2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_129), .Y(n_125) );
INVx2_ASAP7_75t_L g436 ( .A(n_129), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_129), .A2(n_434), .B1(n_716), .B2(n_717), .Y(n_715) );
NAND2x1p5_ASAP7_75t_L g129 ( .A(n_130), .B(n_363), .Y(n_129) );
AND4x1_ASAP7_75t_L g130 ( .A(n_131), .B(n_303), .C(n_318), .D(n_343), .Y(n_130) );
NOR2xp33_ASAP7_75t_SL g131 ( .A(n_132), .B(n_276), .Y(n_131) );
OAI21xp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_184), .B(n_256), .Y(n_132) );
AND2x2_ASAP7_75t_L g306 ( .A(n_133), .B(n_202), .Y(n_306) );
AND2x2_ASAP7_75t_L g319 ( .A(n_133), .B(n_201), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_133), .B(n_185), .Y(n_369) );
INVx1_ASAP7_75t_L g373 ( .A(n_133), .Y(n_373) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_169), .Y(n_133) );
INVx2_ASAP7_75t_L g290 ( .A(n_134), .Y(n_290) );
BUFx2_ASAP7_75t_L g317 ( .A(n_134), .Y(n_317) );
AO21x2_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_142), .B(n_167), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_135), .B(n_168), .Y(n_167) );
INVx3_ASAP7_75t_L g170 ( .A(n_135), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_135), .B(n_200), .Y(n_199) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_135), .A2(n_237), .B(n_244), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_135), .B(n_474), .Y(n_473) );
AO21x2_ASAP7_75t_L g497 ( .A1(n_135), .A2(n_498), .B(n_504), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_135), .B(n_514), .Y(n_513) );
INVx4_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_136), .A2(n_224), .B(n_225), .Y(n_223) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_136), .Y(n_264) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g246 ( .A(n_137), .Y(n_246) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x2_ASAP7_75t_SL g198 ( .A(n_138), .B(n_139), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_163), .Y(n_142) );
INVx5_ASAP7_75t_L g174 ( .A(n_144), .Y(n_174) );
AND2x6_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_145), .Y(n_158) );
BUFx3_ASAP7_75t_L g182 ( .A(n_145), .Y(n_182) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g166 ( .A(n_146), .Y(n_166) );
INVx1_ASAP7_75t_L g232 ( .A(n_146), .Y(n_232) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_148), .Y(n_153) );
INVx3_ASAP7_75t_L g156 ( .A(n_148), .Y(n_156) );
AND2x2_ASAP7_75t_L g165 ( .A(n_148), .B(n_166), .Y(n_165) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_148), .Y(n_180) );
INVx1_ASAP7_75t_L g228 ( .A(n_148), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_154), .C(n_157), .Y(n_149) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_152), .B(n_452), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_152), .B(n_481), .Y(n_480) );
OAI22xp33_ASAP7_75t_L g527 ( .A1(n_152), .A2(n_155), .B1(n_528), .B2(n_529), .Y(n_527) );
INVx4_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g195 ( .A(n_153), .Y(n_195) );
INVx2_ASAP7_75t_L g176 ( .A(n_155), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_155), .B(n_270), .Y(n_269) );
O2A1O1Ixp33_ASAP7_75t_L g510 ( .A1(n_155), .A2(n_210), .B(n_511), .C(n_512), .Y(n_510) );
INVx5_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_156), .B(n_461), .Y(n_460) );
HB1xp67_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx3_ASAP7_75t_L g495 ( .A(n_158), .Y(n_495) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
O2A1O1Ixp33_ASAP7_75t_SL g172 ( .A1(n_160), .A2(n_173), .B(n_174), .C(n_175), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_L g266 ( .A1(n_160), .A2(n_174), .B(n_267), .C(n_268), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_SL g448 ( .A1(n_160), .A2(n_174), .B(n_449), .C(n_450), .Y(n_448) );
O2A1O1Ixp33_ASAP7_75t_SL g456 ( .A1(n_160), .A2(n_174), .B(n_457), .C(n_458), .Y(n_456) );
O2A1O1Ixp33_ASAP7_75t_SL g477 ( .A1(n_160), .A2(n_174), .B(n_478), .C(n_479), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_160), .A2(n_174), .B(n_491), .C(n_492), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_SL g524 ( .A1(n_160), .A2(n_174), .B(n_525), .C(n_526), .Y(n_524) );
INVx4_ASAP7_75t_SL g160 ( .A(n_161), .Y(n_160) );
AND2x4_ASAP7_75t_L g164 ( .A(n_161), .B(n_165), .Y(n_164) );
BUFx3_ASAP7_75t_L g212 ( .A(n_161), .Y(n_212) );
NAND2x1p5_ASAP7_75t_L g239 ( .A(n_161), .B(n_165), .Y(n_239) );
BUFx2_ASAP7_75t_L g205 ( .A(n_164), .Y(n_205) );
INVx1_ASAP7_75t_L g211 ( .A(n_166), .Y(n_211) );
AND2x2_ASAP7_75t_L g257 ( .A(n_169), .B(n_202), .Y(n_257) );
INVx2_ASAP7_75t_L g273 ( .A(n_169), .Y(n_273) );
AND2x2_ASAP7_75t_L g282 ( .A(n_169), .B(n_201), .Y(n_282) );
AND2x2_ASAP7_75t_L g361 ( .A(n_169), .B(n_290), .Y(n_361) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_183), .Y(n_169) );
INVx2_ASAP7_75t_L g191 ( .A(n_174), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_179), .B(n_494), .Y(n_493) );
INVx4_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g459 ( .A(n_180), .Y(n_459) );
INVx2_ASAP7_75t_L g472 ( .A(n_181), .Y(n_472) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_182), .Y(n_197) );
INVx1_ASAP7_75t_L g482 ( .A(n_182), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_185), .B(n_218), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_185), .B(n_288), .Y(n_326) );
INVx1_ASAP7_75t_L g414 ( .A(n_185), .Y(n_414) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_201), .Y(n_185) );
AND2x2_ASAP7_75t_L g272 ( .A(n_186), .B(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g286 ( .A(n_186), .B(n_287), .Y(n_286) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_186), .Y(n_315) );
OR2x2_ASAP7_75t_L g347 ( .A(n_186), .B(n_289), .Y(n_347) );
AND2x2_ASAP7_75t_L g355 ( .A(n_186), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g388 ( .A(n_186), .B(n_357), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_186), .B(n_257), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_186), .B(n_317), .Y(n_413) );
AND2x2_ASAP7_75t_L g419 ( .A(n_186), .B(n_306), .Y(n_419) );
INVx5_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
BUFx2_ASAP7_75t_L g279 ( .A(n_187), .Y(n_279) );
AND2x2_ASAP7_75t_L g309 ( .A(n_187), .B(n_289), .Y(n_309) );
AND2x2_ASAP7_75t_L g342 ( .A(n_187), .B(n_302), .Y(n_342) );
AND2x2_ASAP7_75t_L g362 ( .A(n_187), .B(n_202), .Y(n_362) );
AND2x2_ASAP7_75t_L g396 ( .A(n_187), .B(n_262), .Y(n_396) );
OR2x6_ASAP7_75t_L g187 ( .A(n_188), .B(n_199), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_198), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_196), .C(n_197), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_194), .A2(n_197), .B(n_253), .C(n_254), .Y(n_252) );
O2A1O1Ixp5_ASAP7_75t_L g469 ( .A1(n_194), .A2(n_470), .B(n_471), .C(n_472), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_194), .A2(n_472), .B(n_502), .C(n_503), .Y(n_501) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g214 ( .A(n_198), .Y(n_214) );
INVx1_ASAP7_75t_L g217 ( .A(n_198), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_198), .A2(n_250), .B(n_251), .Y(n_249) );
OA21x2_ASAP7_75t_L g454 ( .A1(n_198), .A2(n_455), .B(n_462), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_L g507 ( .A1(n_198), .A2(n_239), .B(n_508), .C(n_509), .Y(n_507) );
AND2x4_ASAP7_75t_L g302 ( .A(n_201), .B(n_273), .Y(n_302) );
AND2x2_ASAP7_75t_L g313 ( .A(n_201), .B(n_309), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_201), .B(n_289), .Y(n_352) );
INVx2_ASAP7_75t_L g367 ( .A(n_201), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_201), .B(n_301), .Y(n_390) );
AND2x2_ASAP7_75t_L g409 ( .A(n_201), .B(n_361), .Y(n_409) );
INVx5_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_202), .Y(n_308) );
AND2x2_ASAP7_75t_L g316 ( .A(n_202), .B(n_317), .Y(n_316) );
AND2x4_ASAP7_75t_L g357 ( .A(n_202), .B(n_273), .Y(n_357) );
OR2x6_ASAP7_75t_L g202 ( .A(n_203), .B(n_215), .Y(n_202) );
AOI21xp5_ASAP7_75t_SL g203 ( .A1(n_204), .A2(n_206), .B(n_213), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_210), .Y(n_207) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_211), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_214), .B(n_505), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_216), .B(n_217), .Y(n_215) );
AO21x2_ASAP7_75t_L g465 ( .A1(n_217), .A2(n_466), .B(n_473), .Y(n_465) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_220), .B(n_233), .Y(n_219) );
AND2x2_ASAP7_75t_L g280 ( .A(n_220), .B(n_263), .Y(n_280) );
INVx1_ASAP7_75t_SL g220 ( .A(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_221), .B(n_236), .Y(n_260) );
OR2x2_ASAP7_75t_L g293 ( .A(n_221), .B(n_263), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_221), .B(n_263), .Y(n_298) );
AND2x2_ASAP7_75t_L g325 ( .A(n_221), .B(n_262), .Y(n_325) );
AND2x2_ASAP7_75t_L g377 ( .A(n_221), .B(n_235), .Y(n_377) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_222), .B(n_247), .Y(n_285) );
AND2x2_ASAP7_75t_L g321 ( .A(n_222), .B(n_236), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_229), .B(n_230), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_230), .A2(n_242), .B(n_243), .Y(n_241) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx3_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_233), .B(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
OR2x2_ASAP7_75t_L g311 ( .A(n_234), .B(n_293), .Y(n_311) );
OR2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_247), .Y(n_234) );
OAI322xp33_ASAP7_75t_L g276 ( .A1(n_235), .A2(n_277), .A3(n_281), .B1(n_283), .B2(n_286), .C1(n_291), .C2(n_299), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_235), .B(n_262), .Y(n_284) );
OR2x2_ASAP7_75t_L g294 ( .A(n_235), .B(n_248), .Y(n_294) );
AND2x2_ASAP7_75t_L g296 ( .A(n_235), .B(n_248), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_235), .B(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_235), .B(n_263), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_235), .B(n_392), .Y(n_391) );
INVx5_ASAP7_75t_SL g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_236), .B(n_280), .Y(n_406) );
OAI21xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B(n_240), .Y(n_237) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_239), .A2(n_467), .B(n_468), .Y(n_466) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_239), .A2(n_499), .B(n_500), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
INVx2_ASAP7_75t_L g522 ( .A(n_246), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_247), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g274 ( .A(n_247), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_247), .B(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g336 ( .A(n_247), .B(n_263), .Y(n_336) );
AOI211xp5_ASAP7_75t_SL g364 ( .A1(n_247), .A2(n_365), .B(n_368), .C(n_380), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_247), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g402 ( .A(n_247), .B(n_377), .Y(n_402) );
INVx5_ASAP7_75t_SL g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g330 ( .A(n_248), .B(n_263), .Y(n_330) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_248), .Y(n_339) );
AND2x2_ASAP7_75t_L g379 ( .A(n_248), .B(n_377), .Y(n_379) );
AND2x2_ASAP7_75t_SL g410 ( .A(n_248), .B(n_280), .Y(n_410) );
AND2x2_ASAP7_75t_L g417 ( .A(n_248), .B(n_376), .Y(n_417) );
OR2x6_ASAP7_75t_L g248 ( .A(n_249), .B(n_255), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_258), .B1(n_272), .B2(n_274), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_257), .B(n_279), .Y(n_327) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
INVx1_ASAP7_75t_L g275 ( .A(n_260), .Y(n_275) );
OR2x2_ASAP7_75t_L g335 ( .A(n_260), .B(n_336), .Y(n_335) );
OAI221xp5_ASAP7_75t_SL g383 ( .A1(n_260), .A2(n_384), .B1(n_386), .B2(n_387), .C(n_389), .Y(n_383) );
INVx2_ASAP7_75t_L g322 ( .A(n_261), .Y(n_322) );
AND2x2_ASAP7_75t_L g295 ( .A(n_262), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g385 ( .A(n_262), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_262), .B(n_377), .Y(n_398) );
INVx3_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVxp67_ASAP7_75t_L g340 ( .A(n_263), .Y(n_340) );
AND2x2_ASAP7_75t_L g376 ( .A(n_263), .B(n_377), .Y(n_376) );
OA21x2_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_265), .B(n_271), .Y(n_263) );
OA21x2_ASAP7_75t_L g446 ( .A1(n_264), .A2(n_447), .B(n_453), .Y(n_446) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_264), .A2(n_476), .B(n_483), .Y(n_475) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_264), .A2(n_489), .B(n_496), .Y(n_488) );
AND2x2_ASAP7_75t_L g378 ( .A(n_272), .B(n_317), .Y(n_378) );
AND2x2_ASAP7_75t_L g288 ( .A(n_273), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_273), .B(n_346), .Y(n_345) );
NOR2xp33_ASAP7_75t_SL g359 ( .A(n_275), .B(n_322), .Y(n_359) );
INVx1_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g365 ( .A(n_278), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
OR2x2_ASAP7_75t_L g351 ( .A(n_279), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g416 ( .A(n_279), .B(n_361), .Y(n_416) );
INVx2_ASAP7_75t_L g349 ( .A(n_280), .Y(n_349) );
NAND4xp25_ASAP7_75t_SL g412 ( .A(n_281), .B(n_413), .C(n_414), .D(n_415), .Y(n_412) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_282), .B(n_346), .Y(n_381) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx1_ASAP7_75t_SL g418 ( .A(n_285), .Y(n_418) );
O2A1O1Ixp33_ASAP7_75t_SL g380 ( .A1(n_286), .A2(n_349), .B(n_353), .C(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g375 ( .A(n_288), .B(n_367), .Y(n_375) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_289), .Y(n_301) );
INVx1_ASAP7_75t_L g356 ( .A(n_289), .Y(n_356) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_290), .Y(n_333) );
AOI211xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_294), .B(n_295), .C(n_297), .Y(n_291) );
AND2x2_ASAP7_75t_L g312 ( .A(n_292), .B(n_296), .Y(n_312) );
OAI322xp33_ASAP7_75t_SL g350 ( .A1(n_292), .A2(n_351), .A3(n_353), .B1(n_354), .B2(n_358), .C1(n_359), .C2(n_360), .Y(n_350) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g372 ( .A(n_294), .B(n_298), .Y(n_372) );
INVx1_ASAP7_75t_L g353 ( .A(n_296), .Y(n_353) );
INVx1_ASAP7_75t_SL g371 ( .A(n_298), .Y(n_371) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
AOI222xp33_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_310), .B1(n_312), .B2(n_313), .C1(n_314), .C2(n_721), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g304 ( .A(n_305), .B(n_307), .Y(n_304) );
OAI322xp33_ASAP7_75t_L g393 ( .A1(n_305), .A2(n_367), .A3(n_372), .B1(n_394), .B2(n_395), .C1(n_397), .C2(n_398), .Y(n_393) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AOI221xp5_ASAP7_75t_L g343 ( .A1(n_306), .A2(n_320), .B1(n_344), .B2(n_348), .C(n_350), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx1_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
OAI222xp33_ASAP7_75t_L g323 ( .A1(n_311), .A2(n_324), .B1(n_326), .B2(n_327), .C1(n_328), .C2(n_331), .Y(n_323) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_313), .A2(n_320), .B1(n_390), .B2(n_391), .Y(n_389) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
AOI211xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_320), .B(n_323), .C(n_334), .Y(n_318) );
O2A1O1Ixp33_ASAP7_75t_L g399 ( .A1(n_320), .A2(n_357), .B(n_400), .C(n_403), .Y(n_399) );
AND2x4_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
AND2x2_ASAP7_75t_L g329 ( .A(n_321), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_SL g392 ( .A(n_325), .Y(n_392) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_332), .B(n_357), .Y(n_386) );
BUFx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AOI21xp33_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_337), .B(n_341), .Y(n_334) );
OAI221xp5_ASAP7_75t_SL g403 ( .A1(n_335), .A2(n_404), .B1(n_405), .B2(n_406), .C(n_407), .Y(n_403) );
INVxp33_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_339), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_346), .B(n_357), .Y(n_397) );
INVx2_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_357), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
AND2x2_ASAP7_75t_L g408 ( .A(n_361), .B(n_367), .Y(n_408) );
AND4x1_ASAP7_75t_L g363 ( .A(n_364), .B(n_382), .C(n_399), .D(n_411), .Y(n_363) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OAI221xp5_ASAP7_75t_SL g368 ( .A1(n_369), .A2(n_370), .B1(n_372), .B2(n_373), .C(n_374), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_376), .B1(n_378), .B2(n_379), .Y(n_374) );
INVx1_ASAP7_75t_L g404 ( .A(n_375), .Y(n_404) );
INVx1_ASAP7_75t_SL g394 ( .A(n_379), .Y(n_394) );
NOR2xp33_ASAP7_75t_SL g382 ( .A(n_383), .B(n_393), .Y(n_382) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_395), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_402), .A2(n_408), .B1(n_409), .B2(n_410), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_417), .B1(n_418), .B2(n_419), .Y(n_411) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_SL g429 ( .A(n_424), .Y(n_429) );
NOR2x2_ASAP7_75t_L g713 ( .A(n_425), .B(n_439), .Y(n_713) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OR2x2_ASAP7_75t_L g438 ( .A(n_426), .B(n_439), .Y(n_438) );
AOI21xp33_ASAP7_75t_SL g430 ( .A1(n_428), .A2(n_431), .B(n_718), .Y(n_430) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_436), .B1(n_437), .B2(n_440), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx6_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g716 ( .A(n_438), .Y(n_716) );
BUFx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g717 ( .A(n_441), .Y(n_717) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_627), .Y(n_441) );
NOR4xp25_ASAP7_75t_L g442 ( .A(n_443), .B(n_569), .C(n_599), .D(n_609), .Y(n_442) );
OAI211xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_484), .B(n_532), .C(n_559), .Y(n_443) );
OAI222xp33_ASAP7_75t_L g654 ( .A1(n_444), .A2(n_574), .B1(n_655), .B2(n_656), .C1(n_657), .C2(n_658), .Y(n_654) );
OR2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_463), .Y(n_444) );
AOI33xp33_ASAP7_75t_L g580 ( .A1(n_445), .A2(n_567), .A3(n_568), .B1(n_581), .B2(n_586), .B3(n_588), .Y(n_580) );
OAI211xp5_ASAP7_75t_SL g637 ( .A1(n_445), .A2(n_638), .B(n_640), .C(n_642), .Y(n_637) );
OR2x2_ASAP7_75t_L g653 ( .A(n_445), .B(n_639), .Y(n_653) );
INVx1_ASAP7_75t_L g686 ( .A(n_445), .Y(n_686) );
OR2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_454), .Y(n_445) );
INVx2_ASAP7_75t_L g563 ( .A(n_446), .Y(n_563) );
AND2x2_ASAP7_75t_L g579 ( .A(n_446), .B(n_475), .Y(n_579) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_446), .Y(n_614) );
AND2x2_ASAP7_75t_L g643 ( .A(n_446), .B(n_454), .Y(n_643) );
INVx2_ASAP7_75t_L g543 ( .A(n_454), .Y(n_543) );
BUFx3_ASAP7_75t_L g551 ( .A(n_454), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_454), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g562 ( .A(n_454), .B(n_563), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_454), .B(n_464), .Y(n_591) );
AND2x2_ASAP7_75t_L g660 ( .A(n_454), .B(n_594), .Y(n_660) );
INVx2_ASAP7_75t_SL g554 ( .A(n_463), .Y(n_554) );
OR2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_475), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_464), .B(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g596 ( .A(n_464), .Y(n_596) );
AND2x2_ASAP7_75t_L g607 ( .A(n_464), .B(n_563), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_464), .B(n_592), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_464), .B(n_594), .Y(n_639) );
AND2x2_ASAP7_75t_L g698 ( .A(n_464), .B(n_643), .Y(n_698) );
INVx4_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g568 ( .A(n_465), .B(n_475), .Y(n_568) );
AND2x2_ASAP7_75t_L g578 ( .A(n_465), .B(n_579), .Y(n_578) );
BUFx3_ASAP7_75t_L g600 ( .A(n_465), .Y(n_600) );
AND3x2_ASAP7_75t_L g659 ( .A(n_465), .B(n_660), .C(n_661), .Y(n_659) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_475), .Y(n_550) );
INVx1_ASAP7_75t_SL g594 ( .A(n_475), .Y(n_594) );
NAND3xp33_ASAP7_75t_L g606 ( .A(n_475), .B(n_543), .C(n_607), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_485), .B(n_515), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g629 ( .A1(n_485), .A2(n_578), .B(n_630), .C(n_632), .Y(n_629) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_487), .B(n_506), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_487), .B(n_636), .Y(n_635) );
INVx2_ASAP7_75t_SL g646 ( .A(n_487), .Y(n_646) );
AND2x2_ASAP7_75t_L g667 ( .A(n_487), .B(n_517), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_487), .B(n_576), .Y(n_695) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_497), .Y(n_487) );
AND2x2_ASAP7_75t_L g540 ( .A(n_488), .B(n_531), .Y(n_540) );
INVx2_ASAP7_75t_L g547 ( .A(n_488), .Y(n_547) );
AND2x2_ASAP7_75t_L g567 ( .A(n_488), .B(n_517), .Y(n_567) );
AND2x2_ASAP7_75t_L g617 ( .A(n_488), .B(n_506), .Y(n_617) );
INVx1_ASAP7_75t_L g621 ( .A(n_488), .Y(n_621) );
INVx2_ASAP7_75t_SL g531 ( .A(n_497), .Y(n_531) );
BUFx2_ASAP7_75t_L g557 ( .A(n_497), .Y(n_557) );
AND2x2_ASAP7_75t_L g684 ( .A(n_497), .B(n_506), .Y(n_684) );
INVx3_ASAP7_75t_SL g517 ( .A(n_506), .Y(n_517) );
AND2x2_ASAP7_75t_L g539 ( .A(n_506), .B(n_540), .Y(n_539) );
AND2x4_ASAP7_75t_L g546 ( .A(n_506), .B(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g576 ( .A(n_506), .B(n_536), .Y(n_576) );
OR2x2_ASAP7_75t_L g585 ( .A(n_506), .B(n_531), .Y(n_585) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_506), .Y(n_603) );
AND2x2_ASAP7_75t_L g608 ( .A(n_506), .B(n_561), .Y(n_608) );
AND2x2_ASAP7_75t_L g636 ( .A(n_506), .B(n_519), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_506), .B(n_672), .Y(n_671) );
OR2x2_ASAP7_75t_L g674 ( .A(n_506), .B(n_518), .Y(n_674) );
OR2x6_ASAP7_75t_L g506 ( .A(n_507), .B(n_513), .Y(n_506) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
AND2x2_ASAP7_75t_L g598 ( .A(n_517), .B(n_547), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_517), .B(n_540), .Y(n_626) );
AND2x2_ASAP7_75t_L g644 ( .A(n_517), .B(n_561), .Y(n_644) );
OR2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_531), .Y(n_518) );
AND2x2_ASAP7_75t_L g545 ( .A(n_519), .B(n_531), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_519), .B(n_574), .Y(n_573) );
BUFx3_ASAP7_75t_L g583 ( .A(n_519), .Y(n_583) );
OR2x2_ASAP7_75t_L g631 ( .A(n_519), .B(n_551), .Y(n_631) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_523), .B(n_530), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AO21x2_ASAP7_75t_L g536 ( .A1(n_521), .A2(n_537), .B(n_538), .Y(n_536) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g537 ( .A(n_523), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_530), .Y(n_538) );
AND2x2_ASAP7_75t_L g566 ( .A(n_531), .B(n_536), .Y(n_566) );
INVx1_ASAP7_75t_L g574 ( .A(n_531), .Y(n_574) );
AND2x2_ASAP7_75t_L g669 ( .A(n_531), .B(n_547), .Y(n_669) );
AOI222xp33_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_541), .B1(n_544), .B2(n_548), .C1(n_552), .C2(n_555), .Y(n_532) );
INVx1_ASAP7_75t_L g664 ( .A(n_533), .Y(n_664) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_539), .Y(n_533) );
AND2x2_ASAP7_75t_L g560 ( .A(n_534), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g571 ( .A(n_534), .B(n_540), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_534), .B(n_562), .Y(n_587) );
OAI222xp33_ASAP7_75t_L g609 ( .A1(n_534), .A2(n_610), .B1(n_615), .B2(n_616), .C1(n_624), .C2(n_626), .Y(n_609) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g597 ( .A(n_536), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_536), .B(n_617), .Y(n_657) );
AND2x2_ASAP7_75t_L g668 ( .A(n_536), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g676 ( .A(n_539), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g655 ( .A(n_541), .B(n_592), .Y(n_655) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_543), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g613 ( .A(n_543), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
INVx3_ASAP7_75t_L g558 ( .A(n_546), .Y(n_558) );
O2A1O1Ixp33_ASAP7_75t_L g648 ( .A1(n_546), .A2(n_649), .B(n_652), .C(n_654), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_546), .B(n_583), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_546), .B(n_566), .Y(n_688) );
AND2x2_ASAP7_75t_L g561 ( .A(n_547), .B(n_557), .Y(n_561) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
INVx1_ASAP7_75t_L g588 ( .A(n_550), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_551), .B(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g640 ( .A(n_551), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g679 ( .A(n_551), .B(n_579), .Y(n_679) );
INVx1_ASAP7_75t_L g691 ( .A(n_551), .Y(n_691) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_554), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
INVx1_ASAP7_75t_L g672 ( .A(n_557), .Y(n_672) );
A2O1A1Ixp33_ASAP7_75t_SL g559 ( .A1(n_560), .A2(n_562), .B(n_564), .C(n_568), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_560), .A2(n_590), .B1(n_605), .B2(n_608), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_561), .B(n_575), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_561), .B(n_583), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_562), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_SL g625 ( .A(n_562), .Y(n_625) );
AND2x2_ASAP7_75t_L g632 ( .A(n_562), .B(n_612), .Y(n_632) );
INVx2_ASAP7_75t_L g593 ( .A(n_563), .Y(n_593) );
INVxp67_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
NOR4xp25_ASAP7_75t_L g570 ( .A(n_567), .B(n_571), .C(n_572), .D(n_575), .Y(n_570) );
INVx1_ASAP7_75t_SL g641 ( .A(n_568), .Y(n_641) );
AND2x2_ASAP7_75t_L g685 ( .A(n_568), .B(n_686), .Y(n_685) );
OAI211xp5_ASAP7_75t_SL g569 ( .A1(n_570), .A2(n_577), .B(n_580), .C(n_589), .Y(n_569) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_576), .B(n_646), .Y(n_697) );
AOI22xp5_ASAP7_75t_L g696 ( .A1(n_578), .A2(n_697), .B1(n_698), .B2(n_699), .Y(n_696) );
INVx1_ASAP7_75t_SL g651 ( .A(n_579), .Y(n_651) );
AND2x2_ASAP7_75t_L g690 ( .A(n_579), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_583), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_587), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_588), .B(n_613), .Y(n_673) );
OAI21xp5_ASAP7_75t_SL g589 ( .A1(n_590), .A2(n_595), .B(n_597), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx1_ASAP7_75t_L g665 ( .A(n_592), .Y(n_665) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
INVx2_ASAP7_75t_L g693 ( .A(n_593), .Y(n_693) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_594), .Y(n_620) );
OAI21xp33_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_601), .B(n_604), .Y(n_599) );
CKINVDCx16_ASAP7_75t_R g612 ( .A(n_600), .Y(n_612) );
OR2x2_ASAP7_75t_L g650 ( .A(n_600), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AOI21xp33_ASAP7_75t_SL g645 ( .A1(n_603), .A2(n_646), .B(n_647), .Y(n_645) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AOI221xp5_ASAP7_75t_L g633 ( .A1(n_607), .A2(n_634), .B1(n_637), .B2(n_644), .C(n_645), .Y(n_633) );
INVx1_ASAP7_75t_SL g677 ( .A(n_608), .Y(n_677) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
OR2x2_ASAP7_75t_L g624 ( .A(n_612), .B(n_625), .Y(n_624) );
INVxp67_ASAP7_75t_L g661 ( .A(n_614), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_618), .B1(n_621), .B2(n_622), .Y(n_616) );
INVx1_ASAP7_75t_L g656 ( .A(n_617), .Y(n_656) );
INVxp67_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_620), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NOR4xp25_ASAP7_75t_L g627 ( .A(n_628), .B(n_662), .C(n_675), .D(n_687), .Y(n_627) );
NAND3xp33_ASAP7_75t_SL g628 ( .A(n_629), .B(n_633), .C(n_648), .Y(n_628) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_631), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_638), .B(n_643), .Y(n_647) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OAI221xp5_ASAP7_75t_SL g675 ( .A1(n_650), .A2(n_676), .B1(n_677), .B2(n_678), .C(n_680), .Y(n_675) );
O2A1O1Ixp33_ASAP7_75t_L g666 ( .A1(n_652), .A2(n_667), .B(n_668), .C(n_670), .Y(n_666) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g670 ( .A1(n_653), .A2(n_671), .B1(n_673), .B2(n_674), .Y(n_670) );
INVx2_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
A2O1A1Ixp33_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_664), .B(n_665), .C(n_666), .Y(n_662) );
INVx1_ASAP7_75t_L g681 ( .A(n_674), .Y(n_681) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OAI21xp5_ASAP7_75t_SL g680 ( .A1(n_681), .A2(n_682), .B(n_685), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OAI221xp5_ASAP7_75t_SL g687 ( .A1(n_688), .A2(n_689), .B1(n_692), .B2(n_694), .C(n_696), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVxp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
INVx3_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
endmodule