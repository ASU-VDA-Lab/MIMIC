module fake_jpeg_231_n_191 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_191);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_191;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_33),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_32),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_27),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_16),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_31),
.B(n_19),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_35),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_9),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_80),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_73),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_80),
.A2(n_70),
.B1(n_64),
.B2(n_61),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_82),
.A2(n_89),
.B1(n_72),
.B2(n_77),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_54),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_88),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_78),
.B(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_87),
.B(n_1),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_75),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_70),
.B1(n_59),
.B2(n_66),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_59),
.B1(n_61),
.B2(n_73),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_81),
.B1(n_69),
.B2(n_52),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_53),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_62),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_88),
.A2(n_68),
.B1(n_55),
.B2(n_56),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_103),
.B1(n_98),
.B2(n_112),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_95),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_102),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_112),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_86),
.B(n_60),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_71),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_85),
.A2(n_58),
.B1(n_57),
.B2(n_63),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_91),
.B(n_0),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_110),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_113),
.Y(n_119)
);

AND2x4_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_69),
.Y(n_108)
);

NAND2xp33_ASAP7_75t_SL g114 ( 
.A(n_108),
.B(n_72),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_109),
.A2(n_111),
.B(n_76),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_91),
.B(n_0),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_84),
.A2(n_77),
.B1(n_76),
.B2(n_79),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_114),
.Y(n_148)
);

NOR2x1_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_130),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_108),
.A2(n_90),
.B1(n_93),
.B2(n_79),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_125),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_108),
.A2(n_100),
.B1(n_96),
.B2(n_99),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_8),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_108),
.A2(n_90),
.B(n_71),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_6),
.B(n_7),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_71),
.B1(n_3),
.B2(n_4),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_2),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_126),
.B(n_132),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_2),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_127),
.B(n_128),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_100),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_133),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_4),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_5),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_6),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_23),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_124),
.C(n_120),
.Y(n_153)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_137),
.Y(n_155)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

AO21x1_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_10),
.B(n_11),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_142),
.A2(n_141),
.B1(n_150),
.B2(n_139),
.Y(n_156)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_119),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_26),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_8),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_152),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_28),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_153),
.B(n_163),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_142),
.A2(n_120),
.B1(n_10),
.B2(n_11),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_154),
.A2(n_156),
.B1(n_134),
.B2(n_135),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_146),
.C(n_144),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_25),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_146),
.A2(n_144),
.B(n_120),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_162),
.A2(n_167),
.B(n_168),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_9),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_164),
.B(n_166),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_12),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_30),
.B(n_47),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_140),
.A2(n_29),
.B(n_45),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_170),
.A2(n_171),
.B1(n_174),
.B2(n_176),
.Y(n_178)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_165),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_153),
.C(n_168),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_161),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_177),
.B(n_181),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_172),
.A2(n_156),
.B1(n_157),
.B2(n_154),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_173),
.B1(n_17),
.B2(n_16),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_158),
.C(n_162),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_173),
.C(n_22),
.Y(n_184)
);

AOI321xp33_ASAP7_75t_L g181 ( 
.A1(n_169),
.A2(n_159),
.A3(n_164),
.B1(n_160),
.B2(n_34),
.C(n_37),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_182),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_177),
.B(n_180),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_185),
.A2(n_184),
.B(n_183),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_48),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_188),
.A2(n_186),
.B(n_41),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_189),
.B(n_42),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_178),
.Y(n_191)
);


endmodule