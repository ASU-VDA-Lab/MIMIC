module real_jpeg_33952_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx2_ASAP7_75t_L g94 ( 
.A(n_0),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_0),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_1),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_1),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_1),
.B(n_372),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_1),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_2),
.B(n_40),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_2),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_2),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_2),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g96 ( 
.A(n_2),
.B(n_86),
.Y(n_96)
);

AND2x4_ASAP7_75t_SL g108 ( 
.A(n_2),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_2),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_2),
.B(n_37),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_3),
.B(n_23),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_4),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_4),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_4),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_4),
.B(n_118),
.Y(n_117)
);

AND2x4_ASAP7_75t_L g201 ( 
.A(n_4),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_4),
.B(n_212),
.Y(n_211)
);

NAND2x1_ASAP7_75t_SL g232 ( 
.A(n_4),
.B(n_233),
.Y(n_232)
);

NAND2xp33_ASAP7_75t_R g282 ( 
.A(n_4),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_5),
.B(n_86),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_5),
.B(n_193),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_5),
.A2(n_279),
.B(n_281),
.Y(n_278)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_5),
.Y(n_342)
);

NAND2x1_ASAP7_75t_SL g374 ( 
.A(n_5),
.B(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_5),
.B(n_279),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_6),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_6),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_6),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_7),
.Y(n_341)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_8),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_8),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_9),
.B(n_57),
.Y(n_56)
);

AND2x4_ASAP7_75t_SL g65 ( 
.A(n_9),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_9),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_9),
.B(n_53),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_9),
.B(n_86),
.Y(n_85)
);

AND2x4_ASAP7_75t_L g98 ( 
.A(n_9),
.B(n_81),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g151 ( 
.A(n_9),
.B(n_152),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_9),
.B(n_209),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_10),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_10),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_11),
.A2(n_19),
.B(n_22),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_12),
.Y(n_121)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_14),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_14),
.B(n_172),
.Y(n_171)
);

AND2x2_ASAP7_75t_SL g292 ( 
.A(n_14),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_14),
.B(n_35),
.Y(n_302)
);

AND2x2_ASAP7_75t_SL g343 ( 
.A(n_14),
.B(n_344),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_15),
.B(n_86),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_15),
.B(n_79),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_15),
.B(n_386),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_16),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_17),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_17),
.B(n_103),
.Y(n_102)
);

AND2x4_ASAP7_75t_L g126 ( 
.A(n_17),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_17),
.B(n_166),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g289 ( 
.A(n_17),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_17),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_17),
.B(n_333),
.Y(n_332)
);

BUFx12f_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx12f_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

A2O1A1O1Ixp25_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_96),
.B(n_257),
.C(n_422),
.D(n_430),
.Y(n_23)
);

NOR3xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_223),
.C(n_248),
.Y(n_24)
);

NAND2x1_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_176),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_27),
.A2(n_425),
.B(n_426),
.Y(n_424)
);

NOR2x1_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_136),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_28),
.B(n_136),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_99),
.Y(n_28)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_29),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_73),
.C(n_88),
.Y(n_29)
);

INVxp33_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_31),
.B(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_48),
.C(n_64),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_32),
.B(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_45),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_38),
.B1(n_39),
.B2(n_44),
.Y(n_33)
);

INVxp67_ASAP7_75t_SL g44 ( 
.A(n_34),
.Y(n_44)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_37),
.Y(n_393)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_38),
.A2(n_39),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_38),
.A2(n_39),
.B1(n_337),
.B2(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_39),
.B(n_44),
.C(n_95),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_39),
.B(n_102),
.C(n_107),
.Y(n_135)
);

MAJx2_ASAP7_75t_L g336 ( 
.A(n_39),
.B(n_337),
.C(n_343),
.Y(n_336)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_43),
.Y(n_213)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_45),
.B(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_47),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_48),
.B(n_64),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_55),
.C(n_59),
.Y(n_48)
);

OAI22x1_ASAP7_75t_L g156 ( 
.A1(n_49),
.A2(n_50),
.B1(n_59),
.B2(n_60),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_54),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_54),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_55),
.B(n_107),
.C(n_299),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_55),
.A2(n_56),
.B1(n_299),
.B2(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

XNOR2x1_ASAP7_75t_L g155 ( 
.A(n_56),
.B(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_63),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_65),
.B(n_69),
.C(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_65),
.A2(n_214),
.B1(n_215),
.B2(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_65),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_65),
.B(n_133),
.C(n_214),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_67),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_67),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_71),
.Y(n_68)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_69),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_69),
.A2(n_194),
.B1(n_352),
.B2(n_354),
.Y(n_351)
);

INVxp33_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_74),
.B(n_88),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_85),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_78),
.B2(n_84),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_76),
.B(n_78),
.C(n_85),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_76),
.B(n_165),
.C(n_169),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_76),
.A2(n_77),
.B1(n_169),
.B2(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_83),
.Y(n_280)
);

FAx1_ASAP7_75t_SL g251 ( 
.A(n_85),
.B(n_252),
.CI(n_253),
.CON(n_251),
.SN(n_251)
);

NOR3xp33_ASAP7_75t_L g430 ( 
.A(n_85),
.B(n_145),
.C(n_214),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_87),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_96),
.C(n_97),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_89),
.B(n_160),
.Y(n_159)
);

MAJx2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_92),
.C(n_95),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_90),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_90),
.A2(n_145),
.B1(n_214),
.B2(n_215),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_92),
.A2(n_143),
.B1(n_144),
.B2(n_146),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_92),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_92),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_92),
.B(n_151),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_92),
.B(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_94),
.Y(n_209)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_94),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_96),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_97),
.A2(n_98),
.B1(n_117),
.B2(n_122),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_97),
.B(n_164),
.C(n_171),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_97),
.A2(n_98),
.B1(n_171),
.B2(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_98),
.B(n_122),
.C(n_123),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_113),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_100),
.B(n_113),
.C(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_110),
.C(n_111),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_138),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_106),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_108),
.B1(n_130),
.B2(n_133),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_107),
.B(n_130),
.C(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_107),
.B(n_398),
.Y(n_397)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_111),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_124),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_115),
.B(n_135),
.C(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_123),
.Y(n_115)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_134),
.Y(n_124)
);

INVxp33_ASAP7_75t_L g227 ( 
.A(n_125),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_126),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_130),
.A2(n_133),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_130),
.A2(n_133),
.B1(n_192),
.B2(n_353),
.Y(n_352)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_133),
.B(n_192),
.C(n_194),
.Y(n_191)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.C(n_173),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_137),
.B(n_174),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_139),
.B(n_222),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_157),
.C(n_162),
.Y(n_139)
);

INVxp33_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_180),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_147),
.C(n_155),
.Y(n_141)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_142),
.Y(n_270)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XOR2x1_ASAP7_75t_L g271 ( 
.A(n_147),
.B(n_155),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_150),
.B(n_154),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_148),
.A2(n_149),
.B1(n_151),
.B2(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_151),
.B(n_331),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_151),
.A2(n_197),
.B1(n_331),
.B2(n_332),
.Y(n_368)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_154),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_158),
.A2(n_159),
.B1(n_162),
.B2(n_163),
.Y(n_180)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_164),
.B(n_219),
.Y(n_218)
);

INVxp67_ASAP7_75t_SL g188 ( 
.A(n_165),
.Y(n_188)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_170),
.Y(n_387)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_221),
.Y(n_176)
);

NAND2x1p5_ASAP7_75t_L g425 ( 
.A(n_177),
.B(n_221),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.C(n_184),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_179),
.B(n_182),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_184),
.B(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_198),
.C(n_216),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_185),
.A2(n_186),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_191),
.C(n_195),
.Y(n_186)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_187),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_191),
.B(n_195),
.Y(n_322)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_192),
.Y(n_353)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_193),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_198),
.A2(n_217),
.B1(n_218),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_198),
.Y(n_266)
);

MAJx2_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_210),
.C(n_214),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_199),
.A2(n_200),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.C(n_208),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_201),
.B(n_204),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_208),
.B(n_276),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_210),
.A2(n_211),
.B1(n_214),
.B2(n_215),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_211),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_212),
.Y(n_301)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

A2O1A1O1Ixp25_ASAP7_75t_L g423 ( 
.A1(n_224),
.A2(n_249),
.B(n_424),
.C(n_427),
.D(n_428),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_246),
.Y(n_224)
);

NOR2xp67_ASAP7_75t_L g427 ( 
.A(n_225),
.B(n_246),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_229),
.C(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

INVxp33_ASAP7_75t_L g256 ( 
.A(n_230),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_240),
.B1(n_244),
.B2(n_245),
.Y(n_230)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_231),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_236),
.B1(n_238),
.B2(n_239),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_232),
.Y(n_238)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_236),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_238),
.C(n_245),
.Y(n_254)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_240),
.Y(n_245)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_255),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_250),
.B(n_255),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.Y(n_250)
);

BUFx24_ASAP7_75t_SL g432 ( 
.A(n_251),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_252),
.B(n_429),
.Y(n_428)
);

INVxp33_ASAP7_75t_SL g257 ( 
.A(n_258),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_356),
.B(n_419),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_309),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_260),
.A2(n_420),
.B(n_421),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_307),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_261),
.B(n_307),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_267),
.C(n_272),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_263),
.A2(n_268),
.B1(n_269),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_263),
.Y(n_312)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_272),
.B(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_272),
.B(n_311),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_295),
.C(n_303),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_274),
.B(n_318),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.C(n_284),
.Y(n_274)
);

XNOR2x1_ASAP7_75t_L g410 ( 
.A(n_275),
.B(n_411),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_277),
.A2(n_278),
.B1(n_284),
.B2(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NOR2xp67_ASAP7_75t_SL g400 ( 
.A(n_278),
.B(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_282),
.B(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_284),
.Y(n_412)
);

MAJx2_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_289),
.C(n_292),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_285),
.A2(n_286),
.B1(n_289),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_289),
.Y(n_328)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_292),
.B(n_327),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_294),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_304),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_300),
.C(n_302),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_298),
.Y(n_350)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_299),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_300),
.B(n_302),
.Y(n_349)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_305),
.Y(n_306)
);

NAND3xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_313),
.C(n_355),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_310),
.A2(n_313),
.B(n_355),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_319),
.C(n_323),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_316),
.A2(n_317),
.B1(n_320),
.B2(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_320),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_324),
.B(n_416),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_348),
.C(n_351),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_325),
.B(n_406),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_329),
.C(n_336),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_326),
.B(n_362),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_329),
.A2(n_330),
.B1(n_336),
.B2(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_336),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_337),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_338),
.B(n_342),
.Y(n_337)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx5_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_343),
.B(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx5_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_348),
.B(n_351),
.Y(n_406)
);

XOR2x2_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_352),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_413),
.B(n_418),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_404),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_364),
.C(n_380),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_368),
.C(n_369),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_374),
.C(n_379),
.Y(n_370)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx3_ASAP7_75t_SL g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_395),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_383),
.B(n_400),
.C(n_409),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_388),
.C(n_394),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_391),
.Y(n_389)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_397),
.B1(n_400),
.B2(n_403),
.Y(n_395)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_396),
.Y(n_409)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_400),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_407),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_405),
.B(n_408),
.C(n_410),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_410),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_415),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_414),
.B(n_415),
.Y(n_418)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);


endmodule