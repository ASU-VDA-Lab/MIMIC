module fake_jpeg_832_n_108 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_108);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_19),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_30),
.Y(n_50)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_44),
.B(n_45),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_43),
.A2(n_36),
.B1(n_37),
.B2(n_31),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_25),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_31),
.B1(n_36),
.B2(n_45),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_49),
.B1(n_39),
.B2(n_45),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_42),
.A2(n_29),
.B1(n_38),
.B2(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_0),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_39),
.B1(n_32),
.B2(n_2),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_55),
.A2(n_52),
.B(n_4),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_28),
.C(n_26),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_3),
.C(n_5),
.Y(n_75)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_58),
.B(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_64),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_53),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_63),
.B1(n_52),
.B2(n_5),
.Y(n_72)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

NOR2x1_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_1),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_72),
.Y(n_76)
);

OAI32xp33_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_46),
.A3(n_54),
.B1(n_51),
.B2(n_53),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_69),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g69 ( 
.A1(n_64),
.A2(n_52),
.B(n_23),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_75),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_77),
.B(n_79),
.Y(n_93)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_69),
.A2(n_59),
.B1(n_21),
.B2(n_16),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_70),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_84),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_6),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_85),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_87),
.B(n_92),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_85),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_6),
.B(n_7),
.Y(n_94)
);

AOI322xp5_ASAP7_75t_SL g98 ( 
.A1(n_94),
.A2(n_95),
.A3(n_82),
.B1(n_76),
.B2(n_10),
.C1(n_11),
.C2(n_8),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_82),
.C(n_78),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_99),
.C(n_90),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_89),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_101),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_93),
.C(n_91),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_96),
.B1(n_99),
.B2(n_97),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_88),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_88),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_12),
.B(n_13),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_106),
.B(n_9),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_11),
.Y(n_108)
);


endmodule