module real_aes_16915_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_756;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g114 ( .A(n_0), .B(n_115), .Y(n_114) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_1), .A2(n_4), .B1(n_254), .B2(n_532), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g148 ( .A1(n_2), .A2(n_41), .B1(n_149), .B2(n_151), .Y(n_148) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_3), .A2(n_22), .B1(n_151), .B2(n_194), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_5), .A2(n_15), .B1(n_176), .B2(n_245), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_6), .A2(n_58), .B1(n_196), .B2(n_221), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_7), .A2(n_16), .B1(n_149), .B2(n_180), .Y(n_610) );
INVx1_ASAP7_75t_L g115 ( .A(n_8), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g593 ( .A(n_9), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_10), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_11), .A2(n_17), .B1(n_178), .B2(n_220), .Y(n_219) );
BUFx2_ASAP7_75t_L g103 ( .A(n_12), .Y(n_103) );
OR2x2_ASAP7_75t_L g122 ( .A(n_12), .B(n_37), .Y(n_122) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_13), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_14), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_18), .A2(n_97), .B1(n_176), .B2(n_254), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_19), .A2(n_38), .B1(n_212), .B2(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_20), .B(n_177), .Y(n_209) );
OAI21x1_ASAP7_75t_L g165 ( .A1(n_21), .A2(n_55), .B(n_166), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_23), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g511 ( .A(n_24), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_25), .B(n_155), .Y(n_518) );
INVx4_ASAP7_75t_R g573 ( .A(n_26), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g156 ( .A1(n_27), .A2(n_45), .B1(n_157), .B2(n_159), .Y(n_156) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_28), .A2(n_51), .B1(n_159), .B2(n_176), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_29), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_30), .B(n_212), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_31), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_32), .B(n_151), .Y(n_525) );
INVx1_ASAP7_75t_L g534 ( .A(n_33), .Y(n_534) );
A2O1A1Ixp33_ASAP7_75t_SL g591 ( .A1(n_34), .A2(n_149), .B(n_161), .C(n_592), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_35), .A2(n_100), .B1(n_116), .B2(n_860), .Y(n_99) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_36), .A2(n_52), .B1(n_149), .B2(n_159), .Y(n_507) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_37), .Y(n_105) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_39), .A2(n_83), .B1(n_149), .B2(n_193), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_40), .A2(n_44), .B1(n_149), .B2(n_180), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g589 ( .A(n_42), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_43), .A2(n_57), .B1(n_176), .B2(n_231), .Y(n_256) );
INVx1_ASAP7_75t_L g522 ( .A(n_46), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_47), .B(n_149), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_48), .Y(n_543) );
INVx2_ASAP7_75t_L g128 ( .A(n_49), .Y(n_128) );
INVx1_ASAP7_75t_L g109 ( .A(n_50), .Y(n_109) );
BUFx3_ASAP7_75t_L g131 ( .A(n_50), .Y(n_131) );
AOI22xp33_ASAP7_75t_L g132 ( .A1(n_53), .A2(n_133), .B1(n_839), .B2(n_840), .Y(n_132) );
INVx1_ASAP7_75t_L g839 ( .A(n_53), .Y(n_839) );
CKINVDCx5p33_ASAP7_75t_R g574 ( .A(n_54), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_56), .A2(n_85), .B1(n_149), .B2(n_159), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_59), .A2(n_72), .B1(n_157), .B2(n_231), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g613 ( .A(n_60), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g179 ( .A1(n_61), .A2(n_74), .B1(n_149), .B2(n_180), .Y(n_179) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_62), .A2(n_95), .B1(n_176), .B2(n_178), .Y(n_175) );
AND2x4_ASAP7_75t_L g145 ( .A(n_63), .B(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g166 ( .A(n_64), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_65), .Y(n_118) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_66), .A2(n_88), .B1(n_157), .B2(n_159), .Y(n_530) );
AO22x1_ASAP7_75t_L g560 ( .A1(n_67), .A2(n_73), .B1(n_242), .B2(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g146 ( .A(n_68), .Y(n_146) );
AND2x2_ASAP7_75t_L g594 ( .A(n_69), .B(n_163), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_70), .B(n_196), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g587 ( .A(n_71), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_75), .B(n_151), .Y(n_544) );
INVx2_ASAP7_75t_L g155 ( .A(n_76), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_77), .B(n_163), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_78), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_79), .A2(n_96), .B1(n_159), .B2(n_196), .Y(n_195) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_80), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_81), .B(n_173), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_82), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g853 ( .A(n_84), .Y(n_853) );
AOI22xp5_ASAP7_75t_L g846 ( .A1(n_86), .A2(n_134), .B1(n_847), .B2(n_848), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_86), .Y(n_847) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_87), .B(n_163), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_89), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_90), .B(n_163), .Y(n_540) );
INVx1_ASAP7_75t_L g113 ( .A(n_91), .Y(n_113) );
NAND2xp33_ASAP7_75t_L g213 ( .A(n_92), .B(n_177), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g568 ( .A1(n_93), .A2(n_182), .B(n_196), .C(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g575 ( .A(n_94), .B(n_576), .Y(n_575) );
NAND2xp33_ASAP7_75t_L g548 ( .A(n_98), .B(n_158), .Y(n_548) );
BUFx12f_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
BUFx6f_ASAP7_75t_L g861 ( .A(n_101), .Y(n_861) );
AND2x6_ASAP7_75t_SL g101 ( .A(n_102), .B(n_106), .Y(n_101) );
NOR2xp33_ASAP7_75t_L g102 ( .A(n_103), .B(n_104), .Y(n_102) );
INVxp33_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
AND3x2_ASAP7_75t_L g120 ( .A(n_108), .B(n_112), .C(n_121), .Y(n_120) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_114), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g493 ( .A(n_113), .Y(n_493) );
OR2x6_ASAP7_75t_L g116 ( .A(n_117), .B(n_123), .Y(n_116) );
INVxp67_ASAP7_75t_SL g849 ( .A(n_117), .Y(n_849) );
NOR2x1_ASAP7_75t_R g117 ( .A(n_118), .B(n_119), .Y(n_117) );
INVx3_ASAP7_75t_L g845 ( .A(n_119), .Y(n_845) );
INVx4_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_121), .B(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NOR2x1_ASAP7_75t_L g859 ( .A(n_122), .B(n_131), .Y(n_859) );
OAI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_132), .B(n_841), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_125), .Y(n_124) );
BUFx12f_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x6_ASAP7_75t_SL g126 ( .A(n_127), .B(n_129), .Y(n_126) );
BUFx3_ASAP7_75t_L g851 ( .A(n_127), .Y(n_851) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g856 ( .A(n_128), .B(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g840 ( .A(n_133), .Y(n_840) );
OA22x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_490), .B1(n_494), .B2(n_496), .Y(n_133) );
INVx2_ASAP7_75t_L g848 ( .A(n_134), .Y(n_848) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_386), .Y(n_134) );
NOR2x1_ASAP7_75t_L g135 ( .A(n_136), .B(n_338), .Y(n_135) );
NAND3xp33_ASAP7_75t_L g136 ( .A(n_137), .B(n_285), .C(n_323), .Y(n_136) );
AOI221xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_216), .B1(n_236), .B2(n_264), .C(n_270), .Y(n_137) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_138), .A2(n_463), .B1(n_466), .B2(n_467), .Y(n_462) );
INVx2_ASAP7_75t_SL g138 ( .A(n_139), .Y(n_138) );
OR2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_187), .Y(n_139) );
INVx1_ASAP7_75t_L g377 ( .A(n_140), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_169), .Y(n_140) );
INVx1_ASAP7_75t_L g329 ( .A(n_141), .Y(n_329) );
AND2x4_ASAP7_75t_L g372 ( .A(n_141), .B(n_293), .Y(n_372) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_L g300 ( .A(n_142), .B(n_203), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_142), .B(n_269), .Y(n_360) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g268 ( .A(n_143), .B(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g284 ( .A(n_143), .B(n_189), .Y(n_284) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_143), .Y(n_291) );
INVx1_ASAP7_75t_L g347 ( .A(n_143), .Y(n_347) );
AO31x2_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_147), .A3(n_162), .B(n_167), .Y(n_143) );
INVx2_ASAP7_75t_L g184 ( .A(n_144), .Y(n_184) );
AO31x2_ASAP7_75t_L g217 ( .A1(n_144), .A2(n_171), .A3(n_218), .B(n_224), .Y(n_217) );
AO31x2_ASAP7_75t_L g239 ( .A1(n_144), .A2(n_190), .A3(n_240), .B(n_247), .Y(n_239) );
AO31x2_ASAP7_75t_L g608 ( .A1(n_144), .A2(n_235), .A3(n_609), .B(n_612), .Y(n_608) );
BUFx10_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g199 ( .A(n_145), .Y(n_199) );
BUFx10_ASAP7_75t_L g509 ( .A(n_145), .Y(n_509) );
INVx1_ASAP7_75t_L g564 ( .A(n_145), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_152), .B1(n_156), .B2(n_160), .Y(n_147) );
INVx1_ASAP7_75t_L g178 ( .A(n_149), .Y(n_178) );
INVx4_ASAP7_75t_L g180 ( .A(n_149), .Y(n_180) );
INVx1_ASAP7_75t_L g231 ( .A(n_149), .Y(n_231) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_150), .Y(n_151) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_150), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_150), .Y(n_159) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_150), .Y(n_177) );
INVx2_ASAP7_75t_L g194 ( .A(n_150), .Y(n_194) );
INVx1_ASAP7_75t_L g196 ( .A(n_150), .Y(n_196) );
INVx1_ASAP7_75t_L g222 ( .A(n_150), .Y(n_222) );
INVx1_ASAP7_75t_L g243 ( .A(n_150), .Y(n_243) );
INVx1_ASAP7_75t_L g246 ( .A(n_150), .Y(n_246) );
INVx1_ASAP7_75t_L g255 ( .A(n_150), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_151), .B(n_587), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g229 ( .A1(n_152), .A2(n_160), .B1(n_230), .B2(n_232), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_152), .A2(n_160), .B1(n_241), .B2(n_244), .Y(n_240) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_152), .A2(n_160), .B1(n_253), .B2(n_256), .Y(n_252) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g508 ( .A(n_153), .Y(n_508) );
BUFx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g546 ( .A(n_154), .Y(n_546) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx8_ASAP7_75t_L g161 ( .A(n_155), .Y(n_161) );
INVx1_ASAP7_75t_L g182 ( .A(n_155), .Y(n_182) );
INVx1_ASAP7_75t_L g521 ( .A(n_155), .Y(n_521) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g212 ( .A(n_158), .Y(n_212) );
OAI22xp33_ASAP7_75t_L g572 ( .A1(n_158), .A2(n_246), .B1(n_573), .B2(n_574), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_159), .B(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g532 ( .A(n_159), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g174 ( .A1(n_160), .A2(n_175), .B1(n_179), .B2(n_181), .Y(n_174) );
OAI22xp5_ASAP7_75t_L g191 ( .A1(n_160), .A2(n_192), .B1(n_195), .B2(n_197), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_160), .A2(n_211), .B(n_213), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_160), .A2(n_181), .B1(n_219), .B2(n_223), .Y(n_218) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_160), .A2(n_506), .B1(n_507), .B2(n_508), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_160), .A2(n_197), .B1(n_530), .B2(n_531), .Y(n_529) );
OAI22x1_ASAP7_75t_L g609 ( .A1(n_160), .A2(n_197), .B1(n_610), .B2(n_611), .Y(n_609) );
INVx6_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
O2A1O1Ixp5_ASAP7_75t_L g207 ( .A1(n_161), .A2(n_180), .B(n_208), .C(n_209), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_161), .A2(n_548), .B(n_549), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_161), .B(n_560), .Y(n_559) );
A2O1A1Ixp33_ASAP7_75t_L g622 ( .A1(n_161), .A2(n_556), .B(n_560), .C(n_563), .Y(n_622) );
AO31x2_ASAP7_75t_L g504 ( .A1(n_162), .A2(n_505), .A3(n_509), .B(n_510), .Y(n_504) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NOR2x1_ASAP7_75t_L g550 ( .A(n_163), .B(n_551), .Y(n_550) );
INVx4_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_164), .B(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_164), .B(n_186), .Y(n_185) );
BUFx3_ASAP7_75t_L g190 ( .A(n_164), .Y(n_190) );
INVx2_ASAP7_75t_SL g205 ( .A(n_164), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_164), .B(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g526 ( .A(n_164), .B(n_509), .Y(n_526) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g173 ( .A(n_165), .Y(n_173) );
INVx3_ASAP7_75t_L g267 ( .A(n_169), .Y(n_267) );
AND2x2_ASAP7_75t_L g282 ( .A(n_169), .B(n_203), .Y(n_282) );
INVx2_ASAP7_75t_L g288 ( .A(n_169), .Y(n_288) );
AND2x4_ASAP7_75t_L g350 ( .A(n_169), .B(n_189), .Y(n_350) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_169), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_169), .B(n_483), .Y(n_482) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g299 ( .A(n_170), .B(n_189), .Y(n_299) );
AND2x2_ASAP7_75t_L g327 ( .A(n_170), .B(n_328), .Y(n_327) );
BUFx2_ASAP7_75t_L g406 ( .A(n_170), .Y(n_406) );
AO31x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_174), .A3(n_183), .B(n_185), .Y(n_170) );
AO31x2_ASAP7_75t_L g528 ( .A1(n_171), .A2(n_198), .A3(n_529), .B(n_533), .Y(n_528) );
AOI21x1_ASAP7_75t_L g583 ( .A1(n_171), .A2(n_584), .B(n_594), .Y(n_583) );
BUFx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_172), .B(n_511), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_172), .B(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g576 ( .A(n_172), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_172), .B(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g201 ( .A(n_173), .Y(n_201) );
INVx2_ASAP7_75t_L g235 ( .A(n_173), .Y(n_235) );
OAI21xp33_ASAP7_75t_L g563 ( .A1(n_173), .A2(n_558), .B(n_564), .Y(n_563) );
INVx3_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVxp67_ASAP7_75t_SL g561 ( .A(n_177), .Y(n_561) );
O2A1O1Ixp33_ASAP7_75t_L g542 ( .A1(n_180), .A2(n_543), .B(n_544), .C(n_545), .Y(n_542) );
INVx1_ASAP7_75t_SL g181 ( .A(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g197 ( .A(n_182), .Y(n_197) );
AO31x2_ASAP7_75t_L g251 ( .A1(n_183), .A2(n_227), .A3(n_252), .B(n_257), .Y(n_251) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_184), .A2(n_568), .B(n_571), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_188), .B(n_203), .Y(n_187) );
INVx1_ASAP7_75t_L g362 ( .A(n_188), .Y(n_362) );
NAND2x1_ASAP7_75t_L g390 ( .A(n_188), .B(n_282), .Y(n_390) );
BUFx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
OR2x2_ASAP7_75t_L g292 ( .A(n_189), .B(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g328 ( .A(n_189), .Y(n_328) );
INVx1_ASAP7_75t_L g404 ( .A(n_189), .Y(n_404) );
AO31x2_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .A3(n_198), .B(n_200), .Y(n_189) );
INVx2_ASAP7_75t_SL g193 ( .A(n_194), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_194), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_197), .B(n_572), .Y(n_571) );
AO31x2_ASAP7_75t_L g226 ( .A1(n_198), .A2(n_227), .A3(n_229), .B(n_233), .Y(n_226) );
INVx2_ASAP7_75t_SL g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_SL g214 ( .A(n_199), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_201), .B(n_202), .Y(n_200) );
NOR2xp33_ASAP7_75t_SL g224 ( .A(n_201), .B(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g228 ( .A(n_201), .Y(n_228) );
AND2x4_ASAP7_75t_L g343 ( .A(n_203), .B(n_328), .Y(n_343) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
BUFx2_ASAP7_75t_L g365 ( .A(n_204), .Y(n_365) );
OAI21x1_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_215), .Y(n_204) );
OAI21x1_ASAP7_75t_L g269 ( .A1(n_205), .A2(n_206), .B(n_215), .Y(n_269) );
OAI21x1_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_210), .B(n_214), .Y(n_206) );
AND2x4_ASAP7_75t_L g237 ( .A(n_216), .B(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_226), .Y(n_216) );
INVx4_ASAP7_75t_SL g261 ( .A(n_217), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_217), .B(n_263), .Y(n_273) );
BUFx2_ASAP7_75t_L g337 ( .A(n_217), .Y(n_337) );
AND2x2_ASAP7_75t_L g381 ( .A(n_217), .B(n_239), .Y(n_381) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_222), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g259 ( .A(n_226), .Y(n_259) );
OR2x2_ASAP7_75t_L g297 ( .A(n_226), .B(n_239), .Y(n_297) );
INVx2_ASAP7_75t_L g308 ( .A(n_226), .Y(n_308) );
AND2x4_ASAP7_75t_L g311 ( .A(n_226), .B(n_312), .Y(n_311) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_226), .Y(n_352) );
INVx1_ASAP7_75t_L g393 ( .A(n_226), .Y(n_393) );
AO21x2_ASAP7_75t_L g566 ( .A1(n_227), .A2(n_567), .B(n_575), .Y(n_566) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_235), .B(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_249), .Y(n_236) );
INVx2_ASAP7_75t_L g486 ( .A(n_237), .Y(n_486) );
AND2x4_ASAP7_75t_L g447 ( .A(n_238), .B(n_250), .Y(n_447) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g263 ( .A(n_239), .Y(n_263) );
INVx2_ASAP7_75t_L g312 ( .A(n_239), .Y(n_312) );
INVx1_ASAP7_75t_L g368 ( .A(n_239), .Y(n_368) );
AND2x2_ASAP7_75t_L g394 ( .A(n_239), .B(n_319), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_239), .B(n_307), .Y(n_398) );
OAI21xp33_ASAP7_75t_SL g517 ( .A1(n_242), .A2(n_518), .B(n_519), .Y(n_517) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_260), .Y(n_249) );
INVx3_ASAP7_75t_L g375 ( .A(n_250), .Y(n_375) );
AND2x4_ASAP7_75t_L g250 ( .A(n_251), .B(n_259), .Y(n_250) );
INVx2_ASAP7_75t_L g279 ( .A(n_251), .Y(n_279) );
INVx2_ASAP7_75t_L g319 ( .A(n_251), .Y(n_319) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_255), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_259), .B(n_261), .Y(n_320) );
AND2x2_ASAP7_75t_L g348 ( .A(n_259), .B(n_319), .Y(n_348) );
INVx1_ASAP7_75t_L g274 ( .A(n_260), .Y(n_274) );
NAND2x1_ASAP7_75t_L g410 ( .A(n_260), .B(n_384), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_260), .B(n_348), .Y(n_459) );
AND2x4_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx2_ASAP7_75t_L g277 ( .A(n_261), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_261), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g367 ( .A(n_261), .B(n_368), .Y(n_367) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_261), .Y(n_444) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_264), .A2(n_457), .B1(n_458), .B2(n_460), .Y(n_456) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_268), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_266), .B(n_300), .Y(n_335) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x4_ASAP7_75t_L g358 ( .A(n_267), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g457 ( .A(n_267), .B(n_268), .Y(n_457) );
AND2x2_ASAP7_75t_L g330 ( .A(n_268), .B(n_299), .Y(n_330) );
AND2x4_ASAP7_75t_L g349 ( .A(n_268), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g400 ( .A(n_268), .B(n_327), .Y(n_400) );
INVx1_ASAP7_75t_L g293 ( .A(n_269), .Y(n_293) );
AOI31xp33_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_274), .A3(n_275), .B(n_280), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_272), .B(n_315), .Y(n_314) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_272), .Y(n_466) );
OAI21xp33_ASAP7_75t_L g484 ( .A1(n_272), .A2(n_274), .B(n_304), .Y(n_484) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g326 ( .A(n_273), .Y(n_326) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g461 ( .A(n_276), .B(n_297), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx2_ASAP7_75t_L g295 ( .A(n_277), .Y(n_295) );
INVx1_ASAP7_75t_L g316 ( .A(n_278), .Y(n_316) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_278), .Y(n_423) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g305 ( .A(n_279), .Y(n_305) );
OR2x2_ASAP7_75t_L g333 ( .A(n_279), .B(n_308), .Y(n_333) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NOR2x1p5_ASAP7_75t_L g322 ( .A(n_284), .B(n_288), .Y(n_322) );
AOI221xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_294), .B1(n_298), .B2(n_301), .C(n_313), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NOR2x1_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g402 ( .A(n_291), .B(n_305), .Y(n_402) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
OR2x2_ASAP7_75t_L g332 ( .A(n_295), .B(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g419 ( .A(n_295), .B(n_311), .Y(n_419) );
AND2x4_ASAP7_75t_L g336 ( .A(n_296), .B(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g355 ( .A(n_297), .B(n_318), .Y(n_355) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
AND2x4_ASAP7_75t_SL g371 ( .A(n_299), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_SL g412 ( .A(n_299), .Y(n_412) );
INVx2_ASAP7_75t_L g421 ( .A(n_299), .Y(n_421) );
AND2x2_ASAP7_75t_L g435 ( .A(n_299), .B(n_365), .Y(n_435) );
INVx1_ASAP7_75t_L g413 ( .A(n_300), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_309), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_306), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_303), .B(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2x1p5_ASAP7_75t_L g345 ( .A(n_304), .B(n_311), .Y(n_345) );
AND2x2_ASAP7_75t_L g366 ( .A(n_304), .B(n_367), .Y(n_366) );
NAND2x1_ASAP7_75t_L g474 ( .A(n_304), .B(n_336), .Y(n_474) );
INVx3_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_317), .B(n_321), .Y(n_313) );
NAND2x1_ASAP7_75t_L g475 ( .A(n_315), .B(n_419), .Y(n_475) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_316), .B(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
INVx4_ASAP7_75t_L g384 ( .A(n_318), .Y(n_384) );
AND2x2_ASAP7_75t_L g454 ( .A(n_318), .B(n_359), .Y(n_454) );
INVx3_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g351 ( .A(n_319), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g364 ( .A(n_322), .B(n_365), .Y(n_364) );
NOR2x1_ASAP7_75t_L g434 ( .A(n_322), .B(n_435), .Y(n_434) );
AOI322xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_327), .A3(n_329), .B1(n_330), .B2(n_331), .C1(n_334), .C2(n_336), .Y(n_323) );
INVxp67_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g417 ( .A(n_327), .B(n_365), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_327), .B(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g441 ( .A(n_327), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g446 ( .A(n_327), .B(n_431), .Y(n_446) );
INVx1_ASAP7_75t_L g455 ( .A(n_327), .Y(n_455) );
OR2x2_ASAP7_75t_L g341 ( .A(n_329), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g468 ( .A(n_329), .Y(n_468) );
AND2x2_ASAP7_75t_L g471 ( .A(n_330), .B(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NOR3xp33_ASAP7_75t_L g407 ( .A(n_333), .B(n_347), .C(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g449 ( .A(n_333), .Y(n_449) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND3xp33_ASAP7_75t_SL g338 ( .A(n_339), .B(n_353), .C(n_363), .Y(n_338) );
AOI222xp33_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_344), .B1(n_346), .B2(n_348), .C1(n_349), .C2(n_351), .Y(n_339) );
INVxp67_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OAI22x1_ASAP7_75t_L g485 ( .A1(n_342), .A2(n_486), .B1(n_487), .B2(n_488), .Y(n_485) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g346 ( .A(n_343), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_343), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g439 ( .A(n_343), .B(n_405), .Y(n_439) );
AND2x4_ASAP7_75t_L g469 ( .A(n_343), .B(n_406), .Y(n_469) );
AND2x2_ASAP7_75t_L g450 ( .A(n_344), .B(n_417), .Y(n_450) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g442 ( .A(n_347), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_348), .B(n_381), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_348), .B(n_367), .Y(n_465) );
INVx1_ASAP7_75t_L g385 ( .A(n_349), .Y(n_385) );
INVx2_ASAP7_75t_L g429 ( .A(n_351), .Y(n_429) );
INVx1_ASAP7_75t_L g379 ( .A(n_352), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2x1p5_ASAP7_75t_L g357 ( .A(n_358), .B(n_361), .Y(n_357) );
AOI221xp5_ASAP7_75t_SL g445 ( .A1(n_358), .A2(n_446), .B1(n_447), .B2(n_448), .C(n_450), .Y(n_445) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g431 ( .A(n_360), .Y(n_431) );
INVxp67_ASAP7_75t_SL g483 ( .A(n_360), .Y(n_483) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_362), .B(n_468), .Y(n_477) );
AOI221xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_366), .B1(n_369), .B2(n_380), .C(n_382), .Y(n_363) );
OR2x2_ASAP7_75t_L g420 ( .A(n_365), .B(n_421), .Y(n_420) );
AOI32xp33_ASAP7_75t_L g401 ( .A1(n_367), .A2(n_381), .A3(n_402), .B1(n_403), .B2(n_407), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_367), .B(n_423), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_373), .B1(n_376), .B2(n_378), .Y(n_369) );
INVx3_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_372), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OR2x2_ASAP7_75t_L g443 ( .A(n_375), .B(n_444), .Y(n_443) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g436 ( .A(n_379), .B(n_381), .Y(n_436) );
AND2x2_ASAP7_75t_L g489 ( .A(n_379), .B(n_394), .Y(n_489) );
AND2x2_ASAP7_75t_L g448 ( .A(n_380), .B(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_381), .B(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .Y(n_382) );
NOR2x1_ASAP7_75t_L g386 ( .A(n_387), .B(n_451), .Y(n_386) );
NAND4xp75_ASAP7_75t_L g387 ( .A(n_388), .B(n_414), .C(n_432), .D(n_445), .Y(n_387) );
AOI211x1_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_391), .B(n_395), .C(n_409), .Y(n_388) );
INVxp67_ASAP7_75t_L g487 ( .A(n_389), .Y(n_487) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_394), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OAI21xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_399), .B(n_401), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
BUFx2_ASAP7_75t_L g408 ( .A(n_404), .Y(n_408) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g480 ( .A(n_408), .Y(n_480) );
NOR3xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .C(n_413), .Y(n_409) );
INVx2_ASAP7_75t_L g472 ( .A(n_410), .Y(n_472) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NOR2x1_ASAP7_75t_L g414 ( .A(n_415), .B(n_424), .Y(n_414) );
OAI22xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_418), .B1(n_420), .B2(n_422), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B1(n_429), .B2(n_430), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AOI21xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_436), .B(n_437), .Y(n_432) );
INVxp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AOI21xp33_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_440), .B(n_443), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_444), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g464 ( .A(n_447), .Y(n_464) );
NAND4xp75_ASAP7_75t_SL g451 ( .A(n_452), .B(n_462), .C(n_470), .D(n_478), .Y(n_451) );
OA21x2_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_455), .B(n_456), .Y(n_452) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
NOR2xp67_ASAP7_75t_SL g470 ( .A(n_471), .B(n_473), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B(n_476), .Y(n_473) );
INVxp67_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
AOI21x1_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_484), .B(n_485), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx8_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx12f_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_493), .Y(n_492) );
BUFx8_ASAP7_75t_SL g495 ( .A(n_493), .Y(n_495) );
AND2x2_ASAP7_75t_L g858 ( .A(n_493), .B(n_859), .Y(n_858) );
INVx3_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x4_ASAP7_75t_L g496 ( .A(n_497), .B(n_729), .Y(n_496) );
NOR4xp25_ASAP7_75t_L g497 ( .A(n_498), .B(n_629), .C(n_671), .D(n_703), .Y(n_497) );
OAI211xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_535), .B(n_577), .C(n_614), .Y(n_498) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x4_ASAP7_75t_L g501 ( .A(n_502), .B(n_512), .Y(n_501) );
INVx2_ASAP7_75t_L g642 ( .A(n_502), .Y(n_642) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g721 ( .A(n_503), .B(n_514), .Y(n_721) );
BUFx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_504), .B(n_528), .Y(n_580) );
AND2x2_ASAP7_75t_L g603 ( .A(n_504), .B(n_604), .Y(n_603) );
INVx2_ASAP7_75t_SL g628 ( .A(n_504), .Y(n_628) );
OR2x2_ASAP7_75t_L g691 ( .A(n_504), .B(n_528), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_508), .A2(n_524), .B(n_525), .Y(n_523) );
OAI21x1_ASAP7_75t_L g556 ( .A1(n_508), .A2(n_557), .B(n_558), .Y(n_556) );
INVx1_ASAP7_75t_L g551 ( .A(n_509), .Y(n_551) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OR2x2_ASAP7_75t_L g625 ( .A(n_513), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g637 ( .A(n_513), .Y(n_637) );
INVxp67_ASAP7_75t_SL g815 ( .A(n_513), .Y(n_815) );
OR2x2_ASAP7_75t_L g828 ( .A(n_513), .B(n_829), .Y(n_828) );
OR2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_527), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_514), .B(n_582), .Y(n_581) );
INVx3_ASAP7_75t_L g601 ( .A(n_514), .Y(n_601) );
AND2x2_ASAP7_75t_L g648 ( .A(n_514), .B(n_649), .Y(n_648) );
NAND2x1p5_ASAP7_75t_SL g667 ( .A(n_514), .B(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_514), .B(n_602), .Y(n_717) );
INVx1_ASAP7_75t_L g806 ( .A(n_514), .Y(n_806) );
AND2x2_ASAP7_75t_L g835 ( .A(n_514), .B(n_528), .Y(n_835) );
AND2x4_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
OAI21xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_523), .B(n_526), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
BUFx4f_ASAP7_75t_L g590 ( .A(n_521), .Y(n_590) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g602 ( .A(n_528), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_528), .B(n_628), .Y(n_650) );
INVx1_ASAP7_75t_L g670 ( .A(n_528), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_528), .B(n_604), .Y(n_722) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_552), .Y(n_536) );
OR2x2_ASAP7_75t_L g619 ( .A(n_537), .B(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g726 ( .A(n_537), .B(n_675), .Y(n_726) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g635 ( .A(n_538), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_538), .B(n_655), .Y(n_654) );
NOR2x1_ASAP7_75t_L g740 ( .A(n_538), .B(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g598 ( .A(n_539), .Y(n_598) );
BUFx3_ASAP7_75t_L g646 ( .A(n_539), .Y(n_646) );
AND2x2_ASAP7_75t_L g682 ( .A(n_539), .B(n_663), .Y(n_682) );
AND2x2_ASAP7_75t_L g762 ( .A(n_539), .B(n_608), .Y(n_762) );
AND2x2_ASAP7_75t_L g775 ( .A(n_539), .B(n_566), .Y(n_775) );
NAND2x1p5_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
OAI21x1_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_547), .B(n_550), .Y(n_541) );
INVx2_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g715 ( .A(n_552), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_552), .B(n_645), .Y(n_723) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_565), .Y(n_552) );
AND2x2_ASAP7_75t_L g634 ( .A(n_553), .B(n_566), .Y(n_634) );
INVx1_ASAP7_75t_L g742 ( .A(n_553), .Y(n_742) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x4_ASAP7_75t_L g596 ( .A(n_554), .B(n_566), .Y(n_596) );
AND2x2_ASAP7_75t_L g659 ( .A(n_554), .B(n_565), .Y(n_659) );
AOI21x1_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_559), .B(n_562), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_564), .A2(n_585), .B(n_591), .Y(n_584) );
AND2x2_ASAP7_75t_L g617 ( .A(n_565), .B(n_608), .Y(n_617) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g607 ( .A(n_566), .B(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g675 ( .A(n_566), .B(n_608), .Y(n_675) );
INVx1_ASAP7_75t_L g686 ( .A(n_566), .Y(n_686) );
AND2x2_ASAP7_75t_L g749 ( .A(n_566), .B(n_598), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_595), .B1(n_599), .B2(n_605), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_578), .A2(n_648), .B1(n_651), .B2(n_653), .Y(n_647) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
OR2x2_ASAP7_75t_L g727 ( .A(n_580), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g833 ( .A(n_580), .Y(n_833) );
INVx1_ASAP7_75t_L g692 ( .A(n_581), .Y(n_692) );
OR2x2_ASAP7_75t_L g755 ( .A(n_581), .B(n_650), .Y(n_755) );
OR2x2_ASAP7_75t_L g626 ( .A(n_582), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_582), .B(n_601), .Y(n_702) );
AND2x2_ASAP7_75t_L g719 ( .A(n_582), .B(n_646), .Y(n_719) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_582), .Y(n_736) );
INVxp67_ASAP7_75t_L g784 ( .A(n_582), .Y(n_784) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g604 ( .A(n_583), .Y(n_604) );
OAI21xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_588), .B(n_590), .Y(n_585) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_596), .Y(n_694) );
INVx3_ASAP7_75t_L g699 ( .A(n_596), .Y(n_699) );
AND2x2_ASAP7_75t_L g712 ( .A(n_596), .B(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g812 ( .A(n_596), .B(n_774), .Y(n_812) );
INVx1_ASAP7_75t_L g606 ( .A(n_597), .Y(n_606) );
OR2x2_ASAP7_75t_L g789 ( .A(n_597), .B(n_764), .Y(n_789) );
BUFx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g713 ( .A(n_598), .B(n_623), .Y(n_713) );
AND2x2_ASAP7_75t_L g734 ( .A(n_598), .B(n_659), .Y(n_734) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_603), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_600), .B(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g735 ( .A(n_600), .Y(n_735) );
AND2x2_ASAP7_75t_L g777 ( .A(n_600), .B(n_778), .Y(n_777) );
AND2x4_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx2_ASAP7_75t_L g678 ( .A(n_601), .Y(n_678) );
AND2x2_ASAP7_75t_L g709 ( .A(n_601), .B(n_710), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_601), .B(n_668), .Y(n_728) );
AND2x2_ASAP7_75t_L g677 ( .A(n_603), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g793 ( .A(n_603), .Y(n_793) );
AND2x2_ASAP7_75t_L g816 ( .A(n_603), .B(n_806), .Y(n_816) );
INVx1_ASAP7_75t_L g829 ( .A(n_603), .Y(n_829) );
INVx2_ASAP7_75t_L g668 ( .A(n_604), .Y(n_668) );
OR2x2_ASAP7_75t_L g764 ( .A(n_604), .B(n_628), .Y(n_764) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_607), .B(n_645), .Y(n_652) );
INVx2_ASAP7_75t_L g623 ( .A(n_608), .Y(n_623) );
INVx2_ASAP7_75t_L g663 ( .A(n_608), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_608), .B(n_621), .Y(n_685) );
OAI21xp33_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_618), .B(n_624), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_617), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OR2x2_ASAP7_75t_L g758 ( .A(n_620), .B(n_759), .Y(n_758) );
OR2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .Y(n_620) );
INVx2_ASAP7_75t_L g664 ( .A(n_621), .Y(n_664) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g655 ( .A(n_623), .Y(n_655) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g638 ( .A(n_626), .Y(n_638) );
INVxp67_ASAP7_75t_L g809 ( .A(n_626), .Y(n_809) );
OR2x2_ASAP7_75t_L g711 ( .A(n_627), .B(n_668), .Y(n_711) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND4xp25_ASAP7_75t_L g629 ( .A(n_630), .B(n_639), .C(n_647), .D(n_656), .Y(n_629) );
NAND3xp33_ASAP7_75t_L g630 ( .A(n_631), .B(n_636), .C(n_638), .Y(n_630) );
INVx3_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
A2O1A1Ixp33_ASAP7_75t_L g825 ( .A1(n_632), .A2(n_826), .B(n_828), .C(n_830), .Y(n_825) );
OR2x6_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_634), .B(n_682), .Y(n_681) );
NOR3xp33_ASAP7_75t_L g737 ( .A(n_634), .B(n_738), .C(n_740), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_634), .B(n_713), .Y(n_818) );
AOI221xp5_ASAP7_75t_L g830 ( .A1(n_634), .A2(n_739), .B1(n_831), .B2(n_834), .C(n_836), .Y(n_830) );
INVx1_ASAP7_75t_L g821 ( .A(n_635), .Y(n_821) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_643), .Y(n_639) );
AOI221xp5_ASAP7_75t_L g756 ( .A1(n_640), .A2(n_648), .B1(n_683), .B2(n_757), .C(n_760), .Y(n_756) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_642), .B(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g707 ( .A(n_643), .Y(n_707) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2x1p5_ASAP7_75t_L g661 ( .A(n_645), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g822 ( .A(n_645), .B(n_673), .Y(n_822) );
INVx3_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
BUFx2_ASAP7_75t_L g658 ( .A(n_646), .Y(n_658) );
AND3x1_ASAP7_75t_L g831 ( .A(n_646), .B(n_832), .C(n_833), .Y(n_831) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g701 ( .A(n_650), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g771 ( .A(n_653), .Y(n_771) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g747 ( .A(n_655), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g774 ( .A(n_655), .Y(n_774) );
OAI21xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_660), .B(n_665), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
NAND2x1_ASAP7_75t_L g672 ( .A(n_658), .B(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g739 ( .A(n_659), .Y(n_739) );
INVxp67_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx1_ASAP7_75t_L g695 ( .A(n_663), .Y(n_695) );
OR2x2_ASAP7_75t_L g674 ( .A(n_664), .B(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g787 ( .A(n_664), .Y(n_787) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_666), .B(n_814), .Y(n_813) );
OR2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_669), .Y(n_666) );
OR2x2_ASAP7_75t_L g743 ( .A(n_667), .B(n_691), .Y(n_743) );
INVx2_ASAP7_75t_L g832 ( .A(n_667), .Y(n_832) );
INVx1_ASAP7_75t_L g706 ( .A(n_668), .Y(n_706) );
NOR4xp25_ASAP7_75t_L g836 ( .A(n_668), .B(n_699), .C(n_837), .D(n_838), .Y(n_836) );
INVx1_ASAP7_75t_L g838 ( .A(n_669), .Y(n_838) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
BUFx3_ASAP7_75t_L g824 ( .A(n_670), .Y(n_824) );
OAI211xp5_ASAP7_75t_SL g671 ( .A1(n_672), .A2(n_676), .B(n_679), .C(n_687), .Y(n_671) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g811 ( .A(n_674), .Y(n_811) );
INVx2_ASAP7_75t_L g796 ( .A(n_675), .Y(n_796) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI21xp5_ASAP7_75t_L g679 ( .A1(n_677), .A2(n_680), .B(n_683), .Y(n_679) );
OR2x2_ASAP7_75t_L g763 ( .A(n_678), .B(n_764), .Y(n_763) );
AND2x2_ASAP7_75t_L g781 ( .A(n_678), .B(n_782), .Y(n_781) );
INVxp67_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g697 ( .A(n_682), .Y(n_697) );
AND2x4_ASAP7_75t_SL g786 ( .A(n_682), .B(n_787), .Y(n_786) );
INVx3_ASAP7_75t_R g683 ( .A(n_684), .Y(n_683) );
OR2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_685), .Y(n_752) );
INVx1_ASAP7_75t_L g759 ( .A(n_686), .Y(n_759) );
AOI32xp33_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_693), .A3(n_695), .B1(n_696), .B2(n_700), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_690), .B(n_692), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_690), .B(n_706), .Y(n_705) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_690), .Y(n_751) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
OR2x2_ASAP7_75t_L g768 ( .A(n_691), .B(n_706), .Y(n_768) );
INVx2_ASAP7_75t_L g782 ( .A(n_691), .Y(n_782) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_SL g761 ( .A(n_699), .B(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
OAI211xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_707), .B(n_708), .C(n_724), .Y(n_703) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_712), .B(n_714), .Y(n_708) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g765 ( .A(n_713), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_713), .B(n_800), .Y(n_799) );
OAI32xp33_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_716), .A3(n_718), .B1(n_720), .B2(n_723), .Y(n_714) );
INVx1_ASAP7_75t_L g800 ( .A(n_715), .Y(n_800) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
OR2x2_ASAP7_75t_L g792 ( .A(n_717), .B(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
INVxp67_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
NOR2x1_ASAP7_75t_L g729 ( .A(n_730), .B(n_801), .Y(n_729) );
NAND4xp25_ASAP7_75t_L g730 ( .A(n_731), .B(n_756), .C(n_769), .D(n_797), .Y(n_730) );
NOR2xp67_ASAP7_75t_L g731 ( .A(n_732), .B(n_744), .Y(n_731) );
OAI32xp33_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_735), .A3(n_736), .B1(n_737), .B2(n_743), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OR2x2_ASAP7_75t_L g783 ( .A(n_735), .B(n_784), .Y(n_783) );
OAI32xp33_ASAP7_75t_L g788 ( .A1(n_735), .A2(n_789), .A3(n_790), .B1(n_792), .B2(n_794), .Y(n_788) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_736), .B(n_824), .Y(n_823) );
NAND2xp5_ASAP7_75t_SL g802 ( .A(n_738), .B(n_803), .Y(n_802) );
INVx3_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g795 ( .A(n_741), .B(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g827 ( .A(n_741), .Y(n_827) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g791 ( .A(n_742), .Y(n_791) );
OAI22x1_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_750), .B1(n_752), .B2(n_753), .Y(n_744) );
INVx2_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_754), .B(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx3_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
NOR2x1_ASAP7_75t_L g820 ( .A(n_758), .B(n_821), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_763), .B1(n_765), .B2(n_766), .Y(n_760) );
NAND2x1_ASAP7_75t_L g826 ( .A(n_762), .B(n_827), .Y(n_826) );
INVx2_ASAP7_75t_L g837 ( .A(n_762), .Y(n_837) );
INVx2_ASAP7_75t_L g778 ( .A(n_764), .Y(n_778) );
INVx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
NOR3xp33_ASAP7_75t_SL g769 ( .A(n_770), .B(n_779), .C(n_788), .Y(n_769) );
AOI21xp5_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_772), .B(n_776), .Y(n_770) );
NAND2xp33_ASAP7_75t_L g798 ( .A(n_772), .B(n_799), .Y(n_798) );
INVx2_ASAP7_75t_SL g772 ( .A(n_773), .Y(n_772) );
AND2x2_ASAP7_75t_L g773 ( .A(n_774), .B(n_775), .Y(n_773) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
AND2x4_ASAP7_75t_L g834 ( .A(n_778), .B(n_835), .Y(n_834) );
AOI21xp5_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_783), .B(n_785), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
AND2x4_ASAP7_75t_L g805 ( .A(n_782), .B(n_806), .Y(n_805) );
INVxp67_ASAP7_75t_SL g804 ( .A(n_784), .Y(n_804) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVxp67_ASAP7_75t_SL g790 ( .A(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
NAND3xp33_ASAP7_75t_SL g801 ( .A(n_802), .B(n_807), .C(n_819), .Y(n_801) );
AND2x2_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .Y(n_803) );
INVx1_ASAP7_75t_L g810 ( .A(n_806), .Y(n_810) );
AOI222xp33_ASAP7_75t_L g807 ( .A1(n_808), .A2(n_811), .B1(n_812), .B2(n_813), .C1(n_816), .C2(n_817), .Y(n_807) );
AND2x2_ASAP7_75t_L g808 ( .A(n_809), .B(n_810), .Y(n_808) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
O2A1O1Ixp5_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_822), .B(n_823), .C(n_825), .Y(n_819) );
AOI21xp5_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_850), .B(n_852), .Y(n_841) );
OAI21xp5_ASAP7_75t_L g842 ( .A1(n_843), .A2(n_846), .B(n_849), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx2_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
NOR2xp33_ASAP7_75t_L g852 ( .A(n_853), .B(n_854), .Y(n_852) );
INVx6_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
BUFx10_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx3_ASAP7_75t_SL g860 ( .A(n_861), .Y(n_860) );
endmodule