module real_jpeg_29133_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_0),
.B(n_25),
.Y(n_24)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_0),
.B(n_68),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_0),
.B(n_89),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_2),
.A2(n_19),
.B1(n_40),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_45),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_3),
.A2(n_19),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_3),
.A2(n_21),
.B1(n_39),
.B2(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_39),
.Y(n_68)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_4),
.A2(n_7),
.B(n_26),
.Y(n_78)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

AOI21xp33_ASAP7_75t_SL g18 ( 
.A1(n_6),
.A2(n_7),
.B(n_19),
.Y(n_18)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_7),
.A2(n_16),
.B1(n_25),
.B2(n_26),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_7),
.A2(n_16),
.B1(n_21),
.B2(n_50),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_7),
.B(n_51),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_7),
.A2(n_16),
.B1(n_19),
.B2(n_40),
.Y(n_76)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_8),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_70),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_69),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_59),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_13),
.B(n_59),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_32),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_22),
.B1(n_23),
.B2(n_31),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_17),
.B(n_18),
.C(n_21),
.Y(n_15)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_16),
.A2(n_19),
.B(n_36),
.C(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_16),
.B(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_16),
.B(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_17),
.A2(n_19),
.B1(n_40),
.B2(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_19),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_19),
.A2(n_36),
.B1(n_37),
.B2(n_40),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

O2A1O1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_21),
.A2(n_51),
.B(n_55),
.C(n_56),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_21),
.B(n_55),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_28),
.B(n_30),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_24),
.B(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_24),
.B(n_30),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_25),
.A2(n_26),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_25),
.B(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_28),
.B(n_30),
.Y(n_66)
);

INVx5_ASAP7_75t_SL g104 ( 
.A(n_28),
.Y(n_104)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_46),
.B1(n_47),
.B2(n_58),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_33),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_41),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_34),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_35),
.B(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_35),
.Y(n_96)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_38),
.B(n_42),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_44),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_53),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_51),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.C(n_65),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_63),
.B1(n_64),
.B2(n_81),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_60),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_82),
.B(n_107),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_79),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_72),
.B(n_79),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_77),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_74),
.B1(n_77),
.B2(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_77),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_93),
.B(n_106),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_91),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_84),
.B(n_91),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

INVxp33_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_99),
.B(n_105),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_95),
.B(n_97),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_102),
.Y(n_99)
);


endmodule