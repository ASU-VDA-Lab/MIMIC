module real_jpeg_1548_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_0),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_0),
.B(n_35),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_0),
.B(n_53),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_0),
.B(n_43),
.Y(n_199)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_4),
.B(n_27),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_4),
.B(n_31),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_4),
.B(n_59),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_4),
.B(n_66),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_4),
.B(n_50),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_4),
.B(n_53),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_4),
.B(n_35),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_4),
.B(n_43),
.Y(n_212)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_5),
.B(n_31),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_5),
.B(n_66),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_5),
.B(n_27),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_5),
.B(n_50),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_8),
.B(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_8),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_8),
.B(n_66),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_8),
.B(n_27),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_8),
.B(n_50),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_8),
.B(n_53),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_9),
.B(n_35),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_9),
.B(n_53),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_9),
.B(n_50),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_9),
.B(n_27),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_9),
.B(n_43),
.Y(n_105)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_12),
.B(n_35),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_12),
.B(n_43),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_12),
.B(n_53),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_14),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_14),
.B(n_50),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_14),
.B(n_27),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_14),
.B(n_43),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_14),
.B(n_66),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g191 ( 
.A(n_14),
.B(n_35),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_147),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_146),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_128),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_20),
.B(n_128),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_81),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_54),
.C(n_71),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_22),
.B(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.C(n_47),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_23),
.A2(n_24),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_29),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_25),
.B(n_33),
.C(n_38),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

INVx3_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_28),
.B(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_28),
.B(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_31),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_36),
.B(n_110),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_39),
.A2(n_40),
.B1(n_47),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_45),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_41),
.A2(n_45),
.B1(n_46),
.B2(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_41),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_44),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_42),
.B(n_57),
.Y(n_215)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_44),
.B(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_45),
.A2(n_46),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_46),
.B(n_97),
.Y(n_140)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_47),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.C(n_52),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_48),
.A2(n_52),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_48),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_49),
.B(n_159),
.Y(n_158)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_52),
.Y(n_160)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_54),
.A2(n_71),
.B1(n_72),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_54),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_63),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_55),
.B(n_64),
.C(n_69),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_61),
.C(n_62),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_56),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_57),
.B(n_70),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_58),
.B(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_61),
.A2(n_62),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_69),
.Y(n_63)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_79),
.B2(n_80),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_77),
.C(n_79),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_77),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_99),
.B2(n_100),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx24_ASAP7_75t_SL g249 ( 
.A(n_83),
.Y(n_249)
);

FAx1_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_93),
.CI(n_94),
.CON(n_83),
.SN(n_83)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_91),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_96),
.B(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_96),
.A2(n_97),
.B1(n_185),
.B2(n_186),
.Y(n_200)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_116),
.B2(n_117),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_111),
.C(n_115),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_144),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_109),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_105),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_107),
.C(n_109),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_105),
.A2(n_108),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_113),
.B(n_114),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_126),
.B2(n_127),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_132),
.C(n_143),
.Y(n_128)
);

FAx1_ASAP7_75t_SL g168 ( 
.A(n_129),
.B(n_132),
.CI(n_143),
.CON(n_168),
.SN(n_168)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.C(n_138),
.Y(n_132)
);

FAx1_ASAP7_75t_SL g152 ( 
.A(n_133),
.B(n_137),
.CI(n_138),
.CON(n_152),
.SN(n_152)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.C(n_142),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_139),
.A2(n_140),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_141),
.B(n_142),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_246),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_169),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_168),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_151),
.B(n_168),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.C(n_157),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_152),
.B(n_243),
.Y(n_242)
);

BUFx24_ASAP7_75t_SL g247 ( 
.A(n_152),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_153),
.B(n_157),
.Y(n_243)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_154),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_162),
.C(n_166),
.Y(n_157)
);

FAx1_ASAP7_75t_SL g233 ( 
.A(n_158),
.B(n_162),
.CI(n_166),
.CON(n_233),
.SN(n_233)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.C(n_165),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_165),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_180),
.Y(n_179)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_168),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_241),
.B(n_245),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_229),
.B(n_240),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_201),
.B(n_228),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_192),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_173),
.B(n_192),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_183),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_175),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.C(n_178),
.Y(n_175)
);

FAx1_ASAP7_75t_SL g193 ( 
.A(n_176),
.B(n_177),
.CI(n_178),
.CON(n_193),
.SN(n_193)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_179),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_179),
.B(n_181),
.C(n_183),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_187),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_184),
.B(n_188),
.C(n_189),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.C(n_200),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_225),
.Y(n_224)
);

BUFx24_ASAP7_75t_SL g251 ( 
.A(n_193),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_194),
.A2(n_195),
.B1(n_200),
.B2(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_222),
.B(n_227),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_213),
.B(n_221),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_209),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_209),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_207),
.C(n_208),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_210),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_216),
.B(n_220),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_218),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_224),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_230),
.B(n_231),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_236),
.C(n_237),
.Y(n_244)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx24_ASAP7_75t_SL g248 ( 
.A(n_233),
.Y(n_248)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_244),
.Y(n_245)
);


endmodule