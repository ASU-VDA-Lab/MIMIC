module fake_jpeg_14422_n_54 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_54);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_54;

wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_18),
.B1(n_17),
.B2(n_14),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_25),
.A2(n_29),
.B1(n_30),
.B2(n_24),
.Y(n_35)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_24),
.B(n_2),
.Y(n_33)
);

OA21x2_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_0),
.B(n_1),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g30 ( 
.A1(n_23),
.A2(n_12),
.B(n_11),
.C(n_10),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_37),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_28),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_36),
.C(n_5),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_34),
.B(n_4),
.Y(n_43)
);

XNOR2x1_ASAP7_75t_SL g44 ( 
.A(n_43),
.B(n_39),
.Y(n_44)
);

BUFx24_ASAP7_75t_SL g49 ( 
.A(n_44),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_36),
.C(n_6),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_46),
.C(n_47),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_49),
.C(n_48),
.Y(n_52)
);

AO21x1_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_7),
.B(n_8),
.Y(n_53)
);

OAI211xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_8),
.B(n_9),
.C(n_48),
.Y(n_54)
);


endmodule