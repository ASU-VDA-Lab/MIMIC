module real_aes_1367_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_783, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_783;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g227 ( .A(n_0), .B(n_164), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_1), .B(n_104), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_2), .B(n_140), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_3), .B(n_162), .Y(n_505) );
INVx1_ASAP7_75t_L g136 ( .A(n_4), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_5), .B(n_140), .Y(n_185) );
NAND2xp33_ASAP7_75t_SL g247 ( .A(n_6), .B(n_146), .Y(n_247) );
INVx1_ASAP7_75t_L g239 ( .A(n_7), .Y(n_239) );
AOI222xp33_ASAP7_75t_SL g100 ( .A1(n_8), .A2(n_101), .B1(n_106), .B2(n_456), .C1(n_463), .C2(n_470), .Y(n_100) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_8), .A2(n_56), .B1(n_448), .B2(n_449), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_8), .Y(n_448) );
CKINVDCx16_ASAP7_75t_R g104 ( .A(n_9), .Y(n_104) );
AND2x2_ASAP7_75t_L g183 ( .A(n_10), .B(n_169), .Y(n_183) );
AND2x2_ASAP7_75t_L g498 ( .A(n_11), .B(n_245), .Y(n_498) );
AND2x2_ASAP7_75t_L g507 ( .A(n_12), .B(n_126), .Y(n_507) );
INVx2_ASAP7_75t_L g128 ( .A(n_13), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_14), .B(n_162), .Y(n_532) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_15), .Y(n_110) );
AOI221x1_ASAP7_75t_L g242 ( .A1(n_16), .A2(n_148), .B1(n_243), .B2(n_245), .C(n_246), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_17), .B(n_140), .Y(n_207) );
OAI22xp5_ASAP7_75t_SL g771 ( .A1(n_18), .A2(n_68), .B1(n_772), .B2(n_773), .Y(n_771) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_18), .Y(n_773) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_19), .B(n_140), .Y(n_547) );
INVx1_ASAP7_75t_L g114 ( .A(n_20), .Y(n_114) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_21), .A2(n_89), .B1(n_131), .B2(n_140), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_22), .A2(n_148), .B(n_187), .Y(n_186) );
AOI221xp5_ASAP7_75t_SL g216 ( .A1(n_23), .A2(n_37), .B1(n_140), .B2(n_148), .C(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_24), .B(n_164), .Y(n_188) );
OA21x2_ASAP7_75t_L g127 ( .A1(n_25), .A2(n_88), .B(n_128), .Y(n_127) );
OR2x2_ASAP7_75t_L g170 ( .A(n_25), .B(n_88), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_26), .B(n_162), .Y(n_211) );
INVxp67_ASAP7_75t_L g241 ( .A(n_27), .Y(n_241) );
AND2x2_ASAP7_75t_L g180 ( .A(n_28), .B(n_168), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_29), .A2(n_148), .B(n_226), .Y(n_225) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_30), .A2(n_245), .B(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_31), .B(n_162), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_32), .A2(n_148), .B(n_503), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_33), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_34), .B(n_162), .Y(n_561) );
AND2x2_ASAP7_75t_L g138 ( .A(n_35), .B(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g146 ( .A(n_35), .B(n_136), .Y(n_146) );
INVx1_ASAP7_75t_L g152 ( .A(n_35), .Y(n_152) );
OR2x6_ASAP7_75t_L g112 ( .A(n_36), .B(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_38), .B(n_140), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g147 ( .A1(n_39), .A2(n_81), .B1(n_148), .B2(n_150), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_40), .B(n_162), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_41), .B(n_140), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_42), .B(n_164), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_43), .A2(n_148), .B(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g230 ( .A(n_44), .B(n_168), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_45), .B(n_164), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_46), .B(n_168), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_47), .B(n_140), .Y(n_529) );
INVx1_ASAP7_75t_L g134 ( .A(n_48), .Y(n_134) );
INVx1_ASAP7_75t_L g143 ( .A(n_48), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_49), .B(n_162), .Y(n_496) );
AND2x2_ASAP7_75t_L g537 ( .A(n_50), .B(n_168), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_51), .B(n_140), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_52), .B(n_164), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_53), .B(n_164), .Y(n_560) );
AND2x2_ASAP7_75t_L g171 ( .A(n_54), .B(n_168), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_55), .B(n_140), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_56), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_57), .B(n_162), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_58), .B(n_140), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_59), .A2(n_148), .B(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_60), .B(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_SL g212 ( .A(n_61), .B(n_169), .Y(n_212) );
AND2x2_ASAP7_75t_L g553 ( .A(n_62), .B(n_169), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_63), .A2(n_148), .B(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_64), .B(n_162), .Y(n_189) );
AND2x2_ASAP7_75t_SL g155 ( .A(n_65), .B(n_126), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_66), .B(n_164), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_67), .B(n_164), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_68), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_69), .Y(n_778) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_70), .A2(n_91), .B1(n_148), .B2(n_150), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_71), .B(n_162), .Y(n_550) );
INVx1_ASAP7_75t_L g139 ( .A(n_72), .Y(n_139) );
INVx1_ASAP7_75t_L g145 ( .A(n_72), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_73), .B(n_164), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_74), .A2(n_148), .B(n_541), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_75), .A2(n_148), .B(n_516), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_76), .A2(n_148), .B(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g563 ( .A(n_77), .B(n_169), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_78), .B(n_168), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g130 ( .A1(n_79), .A2(n_83), .B1(n_131), .B2(n_140), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_80), .B(n_140), .Y(n_166) );
INVx1_ASAP7_75t_L g115 ( .A(n_82), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_84), .B(n_164), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_85), .B(n_164), .Y(n_219) );
AND2x2_ASAP7_75t_L g519 ( .A(n_86), .B(n_126), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_87), .A2(n_148), .B(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_90), .B(n_162), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_92), .A2(n_148), .B(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_93), .B(n_162), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_94), .B(n_140), .Y(n_229) );
INVxp67_ASAP7_75t_L g244 ( .A(n_95), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_96), .B(n_162), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_97), .A2(n_148), .B(n_209), .Y(n_208) );
BUFx2_ASAP7_75t_L g552 ( .A(n_98), .Y(n_552) );
BUFx2_ASAP7_75t_L g105 ( .A(n_99), .Y(n_105) );
BUFx2_ASAP7_75t_SL g460 ( .A(n_99), .Y(n_460) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
OR2x2_ASAP7_75t_SL g102 ( .A(n_103), .B(n_105), .Y(n_102) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_103), .A2(n_458), .B(n_461), .Y(n_457) );
INVx2_ASAP7_75t_L g468 ( .A(n_103), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_105), .B(n_468), .Y(n_467) );
INVxp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_116), .B(n_450), .Y(n_107) );
BUFx2_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
BUFx3_ASAP7_75t_L g455 ( .A(n_109), .Y(n_455) );
BUFx2_ASAP7_75t_L g462 ( .A(n_109), .Y(n_462) );
BUFx2_ASAP7_75t_L g469 ( .A(n_109), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
AND2x6_ASAP7_75t_SL g474 ( .A(n_110), .B(n_112), .Y(n_474) );
OR2x6_ASAP7_75t_SL g770 ( .A(n_110), .B(n_111), .Y(n_770) );
OR2x2_ASAP7_75t_L g781 ( .A(n_110), .B(n_112), .Y(n_781) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
XNOR2x1_ASAP7_75t_L g117 ( .A(n_118), .B(n_447), .Y(n_117) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_118), .A2(n_473), .B1(n_475), .B2(n_768), .Y(n_472) );
AO22x1_ASAP7_75t_L g775 ( .A1(n_118), .A2(n_475), .B1(n_769), .B2(n_776), .Y(n_775) );
AND3x4_ASAP7_75t_L g118 ( .A(n_119), .B(n_318), .C(n_392), .Y(n_118) );
NOR3xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_260), .C(n_291), .Y(n_119) );
A2O1A1Ixp33_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_193), .B(n_202), .C(n_231), .Y(n_120) );
AOI21x1_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_172), .B(n_191), .Y(n_121) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_122), .A2(n_294), .B1(n_300), .B2(n_303), .Y(n_293) );
AND2x2_ASAP7_75t_L g427 ( .A(n_122), .B(n_195), .Y(n_427) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_156), .Y(n_122) );
BUFx2_ASAP7_75t_L g198 ( .A(n_123), .Y(n_198) );
AND2x2_ASAP7_75t_L g286 ( .A(n_123), .B(n_157), .Y(n_286) );
AND2x2_ASAP7_75t_L g357 ( .A(n_123), .B(n_201), .Y(n_357) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_124), .Y(n_251) );
AOI21x1_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_129), .B(n_155), .Y(n_124) );
INVx2_ASAP7_75t_SL g125 ( .A(n_126), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_126), .A2(n_207), .B(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_126), .A2(n_547), .B(n_548), .Y(n_546) );
BUFx4f_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx3_ASAP7_75t_L g223 ( .A(n_127), .Y(n_223) );
AND2x2_ASAP7_75t_SL g169 ( .A(n_128), .B(n_170), .Y(n_169) );
AND2x4_ASAP7_75t_L g190 ( .A(n_128), .B(n_170), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_147), .Y(n_129) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_131), .A2(n_150), .B1(n_238), .B2(n_240), .Y(n_237) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_137), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g149 ( .A(n_134), .B(n_136), .Y(n_149) );
AND2x4_ASAP7_75t_L g162 ( .A(n_134), .B(n_144), .Y(n_162) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x6_ASAP7_75t_L g148 ( .A(n_138), .B(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g154 ( .A(n_139), .Y(n_154) );
AND2x6_ASAP7_75t_L g164 ( .A(n_139), .B(n_142), .Y(n_164) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_146), .Y(n_140) );
INVx1_ASAP7_75t_L g248 ( .A(n_141), .Y(n_248) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx5_ASAP7_75t_L g165 ( .A(n_146), .Y(n_165) );
AND2x4_ASAP7_75t_L g150 ( .A(n_149), .B(n_151), .Y(n_150) );
NOR2x1p5_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x4_ASAP7_75t_L g250 ( .A(n_156), .B(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AND2x2_ASAP7_75t_L g192 ( .A(n_157), .B(n_182), .Y(n_192) );
OR2x2_ASAP7_75t_L g200 ( .A(n_157), .B(n_201), .Y(n_200) );
AND2x4_ASAP7_75t_L g255 ( .A(n_157), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g302 ( .A(n_157), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_157), .B(n_201), .Y(n_310) );
AND2x2_ASAP7_75t_L g347 ( .A(n_157), .B(n_251), .Y(n_347) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_157), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_157), .B(n_181), .Y(n_388) );
AO21x2_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_167), .B(n_171), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_159), .B(n_166), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_163), .B(n_165), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_164), .B(n_552), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_165), .A2(n_177), .B(n_178), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_165), .A2(n_188), .B(n_189), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_165), .A2(n_210), .B(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_165), .A2(n_218), .B(n_219), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_165), .A2(n_227), .B(n_228), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_165), .A2(n_495), .B(n_496), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_165), .A2(n_504), .B(n_505), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_165), .A2(n_517), .B(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_165), .A2(n_532), .B(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_165), .A2(n_542), .B(n_543), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_165), .A2(n_550), .B(n_551), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_165), .A2(n_560), .B(n_561), .Y(n_559) );
AO21x2_ASAP7_75t_L g173 ( .A1(n_167), .A2(n_174), .B(n_180), .Y(n_173) );
AO21x2_ASAP7_75t_L g201 ( .A1(n_167), .A2(n_174), .B(n_180), .Y(n_201) );
AOI21x1_ASAP7_75t_L g500 ( .A1(n_167), .A2(n_501), .B(n_507), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_168), .Y(n_167) );
OA21x2_ASAP7_75t_L g215 ( .A1(n_168), .A2(n_216), .B(n_220), .Y(n_215) );
AO21x2_ASAP7_75t_L g485 ( .A1(n_168), .A2(n_486), .B(n_487), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_168), .A2(n_514), .B(n_515), .Y(n_513) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g289 ( .A(n_172), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_172), .B(n_250), .Y(n_345) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_172), .Y(n_446) );
AND2x4_ASAP7_75t_L g172 ( .A(n_173), .B(n_181), .Y(n_172) );
AND2x2_ASAP7_75t_L g191 ( .A(n_173), .B(n_192), .Y(n_191) );
OR2x2_ASAP7_75t_L g271 ( .A(n_173), .B(n_182), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_173), .B(n_302), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_175), .B(n_179), .Y(n_174) );
AND2x2_ASAP7_75t_L g338 ( .A(n_181), .B(n_255), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_181), .B(n_250), .Y(n_394) );
INVx5_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g196 ( .A(n_182), .Y(n_196) );
AND2x2_ASAP7_75t_L g265 ( .A(n_182), .B(n_256), .Y(n_265) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_182), .Y(n_285) );
AND2x4_ASAP7_75t_L g292 ( .A(n_182), .B(n_201), .Y(n_292) );
AND2x2_ASAP7_75t_SL g439 ( .A(n_182), .B(n_251), .Y(n_439) );
OR2x6_ASAP7_75t_L g182 ( .A(n_183), .B(n_184), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_190), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_190), .B(n_239), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_190), .B(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_190), .B(n_244), .Y(n_243) );
NOR3xp33_ASAP7_75t_L g246 ( .A(n_190), .B(n_247), .C(n_248), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_190), .A2(n_529), .B(n_530), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_190), .A2(n_539), .B(n_540), .Y(n_538) );
INVx1_ASAP7_75t_L g418 ( .A(n_191), .Y(n_418) );
INVx1_ASAP7_75t_L g360 ( .A(n_192), .Y(n_360) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_197), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
OR2x2_ASAP7_75t_L g282 ( .A(n_196), .B(n_200), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_196), .B(n_251), .Y(n_375) );
AND2x2_ASAP7_75t_L g377 ( .A(n_196), .B(n_199), .Y(n_377) );
AOI32xp33_ASAP7_75t_L g443 ( .A1(n_196), .A2(n_259), .A3(n_414), .B1(n_444), .B2(n_446), .Y(n_443) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
AND2x2_ASAP7_75t_L g269 ( .A(n_198), .B(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g387 ( .A(n_198), .B(n_388), .Y(n_387) );
OR2x2_ASAP7_75t_L g410 ( .A(n_198), .B(n_271), .Y(n_410) );
AND2x2_ASAP7_75t_L g437 ( .A(n_198), .B(n_338), .Y(n_437) );
AND2x2_ASAP7_75t_L g363 ( .A(n_199), .B(n_251), .Y(n_363) );
AND2x2_ASAP7_75t_L g438 ( .A(n_199), .B(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g256 ( .A(n_201), .Y(n_256) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_213), .Y(n_203) );
NOR2x1p5_ASAP7_75t_L g296 ( .A(n_204), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g314 ( .A(n_204), .Y(n_314) );
OR2x2_ASAP7_75t_L g342 ( .A(n_204), .B(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x4_ASAP7_75t_SL g259 ( .A(n_205), .B(n_236), .Y(n_259) );
AND2x4_ASAP7_75t_L g275 ( .A(n_205), .B(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g278 ( .A(n_205), .B(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g306 ( .A(n_205), .B(n_215), .Y(n_306) );
OR2x2_ASAP7_75t_L g331 ( .A(n_205), .B(n_280), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_205), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_205), .B(n_215), .Y(n_366) );
INVx2_ASAP7_75t_L g382 ( .A(n_205), .Y(n_382) );
AND2x2_ASAP7_75t_L g397 ( .A(n_205), .B(n_235), .Y(n_397) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_205), .Y(n_421) );
INVx1_ASAP7_75t_L g426 ( .A(n_205), .Y(n_426) );
OR2x6_ASAP7_75t_L g205 ( .A(n_206), .B(n_212), .Y(n_205) );
AND2x2_ASAP7_75t_L g290 ( .A(n_213), .B(n_275), .Y(n_290) );
AND2x2_ASAP7_75t_L g311 ( .A(n_213), .B(n_259), .Y(n_311) );
INVx1_ASAP7_75t_L g343 ( .A(n_213), .Y(n_343) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_221), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g234 ( .A(n_215), .Y(n_234) );
INVx2_ASAP7_75t_L g280 ( .A(n_215), .Y(n_280) );
BUFx3_ASAP7_75t_L g297 ( .A(n_215), .Y(n_297) );
AND2x2_ASAP7_75t_L g336 ( .A(n_215), .B(n_221), .Y(n_336) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_215), .Y(n_434) );
INVx2_ASAP7_75t_L g249 ( .A(n_221), .Y(n_249) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_221), .Y(n_258) );
INVx1_ASAP7_75t_L g274 ( .A(n_221), .Y(n_274) );
OR2x2_ASAP7_75t_L g279 ( .A(n_221), .B(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g299 ( .A(n_221), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_221), .B(n_276), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_221), .B(n_382), .Y(n_381) );
INVx3_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AOI21x1_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_230), .Y(n_222) );
INVx4_ASAP7_75t_L g245 ( .A(n_223), .Y(n_245) );
AO21x2_ASAP7_75t_L g491 ( .A1(n_223), .A2(n_492), .B(n_498), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_229), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_250), .B(n_252), .Y(n_231) );
AND2x2_ASAP7_75t_SL g232 ( .A(n_233), .B(n_235), .Y(n_232) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_233), .Y(n_442) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVxp67_ASAP7_75t_SL g268 ( .A(n_234), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_234), .B(n_274), .Y(n_316) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_234), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_235), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g321 ( .A(n_235), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g372 ( .A(n_235), .Y(n_372) );
AOI221xp5_ASAP7_75t_L g376 ( .A1(n_235), .A2(n_377), .B1(n_378), .B2(n_383), .C(n_386), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_235), .B(n_426), .Y(n_425) );
AND2x4_ASAP7_75t_L g235 ( .A(n_236), .B(n_249), .Y(n_235) );
INVx3_ASAP7_75t_L g276 ( .A(n_236), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_236), .B(n_280), .Y(n_380) );
AND2x2_ASAP7_75t_L g409 ( .A(n_236), .B(n_382), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_236), .B(n_441), .Y(n_440) );
AND2x4_ASAP7_75t_L g236 ( .A(n_237), .B(n_242), .Y(n_236) );
INVx3_ASAP7_75t_L g556 ( .A(n_245), .Y(n_556) );
AND2x2_ASAP7_75t_L g317 ( .A(n_250), .B(n_292), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_250), .A2(n_270), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g254 ( .A(n_251), .B(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g263 ( .A(n_251), .Y(n_263) );
OR2x2_ASAP7_75t_L g309 ( .A(n_251), .B(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_SL g401 ( .A(n_251), .B(n_292), .Y(n_401) );
OR2x2_ASAP7_75t_L g433 ( .A(n_251), .B(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g445 ( .A(n_251), .B(n_351), .Y(n_445) );
INVxp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_257), .Y(n_253) );
INVx2_ASAP7_75t_L g323 ( .A(n_254), .Y(n_323) );
INVx3_ASAP7_75t_SL g389 ( .A(n_255), .Y(n_389) );
INVxp67_ASAP7_75t_L g339 ( .A(n_257), .Y(n_339) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
AOI322xp5_ASAP7_75t_L g261 ( .A1(n_259), .A2(n_262), .A3(n_266), .B1(n_269), .B2(n_272), .C1(n_277), .C2(n_281), .Y(n_261) );
INVx1_ASAP7_75t_SL g350 ( .A(n_259), .Y(n_350) );
AND2x4_ASAP7_75t_L g435 ( .A(n_259), .B(n_322), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_283), .Y(n_260) );
NOR2x1_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
OR2x2_ASAP7_75t_L g288 ( .A(n_263), .B(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g384 ( .A(n_263), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g412 ( .A(n_263), .B(n_265), .Y(n_412) );
AOI32xp33_ASAP7_75t_L g413 ( .A1(n_263), .A2(n_264), .A3(n_414), .B1(n_416), .B2(n_419), .Y(n_413) );
OR2x2_ASAP7_75t_L g417 ( .A(n_263), .B(n_310), .Y(n_417) );
NAND3xp33_ASAP7_75t_L g373 ( .A(n_264), .B(n_289), .C(n_374), .Y(n_373) );
OAI22xp33_ASAP7_75t_SL g393 ( .A1(n_264), .A2(n_330), .B1(n_394), .B2(n_395), .Y(n_393) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVxp67_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g396 ( .A(n_267), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_271), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
OAI322xp33_ASAP7_75t_L g319 ( .A1(n_275), .A2(n_279), .A3(n_288), .B1(n_320), .B2(n_323), .C1(n_324), .C2(n_325), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_275), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_275), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g298 ( .A(n_276), .B(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g330 ( .A(n_276), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_276), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g391 ( .A(n_279), .Y(n_391) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_280), .Y(n_322) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OAI21xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_287), .B(n_290), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_286), .B(n_334), .Y(n_333) );
AOI322xp5_ASAP7_75t_SL g428 ( .A1(n_286), .A2(n_292), .A3(n_409), .B1(n_427), .B2(n_429), .C1(n_432), .C2(n_435), .Y(n_428) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OAI21xp33_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_293), .B(n_307), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_292), .B(n_302), .Y(n_324) );
INVx2_ASAP7_75t_SL g334 ( .A(n_292), .Y(n_334) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
INVx1_ASAP7_75t_SL g359 ( .A(n_298), .Y(n_359) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_299), .Y(n_329) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g404 ( .A(n_305), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g358 ( .A(n_306), .B(n_359), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_311), .B1(n_312), .B2(n_317), .Y(n_307) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NOR4xp75_ASAP7_75t_L g318 ( .A(n_319), .B(n_332), .C(n_352), .D(n_368), .Y(n_318) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
INVxp67_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_SL g326 ( .A(n_327), .B(n_330), .Y(n_326) );
INVxp67_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_330), .A2(n_407), .B1(n_410), .B2(n_411), .Y(n_406) );
OR2x2_ASAP7_75t_L g371 ( .A(n_331), .B(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g415 ( .A(n_331), .Y(n_415) );
OAI221xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_335), .B1(n_337), .B2(n_339), .C(n_340), .Y(n_332) );
INVx2_ASAP7_75t_L g351 ( .A(n_336), .Y(n_351) );
AND2x2_ASAP7_75t_L g408 ( .A(n_336), .B(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_344), .B1(n_346), .B2(n_348), .Y(n_340) );
INVx1_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g403 ( .A(n_347), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_348), .A2(n_354), .B1(n_370), .B2(n_373), .Y(n_369) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
OAI221xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_358), .B1(n_360), .B2(n_361), .C(n_783), .Y(n_352) );
AND2x2_ASAP7_75t_SL g354 ( .A(n_355), .B(n_357), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g420 ( .A(n_359), .B(n_421), .Y(n_420) );
INVxp67_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx1_ASAP7_75t_L g405 ( .A(n_367), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_376), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
AOI21xp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_389), .B(n_390), .Y(n_386) );
NOR3xp33_ASAP7_75t_SL g392 ( .A(n_393), .B(n_398), .C(n_422), .Y(n_392) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_413), .Y(n_398) );
O2A1O1Ixp33_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_402), .B(n_404), .C(n_406), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x4_ASAP7_75t_L g414 ( .A(n_405), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_417), .B(n_418), .Y(n_416) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
NAND4xp25_ASAP7_75t_SL g422 ( .A(n_423), .B(n_428), .C(n_436), .D(n_443), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_427), .Y(n_423) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
INVxp67_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
OAI21xp5_ASAP7_75t_SL g436 ( .A1(n_437), .A2(n_438), .B(n_440), .Y(n_436) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
INVx1_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
BUFx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
CKINVDCx11_ASAP7_75t_R g458 ( .A(n_459), .Y(n_458) );
CKINVDCx8_ASAP7_75t_R g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_469), .Y(n_465) );
INVxp67_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVxp33_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AOI221xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_771), .B1(n_774), .B2(n_775), .C(n_777), .Y(n_471) );
INVx3_ASAP7_75t_SL g776 ( .A(n_473), .Y(n_776) );
CKINVDCx5p33_ASAP7_75t_R g473 ( .A(n_474), .Y(n_473) );
AND2x4_ASAP7_75t_L g475 ( .A(n_476), .B(n_693), .Y(n_475) );
NOR3xp33_ASAP7_75t_L g476 ( .A(n_477), .B(n_629), .C(n_676), .Y(n_476) );
NAND4xp25_ASAP7_75t_SL g477 ( .A(n_478), .B(n_564), .C(n_582), .D(n_608), .Y(n_477) );
OAI21xp33_ASAP7_75t_SL g478 ( .A1(n_479), .A2(n_523), .B(n_524), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_480), .B(n_508), .Y(n_479) );
INVx1_ASAP7_75t_L g744 ( .A(n_480), .Y(n_744) );
OR2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_488), .Y(n_480) );
INVx2_ASAP7_75t_L g568 ( .A(n_481), .Y(n_568) );
AND2x2_ASAP7_75t_L g588 ( .A(n_481), .B(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g690 ( .A(n_481), .B(n_510), .Y(n_690) );
AND2x2_ASAP7_75t_L g750 ( .A(n_481), .B(n_569), .Y(n_750) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_482), .B(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OR2x2_ASAP7_75t_L g634 ( .A(n_483), .B(n_491), .Y(n_634) );
BUFx3_ASAP7_75t_L g644 ( .A(n_483), .Y(n_644) );
AND2x2_ASAP7_75t_L g707 ( .A(n_483), .B(n_708), .Y(n_707) );
AND2x4_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
AND2x4_ASAP7_75t_L g522 ( .A(n_484), .B(n_485), .Y(n_522) );
INVx1_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g753 ( .A(n_489), .Y(n_753) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_499), .Y(n_489) );
AND2x2_ASAP7_75t_L g521 ( .A(n_490), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g708 ( .A(n_490), .Y(n_708) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g523 ( .A(n_491), .B(n_512), .Y(n_523) );
AND2x2_ASAP7_75t_L g585 ( .A(n_491), .B(n_499), .Y(n_585) );
INVx2_ASAP7_75t_L g590 ( .A(n_491), .Y(n_590) );
AND2x2_ASAP7_75t_L g592 ( .A(n_491), .B(n_500), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_497), .Y(n_492) );
INVx1_ASAP7_75t_L g570 ( .A(n_499), .Y(n_570) );
INVx2_ASAP7_75t_L g574 ( .A(n_499), .Y(n_574) );
AND2x4_ASAP7_75t_SL g605 ( .A(n_499), .B(n_512), .Y(n_605) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_499), .Y(n_637) );
INVx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_500), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_506), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_521), .Y(n_508) );
AND2x2_ASAP7_75t_L g671 ( .A(n_509), .B(n_616), .Y(n_671) );
INVx2_ASAP7_75t_SL g759 ( .A(n_509), .Y(n_759) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_520), .Y(n_510) );
NAND2x1p5_ASAP7_75t_L g572 ( .A(n_511), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g679 ( .A(n_511), .B(n_592), .Y(n_679) );
INVx4_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx2_ASAP7_75t_L g567 ( .A(n_512), .Y(n_567) );
AND2x4_ASAP7_75t_L g569 ( .A(n_512), .B(n_570), .Y(n_569) );
NOR2x1_ASAP7_75t_L g589 ( .A(n_512), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g662 ( .A(n_512), .Y(n_662) );
AND2x2_ASAP7_75t_L g681 ( .A(n_512), .B(n_620), .Y(n_681) );
AND2x2_ASAP7_75t_L g712 ( .A(n_512), .B(n_621), .Y(n_712) );
OR2x6_ASAP7_75t_L g512 ( .A(n_513), .B(n_519), .Y(n_512) );
AND2x2_ASAP7_75t_L g651 ( .A(n_521), .B(n_605), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_521), .B(n_662), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_521), .A2(n_762), .B1(n_764), .B2(n_765), .Y(n_761) );
AND2x2_ASAP7_75t_L g764 ( .A(n_521), .B(n_571), .Y(n_764) );
INVx3_ASAP7_75t_L g617 ( .A(n_522), .Y(n_617) );
AND2x2_ASAP7_75t_L g620 ( .A(n_522), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g636 ( .A(n_523), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g645 ( .A(n_523), .Y(n_645) );
AND2x4_ASAP7_75t_SL g524 ( .A(n_525), .B(n_534), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_525), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g696 ( .A(n_525), .B(n_697), .Y(n_696) );
NOR3xp33_ASAP7_75t_L g748 ( .A(n_525), .B(n_658), .C(n_749), .Y(n_748) );
OR2x2_ASAP7_75t_L g766 ( .A(n_525), .B(n_660), .Y(n_766) );
INVx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
OR2x2_ASAP7_75t_L g581 ( .A(n_527), .B(n_545), .Y(n_581) );
INVx1_ASAP7_75t_L g598 ( .A(n_527), .Y(n_598) );
INVx2_ASAP7_75t_L g611 ( .A(n_527), .Y(n_611) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_527), .Y(n_626) );
AND2x2_ASAP7_75t_L g640 ( .A(n_527), .B(n_613), .Y(n_640) );
AND2x2_ASAP7_75t_L g719 ( .A(n_527), .B(n_536), .Y(n_719) );
AOI221xp5_ASAP7_75t_L g582 ( .A1(n_534), .A2(n_583), .B1(n_586), .B2(n_593), .C(n_599), .Y(n_582) );
AOI221xp5_ASAP7_75t_L g711 ( .A1(n_534), .A2(n_712), .B1(n_713), .B2(n_714), .C(n_715), .Y(n_711) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_544), .Y(n_534) );
INVx2_ASAP7_75t_L g653 ( .A(n_535), .Y(n_653) );
AND2x2_ASAP7_75t_L g713 ( .A(n_535), .B(n_597), .Y(n_713) );
AND2x2_ASAP7_75t_L g723 ( .A(n_535), .B(n_609), .Y(n_723) );
OR2x2_ASAP7_75t_L g763 ( .A(n_535), .B(n_647), .Y(n_763) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_SL g580 ( .A(n_536), .B(n_581), .Y(n_580) );
NAND2x1_ASAP7_75t_L g596 ( .A(n_536), .B(n_545), .Y(n_596) );
INVx4_ASAP7_75t_L g625 ( .A(n_536), .Y(n_625) );
OR2x2_ASAP7_75t_L g667 ( .A(n_536), .B(n_554), .Y(n_667) );
OR2x6_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
AND2x2_ASAP7_75t_L g718 ( .A(n_544), .B(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_554), .Y(n_544) );
INVx2_ASAP7_75t_SL g606 ( .A(n_545), .Y(n_606) );
NOR2x1_ASAP7_75t_SL g612 ( .A(n_545), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g627 ( .A(n_545), .B(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g658 ( .A(n_545), .B(n_625), .Y(n_658) );
AND2x2_ASAP7_75t_L g665 ( .A(n_545), .B(n_611), .Y(n_665) );
BUFx2_ASAP7_75t_L g699 ( .A(n_545), .Y(n_699) );
AND2x2_ASAP7_75t_L g710 ( .A(n_545), .B(n_625), .Y(n_710) );
OR2x6_ASAP7_75t_L g545 ( .A(n_546), .B(n_553), .Y(n_545) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_554), .Y(n_578) );
AND2x2_ASAP7_75t_L g597 ( .A(n_554), .B(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g628 ( .A(n_554), .Y(n_628) );
AND2x2_ASAP7_75t_L g654 ( .A(n_554), .B(n_610), .Y(n_654) );
INVx3_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AO21x2_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B(n_563), .Y(n_555) );
AO21x1_ASAP7_75t_SL g613 ( .A1(n_556), .A2(n_557), .B(n_563), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_562), .Y(n_557) );
OAI31xp33_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_569), .A3(n_571), .B(n_575), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx2_ASAP7_75t_L g673 ( .A(n_567), .Y(n_673) );
NOR2xp67_ASAP7_75t_L g583 ( .A(n_568), .B(n_584), .Y(n_583) );
AOI322xp5_ASAP7_75t_L g663 ( .A1(n_568), .A2(n_657), .A3(n_664), .B1(n_668), .B2(n_669), .C1(n_671), .C2(n_672), .Y(n_663) );
AND2x2_ASAP7_75t_L g735 ( .A(n_568), .B(n_712), .Y(n_735) );
AOI221xp5_ASAP7_75t_SL g648 ( .A1(n_569), .A2(n_649), .B1(n_651), .B2(n_652), .C(n_655), .Y(n_648) );
INVx2_ASAP7_75t_L g668 ( .A(n_569), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_571), .B(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_571), .B(n_664), .Y(n_767) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OR2x2_ASAP7_75t_L g642 ( .A(n_572), .B(n_617), .Y(n_642) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g621 ( .A(n_574), .B(n_590), .Y(n_621) );
AND2x4_ASAP7_75t_L g575 ( .A(n_576), .B(n_579), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g692 ( .A(n_578), .Y(n_692) );
O2A1O1Ixp5_ASAP7_75t_L g683 ( .A1(n_579), .A2(n_684), .B(n_686), .C(n_688), .Y(n_683) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_580), .A2(n_716), .B1(n_717), .B2(n_720), .Y(n_715) );
OR2x2_ASAP7_75t_L g670 ( .A(n_581), .B(n_667), .Y(n_670) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_587), .B(n_591), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g603 ( .A(n_590), .Y(n_603) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_592), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .Y(n_594) );
INVx3_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g646 ( .A(n_596), .B(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_596), .B(n_597), .Y(n_689) );
OR2x2_ASAP7_75t_L g691 ( .A(n_596), .B(n_692), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_596), .B(n_740), .Y(n_739) );
BUFx2_ASAP7_75t_L g607 ( .A(n_598), .Y(n_607) );
NOR4xp25_ASAP7_75t_L g599 ( .A(n_600), .B(n_604), .C(n_606), .D(n_607), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g727 ( .A(n_601), .B(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g755 ( .A(n_601), .B(n_604), .Y(n_755) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g685 ( .A(n_603), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_604), .B(n_633), .Y(n_720) );
AOI321xp33_ASAP7_75t_L g722 ( .A1(n_604), .A2(n_723), .A3(n_724), .B1(n_725), .B2(n_727), .C(n_730), .Y(n_722) );
INVx2_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_SL g684 ( .A(n_605), .B(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_605), .B(n_644), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_606), .B(n_628), .Y(n_733) );
OR2x2_ASAP7_75t_L g760 ( .A(n_607), .B(n_644), .Y(n_760) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_614), .B(n_618), .Y(n_608) );
AND2x2_ASAP7_75t_L g649 ( .A(n_609), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_612), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g675 ( .A(n_611), .B(n_613), .Y(n_675) );
INVx2_ASAP7_75t_L g660 ( .A(n_612), .Y(n_660) );
INVx1_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_615), .B(n_731), .Y(n_730) );
OR2x2_ASAP7_75t_L g716 ( .A(n_616), .B(n_668), .Y(n_716) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g674 ( .A(n_617), .B(n_675), .Y(n_674) );
NOR2x1_ASAP7_75t_L g752 ( .A(n_617), .B(n_753), .Y(n_752) );
NOR2xp67_ASAP7_75t_L g618 ( .A(n_619), .B(n_622), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g703 ( .A(n_621), .Y(n_703) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_627), .Y(n_623) );
NOR2xp67_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_625), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g650 ( .A(n_625), .Y(n_650) );
BUFx2_ASAP7_75t_L g732 ( .A(n_625), .Y(n_732) );
INVxp67_ASAP7_75t_L g740 ( .A(n_628), .Y(n_740) );
NAND3xp33_ASAP7_75t_L g629 ( .A(n_630), .B(n_648), .C(n_663), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_638), .B(n_641), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_635), .Y(n_631) );
INVx2_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
OR2x2_ASAP7_75t_L g661 ( .A(n_634), .B(n_662), .Y(n_661) );
INVx2_ASAP7_75t_L g714 ( .A(n_635), .Y(n_714) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g729 ( .A(n_637), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_638), .A2(n_735), .B(n_736), .Y(n_734) );
INVx1_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
INVx2_ASAP7_75t_SL g647 ( .A(n_640), .Y(n_647) );
AND2x2_ASAP7_75t_L g709 ( .A(n_640), .B(n_710), .Y(n_709) );
AOI21xp33_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_643), .B(n_646), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_642), .A2(n_689), .B1(n_690), .B2(n_691), .Y(n_688) );
OR2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
INVx1_ASAP7_75t_L g678 ( .A(n_644), .Y(n_678) );
OR2x2_ASAP7_75t_L g726 ( .A(n_647), .B(n_658), .Y(n_726) );
NOR4xp25_ASAP7_75t_L g758 ( .A(n_650), .B(n_699), .C(n_759), .D(n_760), .Y(n_758) );
AND2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
OR2x2_ASAP7_75t_L g659 ( .A(n_653), .B(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_653), .B(n_675), .Y(n_757) );
AOI21xp33_ASAP7_75t_SL g655 ( .A1(n_656), .A2(n_659), .B(n_661), .Y(n_655) );
INVx2_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
OR2x2_ASAP7_75t_L g746 ( .A(n_658), .B(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g754 ( .A(n_660), .Y(n_754) );
AND2x4_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
INVxp67_ASAP7_75t_L g682 ( .A(n_665), .Y(n_682) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
OR2x2_ASAP7_75t_L g698 ( .A(n_667), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
AND2x2_ASAP7_75t_L g701 ( .A(n_673), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g747 ( .A(n_675), .Y(n_747) );
A2O1A1Ixp33_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_680), .B(n_682), .C(n_683), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
INVx1_ASAP7_75t_L g737 ( .A(n_679), .Y(n_737) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVxp67_ASAP7_75t_L g741 ( .A(n_684), .Y(n_741) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NOR3xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_721), .C(n_742), .Y(n_693) );
OAI211xp5_ASAP7_75t_SL g694 ( .A1(n_695), .A2(n_700), .B(n_704), .C(n_711), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
INVxp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
OAI21xp5_ASAP7_75t_SL g704 ( .A1(n_705), .A2(n_707), .B(n_709), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
O2A1O1Ixp33_ASAP7_75t_L g743 ( .A1(n_707), .A2(n_744), .B(n_745), .C(n_748), .Y(n_743) );
BUFx2_ASAP7_75t_L g724 ( .A(n_708), .Y(n_724) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_734), .Y(n_721) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_731), .A2(n_737), .B1(n_738), .B2(n_741), .Y(n_736) );
OR2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
NAND4xp25_ASAP7_75t_L g742 ( .A(n_743), .B(n_751), .C(n_761), .D(n_767), .Y(n_742) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
AOI221xp5_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_754), .B1(n_755), .B2(n_756), .C(n_758), .Y(n_751) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
CKINVDCx11_ASAP7_75t_R g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g774 ( .A(n_771), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g777 ( .A(n_778), .B(n_779), .Y(n_777) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx3_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
endmodule