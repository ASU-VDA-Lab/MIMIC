module fake_jpeg_28538_n_141 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_141);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_34),
.Y(n_42)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

BUFx2_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_36),
.A2(n_26),
.B1(n_13),
.B2(n_18),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_45),
.B1(n_53),
.B2(n_15),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_20),
.C(n_13),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_48),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_20),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_49),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_22),
.B1(n_24),
.B2(n_21),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_18),
.B(n_16),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_16),
.Y(n_49)
);

OAI21xp33_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_28),
.B(n_21),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_17),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_31),
.A2(n_25),
.B1(n_19),
.B2(n_28),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_50),
.A2(n_25),
.B1(n_15),
.B2(n_14),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_55),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_30),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_63),
.Y(n_85)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_47),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_59),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_30),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_60),
.B(n_73),
.Y(n_82)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_67),
.Y(n_79)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_17),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_68),
.B(n_74),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_72),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_34),
.B1(n_14),
.B2(n_16),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_4),
.B1(n_7),
.B2(n_9),
.Y(n_87)
);

INVxp33_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_41),
.B(n_16),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_9),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_16),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_7),
.Y(n_76)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_0),
.B(n_1),
.C(n_4),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_80),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_60),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_63),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_86),
.A2(n_87),
.B1(n_54),
.B2(n_75),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_81),
.A2(n_65),
.B(n_58),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_101),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_70),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_94),
.B(n_96),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_65),
.B(n_58),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_95),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_56),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_97),
.Y(n_110)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_99),
.B(n_104),
.Y(n_113)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_59),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_78),
.A2(n_59),
.B(n_72),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_103),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_61),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_77),
.B(n_92),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_92),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_112),
.B(n_114),
.Y(n_116)
);

NOR4xp25_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_88),
.C(n_80),
.D(n_84),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_113),
.A2(n_83),
.B1(n_99),
.B2(n_95),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_117),
.A2(n_122),
.B1(n_123),
.B2(n_91),
.Y(n_126)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_118),
.A2(n_119),
.B(n_120),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_77),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

FAx1_ASAP7_75t_SL g121 ( 
.A(n_111),
.B(n_96),
.CI(n_94),
.CON(n_121),
.SN(n_121)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_111),
.C(n_101),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_102),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_109),
.A2(n_103),
.B1(n_102),
.B2(n_83),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_SL g124 ( 
.A1(n_123),
.A2(n_108),
.B(n_83),
.C(n_93),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_124),
.A2(n_117),
.B(n_120),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_126),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_82),
.B1(n_115),
.B2(n_110),
.Y(n_127)
);

FAx1_ASAP7_75t_SL g130 ( 
.A(n_127),
.B(n_128),
.CI(n_122),
.CON(n_130),
.SN(n_130)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_118),
.A2(n_115),
.B1(n_98),
.B2(n_87),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_124),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_132),
.A2(n_124),
.B(n_121),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_129),
.A2(n_121),
.B(n_79),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_133),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_136),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_134),
.A2(n_132),
.B(n_131),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_137),
.B(n_10),
.Y(n_139)
);

AOI322xp5_ASAP7_75t_SL g140 ( 
.A1(n_139),
.A2(n_10),
.A3(n_11),
.B1(n_138),
.B2(n_97),
.C1(n_89),
.C2(n_67),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_11),
.Y(n_141)
);


endmodule