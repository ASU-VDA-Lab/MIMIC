module fake_jpeg_23850_n_173 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_173);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx5p33_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_16),
.B(n_0),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_22),
.B1(n_15),
.B2(n_20),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_40),
.B1(n_35),
.B2(n_19),
.Y(n_62)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_54),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_32),
.A2(n_15),
.B1(n_22),
.B2(n_27),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_35),
.B1(n_28),
.B2(n_30),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_33),
.B(n_19),
.Y(n_49)
);

OAI21xp33_ASAP7_75t_L g75 ( 
.A1(n_49),
.A2(n_55),
.B(n_3),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_23),
.B1(n_29),
.B2(n_20),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_56),
.B1(n_27),
.B2(n_17),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_16),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g55 ( 
.A1(n_33),
.A2(n_0),
.B(n_2),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_23),
.B1(n_29),
.B2(n_17),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_60),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_26),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_59),
.B(n_63),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_57),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_50),
.B1(n_47),
.B2(n_44),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_30),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_69),
.B(n_28),
.Y(n_79)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_66),
.Y(n_93)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_53),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_45),
.B(n_2),
.Y(n_68)
);

OAI21xp33_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_72),
.B(n_75),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_30),
.B1(n_26),
.B2(n_4),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_26),
.B(n_31),
.C(n_34),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_70),
.B(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_R g72 ( 
.A(n_54),
.B(n_28),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_2),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_3),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_14),
.Y(n_74)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_86),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_84),
.B1(n_47),
.B2(n_50),
.Y(n_101)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_80),
.B(n_91),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_73),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_43),
.C(n_48),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_85),
.C(n_79),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_43),
.C(n_44),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_52),
.B(n_44),
.Y(n_87)
);

NOR3xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_58),
.C(n_61),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_89),
.Y(n_97)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_63),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_99),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_87),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_85),
.C(n_83),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_71),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_108),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_101),
.A2(n_107),
.B1(n_43),
.B2(n_53),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_72),
.Y(n_104)
);

A2O1A1O1Ixp25_ASAP7_75t_L g122 ( 
.A1(n_104),
.A2(n_81),
.B(n_73),
.C(n_89),
.D(n_53),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_105),
.A2(n_107),
.B(n_88),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_98),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_50),
.B1(n_47),
.B2(n_52),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_110),
.B(n_108),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_115),
.B(n_122),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_113),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_100),
.A2(n_78),
.B1(n_110),
.B2(n_92),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_119),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_91),
.B1(n_84),
.B2(n_93),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_118),
.A2(n_103),
.B1(n_99),
.B2(n_104),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_103),
.B(n_93),
.Y(n_119)
);

OAI32xp33_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_81),
.A3(n_73),
.B1(n_68),
.B2(n_89),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_123),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_90),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_95),
.B(n_77),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_125),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_53),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_123),
.Y(n_130)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_131),
.A2(n_132),
.B1(n_135),
.B2(n_137),
.Y(n_143)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_111),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_13),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_113),
.C(n_122),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_142),
.C(n_144),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_136),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_141),
.A2(n_147),
.B(n_127),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_112),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_99),
.C(n_102),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_97),
.C(n_21),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_128),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_13),
.C(n_5),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_4),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_141),
.B(n_128),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_153),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_146),
.A2(n_137),
.B1(n_133),
.B2(n_132),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_150),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_143),
.A2(n_127),
.B(n_129),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_154),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_155),
.B(n_154),
.Y(n_159)
);

OAI21x1_ASAP7_75t_L g157 ( 
.A1(n_152),
.A2(n_139),
.B(n_142),
.Y(n_157)
);

AOI21x1_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_7),
.B(n_9),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_159),
.B(n_7),
.Y(n_164)
);

A2O1A1O1Ixp25_ASAP7_75t_L g160 ( 
.A1(n_151),
.A2(n_4),
.B(n_6),
.C(n_7),
.D(n_8),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_160),
.A2(n_12),
.B(n_10),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_151),
.C(n_9),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_162),
.A2(n_163),
.B(n_10),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_11),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_166),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_156),
.A2(n_10),
.B1(n_11),
.B2(n_159),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_168),
.Y(n_171)
);

INVxp33_ASAP7_75t_L g170 ( 
.A(n_169),
.Y(n_170)
);

AO21x1_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_162),
.B(n_158),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_170),
.Y(n_173)
);


endmodule