module fake_netlist_1_5846_n_30 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_30);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NAND2xp5_ASAP7_75t_L g14 ( .A(n_2), .B(n_5), .Y(n_14) );
BUFx6f_ASAP7_75t_L g15 ( .A(n_2), .Y(n_15) );
AND2x4_ASAP7_75t_L g16 ( .A(n_3), .B(n_8), .Y(n_16) );
AND3x2_ASAP7_75t_L g17 ( .A(n_11), .B(n_0), .C(n_3), .Y(n_17) );
AND2x4_ASAP7_75t_L g18 ( .A(n_9), .B(n_1), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_1), .B(n_7), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_16), .Y(n_20) );
AOI22xp33_ASAP7_75t_L g21 ( .A1(n_16), .A2(n_0), .B1(n_4), .B2(n_6), .Y(n_21) );
OAI21x1_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_19), .B(n_14), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
AND2x4_ASAP7_75t_L g24 ( .A(n_23), .B(n_20), .Y(n_24) );
OAI33xp33_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_20), .A3(n_22), .B1(n_17), .B2(n_15), .B3(n_18), .Y(n_25) );
XOR2x2_ASAP7_75t_L g26 ( .A(n_25), .B(n_24), .Y(n_26) );
NAND3xp33_ASAP7_75t_SL g27 ( .A(n_26), .B(n_18), .C(n_15), .Y(n_27) );
HB1xp67_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_28), .B(n_15), .Y(n_29) );
AOI22x1_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_10), .B1(n_12), .B2(n_13), .Y(n_30) );
endmodule