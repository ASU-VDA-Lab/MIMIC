module real_jpeg_5453_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_1),
.B(n_226),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_1),
.B(n_259),
.C(n_262),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_L g264 ( 
.A1(n_1),
.A2(n_71),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_1),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_1),
.B(n_140),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_1),
.A2(n_24),
.B1(n_302),
.B2(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_1),
.B(n_192),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_1),
.A2(n_225),
.B(n_390),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_2),
.A2(n_73),
.B1(n_77),
.B2(n_78),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_2),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_2),
.A2(n_77),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_2),
.A2(n_77),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_3),
.A2(n_115),
.B1(n_117),
.B2(n_118),
.Y(n_114)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_3),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_3),
.A2(n_117),
.B1(n_152),
.B2(n_154),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_3),
.A2(n_101),
.B1(n_117),
.B2(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_3),
.A2(n_71),
.B1(n_117),
.B2(n_335),
.Y(n_374)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_5),
.A2(n_101),
.B1(n_103),
.B2(n_104),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_5),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_5),
.A2(n_103),
.B1(n_277),
.B2(n_279),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_5),
.A2(n_103),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_5),
.A2(n_103),
.B1(n_142),
.B2(n_220),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_6),
.A2(n_25),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_6),
.A2(n_45),
.B1(n_69),
.B2(n_71),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_6),
.A2(n_45),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_7),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_7),
.A2(n_35),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_8),
.Y(n_150)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_8),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_8),
.Y(n_237)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_9),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_10),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_10),
.Y(n_92)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_10),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_10),
.Y(n_99)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_10),
.Y(n_223)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_11),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_12),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_12),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_12),
.A2(n_109),
.B1(n_204),
.B2(n_208),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_12),
.A2(n_26),
.B1(n_109),
.B2(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_12),
.A2(n_109),
.B1(n_163),
.B2(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_13),
.Y(n_86)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_13),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_13),
.Y(n_102)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_13),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_13),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_13),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_13),
.Y(n_216)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_13),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_14),
.A2(n_101),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_14),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_14),
.A2(n_163),
.B1(n_241),
.B2(n_268),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_14),
.A2(n_241),
.B1(n_303),
.B2(n_305),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_14),
.A2(n_185),
.B1(n_241),
.B2(n_343),
.Y(n_342)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_15),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_246),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_244),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_196),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_19),
.B(n_196),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_145),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_81),
.C(n_112),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_22),
.B(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_50),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_23),
.B(n_50),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_31),
.B(n_39),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_24),
.A2(n_149),
.B(n_151),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_24),
.B(n_44),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_24),
.A2(n_31),
.B1(n_228),
.B2(n_234),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_24),
.A2(n_173),
.B(n_284),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_24),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_24),
.A2(n_41),
.B1(n_290),
.B2(n_302),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_24),
.A2(n_39),
.B(n_151),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_29),
.Y(n_24)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_25),
.Y(n_230)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_28),
.Y(n_158)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_30),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_30),
.Y(n_364)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_34),
.Y(n_153)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_36),
.Y(n_291)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_37),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_42),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_67),
.B1(n_72),
.B2(n_79),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_51),
.A2(n_160),
.B(n_166),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_51),
.A2(n_371),
.B(n_372),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_51),
.A2(n_166),
.B(n_374),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_52),
.A2(n_80),
.B1(n_161),
.B2(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_52),
.A2(n_80),
.B1(n_264),
.B2(n_267),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_52),
.A2(n_80),
.B1(n_267),
.B2(n_276),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_52),
.A2(n_80),
.B1(n_276),
.B2(n_347),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_62),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_57),
.B1(n_58),
.B2(n_61),
.Y(n_53)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_54),
.Y(n_281)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_55),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_55),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_55),
.Y(n_278)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g336 ( 
.A(n_56),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_58),
.B1(n_63),
.B2(n_65),
.Y(n_62)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_63),
.Y(n_262)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_68),
.B(n_80),
.Y(n_166)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_72),
.Y(n_179)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_73),
.Y(n_348)
);

INVx5_ASAP7_75t_SL g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_75),
.Y(n_257)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g123 ( 
.A1(n_76),
.A2(n_124),
.B1(n_127),
.B2(n_128),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_76),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_79),
.B(n_265),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_79),
.B(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_81),
.A2(n_82),
.B1(n_112),
.B2(n_113),
.Y(n_198)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_100),
.B1(n_106),
.B2(n_111),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_83),
.A2(n_106),
.B(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_83),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_83),
.A2(n_111),
.B1(n_389),
.B2(n_393),
.Y(n_388)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_93),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_93)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_94),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_95),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g341 ( 
.A(n_95),
.Y(n_341)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g207 ( 
.A(n_96),
.Y(n_207)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_96),
.Y(n_345)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_98),
.Y(n_208)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_98),
.Y(n_331)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_99),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_100),
.Y(n_243)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_105),
.Y(n_191)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_110),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_111),
.Y(n_192)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_121),
.B(n_139),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_114),
.B(n_123),
.Y(n_209)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_121),
.A2(n_123),
.B1(n_356),
.B2(n_357),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_121),
.A2(n_123),
.B1(n_357),
.B2(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_122),
.B(n_141),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_122),
.A2(n_203),
.B(n_209),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_122),
.A2(n_140),
.B1(n_340),
.B2(n_342),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_129),
.Y(n_122)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_123),
.A2(n_182),
.B(n_186),
.Y(n_181)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_124),
.Y(n_333)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_126),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_126),
.Y(n_327)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_132),
.B1(n_134),
.B2(n_137),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_134),
.Y(n_183)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_142),
.Y(n_220)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_168),
.B1(n_194),
.B2(n_195),
.Y(n_145)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_159),
.B2(n_167),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

INVx3_ASAP7_75t_SL g152 ( 
.A(n_153),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_157),
.Y(n_304)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_158),
.Y(n_233)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_158),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_159),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_180),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_177),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_170),
.A2(n_177),
.B1(n_178),
.B2(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_172),
.A2(n_229),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

INVx5_ASAP7_75t_L g310 ( 
.A(n_175),
.Y(n_310)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_187),
.B1(n_188),
.B2(n_193),
.Y(n_180)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_192),
.A2(n_239),
.B1(n_242),
.B2(n_243),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.C(n_201),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_197),
.B(n_199),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_201),
.B(n_403),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_210),
.C(n_238),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_202),
.B(n_238),
.Y(n_399)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_203),
.Y(n_386)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

OAI32xp33_ASAP7_75t_L g322 ( 
.A1(n_208),
.A2(n_323),
.A3(n_325),
.B1(n_328),
.B2(n_332),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_210),
.B(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_227),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_211),
.B(n_227),
.Y(n_382)
);

OAI32xp33_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_215),
.A3(n_217),
.B1(n_219),
.B2(n_224),
.Y(n_211)
);

INVx4_ASAP7_75t_SL g212 ( 
.A(n_213),
.Y(n_212)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVxp33_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_232),
.Y(n_285)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_235),
.Y(n_234)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_239),
.Y(n_393)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_395),
.B(n_408),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_378),
.B(n_394),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_350),
.B(n_377),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_318),
.B(n_349),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_286),
.B(n_317),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_271),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_253),
.B(n_271),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_263),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_254),
.B(n_263),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_265),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_265),
.B(n_329),
.Y(n_328)
);

OAI21xp33_ASAP7_75t_SL g340 ( 
.A1(n_265),
.A2(n_328),
.B(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_270),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_283),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_275),
.B2(n_282),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_273),
.B(n_282),
.C(n_283),
.Y(n_319)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_275),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_284),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_298),
.B(n_316),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_297),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_297),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_289),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_291),
.B(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_299),
.A2(n_308),
.B(n_315),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_300),
.B(n_301),
.Y(n_315)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx4_ASAP7_75t_SL g305 ( 
.A(n_306),
.Y(n_305)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_311),
.Y(n_308)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_319),
.B(n_320),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_338),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_321),
.B(n_339),
.C(n_346),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_337),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_322),
.B(n_337),
.Y(n_369)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx6_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx5_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_346),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_342),
.Y(n_356)
);

INVx5_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx6_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_347),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_351),
.B(n_352),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_353),
.A2(n_354),
.B1(n_367),
.B2(n_368),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_353),
.B(n_370),
.C(n_375),
.Y(n_379)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_355),
.B(n_358),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_355),
.B(n_359),
.C(n_366),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_359),
.A2(n_360),
.B1(n_365),
.B2(n_366),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx8_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_365),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_369),
.A2(n_370),
.B1(n_375),
.B2(n_376),
.Y(n_368)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_369),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_370),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_379),
.B(n_380),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_384),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_383),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_382),
.B(n_383),
.C(n_384),
.Y(n_405)
);

BUFx24_ASAP7_75t_SL g411 ( 
.A(n_384),
.Y(n_411)
);

FAx1_ASAP7_75t_SL g384 ( 
.A(n_385),
.B(n_387),
.CI(n_388),
.CON(n_384),
.SN(n_384)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_385),
.B(n_387),
.C(n_388),
.Y(n_400)
);

INVx5_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_396),
.B(n_404),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_396),
.A2(n_409),
.B(n_410),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_402),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_397),
.B(n_402),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_400),
.C(n_401),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_398),
.B(n_407),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_400),
.B(n_401),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_406),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_405),
.B(n_406),
.Y(n_409)
);


endmodule