module fake_ariane_460_n_1942 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1942);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1942;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_604;
wire n_677;
wire n_439;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_65),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_61),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_36),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_38),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_124),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_77),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_3),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_195),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_51),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_56),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_35),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_147),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_46),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_44),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_187),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_140),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_17),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_104),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_74),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_113),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_100),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_12),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_184),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_39),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_137),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_50),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_0),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_153),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_120),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_4),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_61),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_54),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_32),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_145),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_150),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_106),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_115),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_86),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_11),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_23),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_46),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_85),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_110),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_107),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_158),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_109),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_102),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_149),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_103),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_108),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_79),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_14),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_112),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_63),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_155),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_73),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_173),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_36),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_15),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_186),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_141),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_99),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_45),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_114),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_81),
.Y(n_263)
);

BUFx5_ASAP7_75t_L g264 ( 
.A(n_91),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_30),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_144),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_131),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_57),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_176),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_64),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_133),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_143),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_121),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_16),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_26),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_159),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_10),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_160),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_126),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_47),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_10),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_22),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_90),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_95),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_6),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_181),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g287 ( 
.A(n_146),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_134),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_125),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_4),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_1),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_12),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_40),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_40),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_142),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_84),
.Y(n_296)
);

BUFx5_ASAP7_75t_L g297 ( 
.A(n_190),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_67),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_60),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_2),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_37),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_170),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_192),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_67),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_87),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_65),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_127),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_55),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_48),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_6),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_7),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_16),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_70),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_17),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_138),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_171),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_38),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_130),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_57),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_32),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_156),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_44),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_11),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_37),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_136),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_2),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_23),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_73),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_70),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_82),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_180),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_39),
.Y(n_332)
);

BUFx10_ASAP7_75t_L g333 ( 
.A(n_20),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_167),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_80),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_163),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_60),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_9),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_14),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_111),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_71),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_18),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_72),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_162),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_78),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_50),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_129),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_69),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_196),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_15),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_20),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_123),
.Y(n_352)
);

BUFx10_ASAP7_75t_L g353 ( 
.A(n_54),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_132),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_189),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_193),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_88),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_89),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_96),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_3),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_24),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_117),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_179),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_168),
.Y(n_364)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_164),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_94),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_41),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_71),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_98),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_22),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_27),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_52),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_45),
.Y(n_373)
);

INVx2_ASAP7_75t_SL g374 ( 
.A(n_93),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_175),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_119),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_28),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_83),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_53),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_152),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_178),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_8),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_166),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_118),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_42),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_58),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_13),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_41),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_174),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_75),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_197),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_311),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_197),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_197),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_310),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_273),
.Y(n_396)
);

CKINVDCx14_ASAP7_75t_R g397 ( 
.A(n_263),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_342),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_197),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_229),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_197),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_198),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_198),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_198),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_198),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_282),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_303),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_340),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_362),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_369),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_250),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_198),
.Y(n_412)
);

NOR2xp67_ASAP7_75t_L g413 ( 
.A(n_225),
.B(n_0),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_320),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_252),
.Y(n_415)
);

NOR2xp67_ASAP7_75t_L g416 ( 
.A(n_225),
.B(n_1),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_265),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_373),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_257),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_268),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_275),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_373),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_373),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_200),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_373),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_R g426 ( 
.A(n_262),
.B(n_151),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_317),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_209),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_373),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_350),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_333),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_277),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_298),
.Y(n_433)
);

INVxp33_ASAP7_75t_SL g434 ( 
.A(n_200),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_333),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_298),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_203),
.B(n_5),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_351),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_312),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_367),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_359),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_312),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_382),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_264),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_281),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_382),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_290),
.Y(n_447)
);

INVxp33_ASAP7_75t_SL g448 ( 
.A(n_204),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_204),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_206),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_292),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_333),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_202),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_202),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_299),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_389),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_242),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_300),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_301),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_264),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_264),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_242),
.Y(n_462)
);

OR2x2_ASAP7_75t_L g463 ( 
.A(n_209),
.B(n_7),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_255),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_263),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_206),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_263),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_306),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_308),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_353),
.B(n_9),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_255),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_313),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_370),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_322),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_384),
.Y(n_475)
);

BUFx6f_ASAP7_75t_SL g476 ( 
.A(n_287),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_287),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_384),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_199),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_212),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_370),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_372),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_220),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_287),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_372),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_326),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_233),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_264),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_222),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_428),
.B(n_318),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_444),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_453),
.B(n_207),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_444),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_444),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_453),
.B(n_217),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_481),
.B(n_251),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_454),
.B(n_221),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_418),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_391),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_460),
.A2(n_235),
.B(n_223),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_424),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_391),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_418),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_460),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_454),
.B(n_236),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_418),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_473),
.B(n_233),
.Y(n_507)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_407),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_482),
.B(n_251),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_460),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_393),
.Y(n_511)
);

BUFx8_ASAP7_75t_L g512 ( 
.A(n_476),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_461),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_400),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_393),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_449),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_419),
.Y(n_517)
);

OR2x2_ASAP7_75t_L g518 ( 
.A(n_473),
.B(n_319),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_394),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_461),
.Y(n_520)
);

NAND2xp33_ASAP7_75t_L g521 ( 
.A(n_426),
.B(n_264),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_457),
.B(n_241),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_461),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_394),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_457),
.B(n_244),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_485),
.B(n_237),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_488),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_462),
.B(n_246),
.Y(n_528)
);

NOR2x1_ASAP7_75t_L g529 ( 
.A(n_462),
.B(n_218),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_488),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_399),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_399),
.Y(n_532)
);

OR2x6_ASAP7_75t_L g533 ( 
.A(n_470),
.B(n_289),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_401),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_464),
.B(n_471),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_488),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_401),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_395),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_402),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_402),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_403),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_403),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_479),
.B(n_254),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_404),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_404),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_405),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_405),
.Y(n_547)
);

OA21x2_ASAP7_75t_L g548 ( 
.A1(n_412),
.A2(n_248),
.B(n_247),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_464),
.B(n_253),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_412),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_422),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_422),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_423),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_423),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_409),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_425),
.Y(n_556)
);

BUFx8_ASAP7_75t_L g557 ( 
.A(n_476),
.Y(n_557)
);

BUFx8_ASAP7_75t_L g558 ( 
.A(n_476),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_479),
.B(n_261),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_425),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_429),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_429),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_471),
.Y(n_563)
);

OA21x2_ASAP7_75t_L g564 ( 
.A1(n_475),
.A2(n_478),
.B(n_437),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_450),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_475),
.B(n_258),
.Y(n_566)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_487),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_478),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_433),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_496),
.B(n_397),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_496),
.B(n_467),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_496),
.B(n_411),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_568),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_535),
.B(n_467),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_568),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_535),
.Y(n_576)
);

BUFx8_ASAP7_75t_SL g577 ( 
.A(n_517),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_513),
.Y(n_578)
);

OR2x6_ASAP7_75t_L g579 ( 
.A(n_533),
.B(n_463),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_533),
.A2(n_476),
.B1(n_416),
.B2(n_413),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_535),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_518),
.Y(n_582)
);

OR2x6_ASAP7_75t_L g583 ( 
.A(n_533),
.B(n_463),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_518),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_504),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_504),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_518),
.B(n_406),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_496),
.B(n_415),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_510),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_513),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_513),
.Y(n_591)
);

BUFx4f_ASAP7_75t_L g592 ( 
.A(n_564),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_496),
.B(n_417),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_490),
.B(n_420),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_520),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_504),
.Y(n_596)
);

NAND3xp33_ASAP7_75t_L g597 ( 
.A(n_509),
.B(n_432),
.C(n_421),
.Y(n_597)
);

NAND3xp33_ASAP7_75t_L g598 ( 
.A(n_501),
.B(n_447),
.C(n_445),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_520),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_529),
.B(n_451),
.Y(n_600)
);

NAND2xp33_ASAP7_75t_R g601 ( 
.A(n_538),
.B(n_398),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_529),
.B(n_455),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_491),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_491),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_533),
.B(n_507),
.Y(n_605)
);

INVx6_ASAP7_75t_L g606 ( 
.A(n_512),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_504),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_555),
.Y(n_608)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_504),
.Y(n_609)
);

OR2x6_ASAP7_75t_L g610 ( 
.A(n_533),
.B(n_413),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_491),
.Y(n_611)
);

BUFx8_ASAP7_75t_SL g612 ( 
.A(n_517),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_533),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_535),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_491),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_535),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_501),
.B(n_458),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_508),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_516),
.B(n_459),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_504),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_SL g621 ( 
.A(n_512),
.B(n_465),
.Y(n_621)
);

NAND2xp33_ASAP7_75t_L g622 ( 
.A(n_504),
.B(n_264),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_493),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_569),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_507),
.B(n_468),
.Y(n_625)
);

NOR3xp33_ASAP7_75t_L g626 ( 
.A(n_516),
.B(n_256),
.C(n_469),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_493),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_520),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_521),
.A2(n_416),
.B1(n_414),
.B2(n_392),
.Y(n_629)
);

OAI22xp33_ASAP7_75t_SL g630 ( 
.A1(n_565),
.A2(n_434),
.B1(n_448),
.B2(n_435),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_565),
.B(n_472),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_520),
.Y(n_632)
);

OAI22xp33_ASAP7_75t_L g633 ( 
.A1(n_514),
.A2(n_452),
.B1(n_431),
.B2(n_474),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_493),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_493),
.Y(n_635)
);

OR2x6_ASAP7_75t_L g636 ( 
.A(n_526),
.B(n_489),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_507),
.B(n_486),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_520),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_510),
.Y(n_639)
);

NAND3xp33_ASAP7_75t_L g640 ( 
.A(n_521),
.B(n_466),
.C(n_211),
.Y(n_640)
);

INVx4_ASAP7_75t_L g641 ( 
.A(n_504),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_512),
.B(n_201),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_494),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_512),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_494),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_569),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_499),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_512),
.B(n_201),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_526),
.B(n_441),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_510),
.B(n_480),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_543),
.B(n_559),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_494),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_499),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_514),
.B(n_489),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_502),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_502),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_494),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_527),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_523),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_510),
.B(n_480),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_526),
.B(n_456),
.Y(n_661)
);

INVx4_ASAP7_75t_L g662 ( 
.A(n_527),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_557),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_563),
.Y(n_664)
);

OAI22xp33_ASAP7_75t_L g665 ( 
.A1(n_538),
.A2(n_208),
.B1(n_215),
.B2(n_211),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_527),
.Y(n_666)
);

AND2x6_ASAP7_75t_L g667 ( 
.A(n_557),
.B(n_321),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_511),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_538),
.B(n_477),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_536),
.B(n_483),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_543),
.B(n_483),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_557),
.B(n_205),
.Y(n_672)
);

OR2x2_ASAP7_75t_L g673 ( 
.A(n_508),
.B(n_208),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_557),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_536),
.B(n_564),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_564),
.A2(n_280),
.B1(n_379),
.B2(n_361),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_557),
.B(n_205),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g678 ( 
.A(n_567),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_523),
.Y(n_679)
);

OAI22xp5_ASAP7_75t_SL g680 ( 
.A1(n_567),
.A2(n_440),
.B1(n_438),
.B2(n_427),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_523),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_543),
.B(n_215),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_536),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_536),
.Y(n_684)
);

AND3x2_ASAP7_75t_L g685 ( 
.A(n_559),
.B(n_274),
.C(n_270),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_523),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_536),
.B(n_344),
.Y(n_687)
);

NAND2xp33_ASAP7_75t_L g688 ( 
.A(n_527),
.B(n_264),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_530),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_530),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_492),
.B(n_484),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_530),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_558),
.B(n_210),
.Y(n_693)
);

BUFx2_ASAP7_75t_L g694 ( 
.A(n_558),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_564),
.B(n_210),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_564),
.B(n_213),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_559),
.B(n_224),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_563),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_511),
.Y(n_699)
);

INVx5_ASAP7_75t_L g700 ( 
.A(n_527),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_530),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_558),
.B(n_213),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_540),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_548),
.A2(n_338),
.B1(n_332),
.B2(n_341),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_558),
.B(n_214),
.Y(n_705)
);

BUFx10_ASAP7_75t_L g706 ( 
.A(n_563),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_515),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_558),
.Y(n_708)
);

INVx1_ASAP7_75t_SL g709 ( 
.A(n_495),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_495),
.B(n_214),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_497),
.B(n_396),
.Y(n_711)
);

NAND3xp33_ASAP7_75t_L g712 ( 
.A(n_497),
.B(n_228),
.C(n_224),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_548),
.A2(n_304),
.B1(n_309),
.B2(n_328),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_515),
.Y(n_714)
);

NOR2x1p5_ASAP7_75t_L g715 ( 
.A(n_505),
.B(n_228),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_563),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_527),
.B(n_216),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_527),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_505),
.B(n_408),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_636),
.B(n_410),
.Y(n_720)
);

INVxp67_ASAP7_75t_L g721 ( 
.A(n_678),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_613),
.B(n_216),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_576),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_709),
.B(n_522),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_613),
.B(n_527),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_691),
.B(n_522),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_581),
.Y(n_727)
);

BUFx10_ASAP7_75t_L g728 ( 
.A(n_669),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_614),
.Y(n_729)
);

AND2x4_ASAP7_75t_SL g730 ( 
.A(n_608),
.B(n_430),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_637),
.A2(n_289),
.B1(n_365),
.B2(n_374),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_631),
.B(n_219),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_651),
.B(n_525),
.Y(n_733)
);

NAND2x1p5_ASAP7_75t_L g734 ( 
.A(n_674),
.B(n_563),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_616),
.Y(n_735)
);

INVx8_ASAP7_75t_L g736 ( 
.A(n_667),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_589),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_595),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_571),
.B(n_525),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_577),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_651),
.B(n_528),
.Y(n_741)
);

BUFx8_ASAP7_75t_L g742 ( 
.A(n_582),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_589),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_595),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_639),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_592),
.A2(n_676),
.B1(n_610),
.B2(n_636),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_671),
.B(n_528),
.Y(n_747)
);

BUFx6f_ASAP7_75t_SL g748 ( 
.A(n_582),
.Y(n_748)
);

A2O1A1Ixp33_ASAP7_75t_L g749 ( 
.A1(n_592),
.A2(n_500),
.B(n_566),
.C(n_549),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_671),
.B(n_549),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_625),
.B(n_566),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_605),
.B(n_563),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_592),
.B(n_563),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_588),
.B(n_329),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_579),
.A2(n_365),
.B1(n_374),
.B2(n_380),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_570),
.B(n_563),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_574),
.B(n_219),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_594),
.B(n_337),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_636),
.B(n_540),
.Y(n_759)
);

NAND2xp33_ASAP7_75t_SL g760 ( 
.A(n_708),
.B(n_230),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_585),
.B(n_500),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_636),
.B(n_540),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_599),
.Y(n_763)
);

AND2x2_ASAP7_75t_SL g764 ( 
.A(n_694),
.B(n_548),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_711),
.B(n_540),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_599),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_572),
.B(n_339),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_610),
.A2(n_548),
.B1(n_546),
.B2(n_560),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_574),
.B(n_226),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_600),
.B(n_226),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_593),
.B(n_719),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_602),
.B(n_343),
.Y(n_772)
);

NAND2xp33_ASAP7_75t_L g773 ( 
.A(n_667),
.B(n_227),
.Y(n_773)
);

NOR2xp67_ASAP7_75t_SL g774 ( 
.A(n_606),
.B(n_674),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_628),
.Y(n_775)
);

OR2x6_ASAP7_75t_L g776 ( 
.A(n_579),
.B(n_433),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_573),
.B(n_540),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_584),
.Y(n_778)
);

OAI22xp33_ASAP7_75t_L g779 ( 
.A1(n_579),
.A2(n_583),
.B1(n_610),
.B2(n_584),
.Y(n_779)
);

NAND2xp33_ASAP7_75t_SL g780 ( 
.A(n_708),
.B(n_230),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_585),
.B(n_500),
.Y(n_781)
);

AO221x1_ASAP7_75t_L g782 ( 
.A1(n_665),
.A2(n_633),
.B1(n_694),
.B2(n_680),
.C(n_618),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_606),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_579),
.B(n_285),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_585),
.B(n_227),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_578),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_578),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_575),
.B(n_624),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_597),
.B(n_346),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_618),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_632),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_646),
.B(n_541),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_673),
.B(n_232),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_580),
.B(n_541),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_649),
.B(n_661),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_703),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_650),
.B(n_541),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_660),
.B(n_541),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_632),
.Y(n_799)
);

NAND2x1p5_ASAP7_75t_L g800 ( 
.A(n_644),
.B(n_548),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_585),
.B(n_607),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_638),
.Y(n_802)
);

OR2x2_ASAP7_75t_SL g803 ( 
.A(n_673),
.B(n_291),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_590),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_638),
.B(n_541),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_583),
.A2(n_380),
.B1(n_234),
.B2(n_232),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_654),
.Y(n_807)
);

OR2x6_ASAP7_75t_L g808 ( 
.A(n_583),
.B(n_436),
.Y(n_808)
);

NOR2xp67_ASAP7_75t_L g809 ( 
.A(n_598),
.B(n_519),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_683),
.B(n_519),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_640),
.B(n_234),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_606),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_654),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_683),
.B(n_524),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_590),
.Y(n_815)
);

NOR2x1p5_ASAP7_75t_L g816 ( 
.A(n_587),
.B(n_231),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_587),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_610),
.A2(n_562),
.B1(n_524),
.B2(n_560),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_684),
.B(n_531),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_684),
.B(n_531),
.Y(n_820)
);

INVxp67_ASAP7_75t_SL g821 ( 
.A(n_585),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_647),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_607),
.B(n_620),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_607),
.B(n_349),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_710),
.B(n_348),
.Y(n_825)
);

NAND3xp33_ASAP7_75t_L g826 ( 
.A(n_629),
.B(n_238),
.C(n_231),
.Y(n_826)
);

NAND2x1p5_ASAP7_75t_L g827 ( 
.A(n_644),
.B(n_532),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_583),
.B(n_532),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_617),
.B(n_238),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_702),
.B(n_349),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_687),
.B(n_534),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_603),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_619),
.B(n_354),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_653),
.Y(n_834)
);

NOR3xp33_ASAP7_75t_L g835 ( 
.A(n_630),
.B(n_314),
.C(n_294),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_655),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_626),
.B(n_354),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_670),
.B(n_534),
.Y(n_838)
);

BUFx8_ASAP7_75t_L g839 ( 
.A(n_577),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_663),
.B(n_355),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_682),
.B(n_239),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_656),
.B(n_537),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_715),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_668),
.B(n_537),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_699),
.B(n_539),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_704),
.A2(n_562),
.B1(n_544),
.B2(n_556),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_707),
.Y(n_847)
);

NOR3xp33_ASAP7_75t_L g848 ( 
.A(n_712),
.B(n_324),
.C(n_323),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_714),
.B(n_539),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_690),
.B(n_544),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_604),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_682),
.B(n_239),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_697),
.B(n_353),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_690),
.B(n_545),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_607),
.B(n_355),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_697),
.B(n_293),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_692),
.B(n_545),
.Y(n_857)
);

NAND2x1p5_ASAP7_75t_L g858 ( 
.A(n_663),
.B(n_546),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_703),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_692),
.B(n_551),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_591),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_607),
.B(n_357),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_591),
.B(n_604),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_642),
.A2(n_383),
.B1(n_366),
.B2(n_358),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_611),
.B(n_551),
.Y(n_865)
);

AND2x2_ASAP7_75t_SL g866 ( 
.A(n_621),
.B(n_266),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_716),
.B(n_357),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_615),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_615),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_648),
.B(n_293),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_623),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_623),
.B(n_553),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_627),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_627),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_634),
.B(n_553),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_672),
.B(n_360),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_677),
.B(n_360),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_601),
.B(n_368),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_685),
.B(n_327),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_693),
.B(n_368),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_705),
.B(n_371),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_634),
.B(n_554),
.Y(n_882)
);

OAI22xp33_ASAP7_75t_L g883 ( 
.A1(n_695),
.A2(n_377),
.B1(n_371),
.B2(n_385),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_635),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_635),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_643),
.B(n_554),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_796),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_796),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_723),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_749),
.A2(n_675),
.B(n_696),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_801),
.A2(n_596),
.B(n_586),
.Y(n_891)
);

INVxp67_ASAP7_75t_L g892 ( 
.A(n_778),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_761),
.A2(n_645),
.B(n_643),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_795),
.B(n_436),
.Y(n_894)
);

O2A1O1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_726),
.A2(n_717),
.B(n_664),
.C(n_698),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_761),
.A2(n_652),
.B(n_645),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_801),
.A2(n_596),
.B(n_586),
.Y(n_897)
);

OAI21xp33_ASAP7_75t_L g898 ( 
.A1(n_841),
.A2(n_385),
.B(n_377),
.Y(n_898)
);

OAI22xp5_ASAP7_75t_L g899 ( 
.A1(n_751),
.A2(n_606),
.B1(n_716),
.B2(n_658),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_779),
.B(n_620),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_751),
.B(n_713),
.Y(n_901)
);

AO21x1_ASAP7_75t_L g902 ( 
.A1(n_753),
.A2(n_688),
.B(n_622),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_721),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_730),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_823),
.A2(n_596),
.B(n_586),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_823),
.A2(n_641),
.B(n_609),
.Y(n_906)
);

NAND2xp33_ASAP7_75t_L g907 ( 
.A(n_733),
.B(n_667),
.Y(n_907)
);

OAI22xp5_ASAP7_75t_L g908 ( 
.A1(n_746),
.A2(n_662),
.B1(n_609),
.B2(n_641),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_771),
.A2(n_664),
.B1(n_698),
.B2(n_658),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_739),
.B(n_724),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_753),
.A2(n_641),
.B(n_609),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_797),
.A2(n_662),
.B(n_658),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_779),
.B(n_620),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_817),
.B(n_439),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_739),
.B(n_652),
.Y(n_915)
);

OAI21xp33_ASAP7_75t_L g916 ( 
.A1(n_841),
.A2(n_387),
.B(n_386),
.Y(n_916)
);

AO21x1_ASAP7_75t_L g917 ( 
.A1(n_771),
.A2(n_688),
.B(n_622),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_839),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_746),
.B(n_620),
.Y(n_919)
);

NAND3xp33_ASAP7_75t_L g920 ( 
.A(n_790),
.B(n_387),
.C(n_386),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_798),
.A2(n_662),
.B(n_718),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_741),
.B(n_657),
.Y(n_922)
);

INVx4_ASAP7_75t_L g923 ( 
.A(n_776),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_852),
.A2(n_664),
.B(n_698),
.C(n_701),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_778),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_783),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_821),
.A2(n_666),
.B(n_620),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_790),
.B(n_657),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_781),
.A2(n_681),
.B(n_679),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_747),
.B(n_750),
.Y(n_930)
);

O2A1O1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_852),
.A2(n_689),
.B(n_686),
.C(n_681),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_781),
.A2(n_666),
.B(n_700),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_772),
.B(n_659),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_776),
.A2(n_666),
.B1(n_689),
.B2(n_679),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_805),
.A2(n_666),
.B(n_700),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_807),
.B(n_813),
.Y(n_936)
);

NOR3xp33_ASAP7_75t_L g937 ( 
.A(n_856),
.B(n_789),
.C(n_758),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_776),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_772),
.B(n_659),
.Y(n_939)
);

A2O1A1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_754),
.A2(n_278),
.B(n_335),
.C(n_284),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_783),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_754),
.B(n_667),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_752),
.A2(n_700),
.B(n_556),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_765),
.A2(n_666),
.B(n_700),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_853),
.B(n_706),
.Y(n_945)
);

O2A1O1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_856),
.A2(n_286),
.B(n_288),
.C(n_315),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_727),
.B(n_667),
.Y(n_947)
);

NOR2xp67_ASAP7_75t_L g948 ( 
.A(n_878),
.B(n_439),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_729),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_735),
.B(n_667),
.Y(n_950)
);

AOI22xp33_ASAP7_75t_L g951 ( 
.A1(n_782),
.A2(n_353),
.B1(n_547),
.B2(n_542),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_783),
.Y(n_952)
);

AOI21xp33_ASAP7_75t_L g953 ( 
.A1(n_758),
.A2(n_388),
.B(n_356),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_822),
.B(n_700),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_834),
.Y(n_955)
);

A2O1A1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_789),
.A2(n_330),
.B(n_352),
.C(n_364),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_836),
.B(n_706),
.Y(n_957)
);

NOR2x1_ASAP7_75t_L g958 ( 
.A(n_720),
.B(n_336),
.Y(n_958)
);

O2A1O1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_883),
.A2(n_561),
.B(n_550),
.C(n_547),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_847),
.B(n_706),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_738),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_788),
.B(n_388),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_870),
.A2(n_358),
.B1(n_363),
.B2(n_366),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_793),
.B(n_363),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_744),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_763),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_863),
.A2(n_375),
.B(n_376),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_742),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_832),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_808),
.A2(n_383),
.B1(n_376),
.B2(n_378),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_883),
.B(n_375),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_784),
.B(n_378),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_720),
.B(n_442),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_777),
.A2(n_381),
.B(n_267),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_756),
.A2(n_561),
.B(n_550),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_870),
.B(n_442),
.Y(n_976)
);

OAI21xp5_ASAP7_75t_L g977 ( 
.A1(n_859),
.A2(n_561),
.B(n_550),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_792),
.A2(n_269),
.B(n_240),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_783),
.Y(n_979)
);

AOI22xp33_ASAP7_75t_L g980 ( 
.A1(n_866),
.A2(n_547),
.B1(n_542),
.B2(n_443),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_812),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_757),
.B(n_13),
.Y(n_982)
);

INVx3_ASAP7_75t_L g983 ( 
.A(n_812),
.Y(n_983)
);

AOI22xp5_ASAP7_75t_L g984 ( 
.A1(n_876),
.A2(n_307),
.B1(n_245),
.B2(n_249),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_838),
.A2(n_271),
.B(n_260),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_766),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_736),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_775),
.A2(n_542),
.B(n_503),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_851),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_850),
.A2(n_857),
.B(n_854),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_860),
.A2(n_259),
.B(n_243),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_769),
.B(n_18),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_742),
.B(n_806),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_818),
.B(n_552),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_876),
.B(n_443),
.Y(n_995)
);

INVx2_ASAP7_75t_SL g996 ( 
.A(n_728),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_810),
.A2(n_272),
.B(n_276),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_877),
.B(n_880),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_791),
.A2(n_498),
.B(n_503),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_814),
.A2(n_325),
.B(n_283),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_803),
.B(n_19),
.Y(n_1001)
);

NAND2xp33_ASAP7_75t_L g1002 ( 
.A(n_736),
.B(n_552),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_819),
.A2(n_331),
.B(n_295),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_820),
.A2(n_279),
.B(n_296),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_831),
.A2(n_345),
.B(n_305),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_877),
.B(n_880),
.Y(n_1006)
);

INVx1_ASAP7_75t_SL g1007 ( 
.A(n_740),
.Y(n_1007)
);

AOI21xp33_ASAP7_75t_L g1008 ( 
.A1(n_829),
.A2(n_446),
.B(n_506),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_725),
.A2(n_347),
.B(n_316),
.Y(n_1009)
);

AND2x4_ASAP7_75t_SL g1010 ( 
.A(n_808),
.B(n_612),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_881),
.A2(n_506),
.B(n_498),
.C(n_446),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_725),
.A2(n_390),
.B(n_302),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_881),
.B(n_506),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_829),
.A2(n_552),
.B(n_334),
.C(n_321),
.Y(n_1014)
);

NAND2xp33_ASAP7_75t_L g1015 ( 
.A(n_736),
.B(n_552),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_818),
.A2(n_755),
.B1(n_762),
.B2(n_759),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_861),
.A2(n_799),
.B(n_802),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_865),
.A2(n_334),
.B(n_321),
.Y(n_1018)
);

INVx1_ASAP7_75t_SL g1019 ( 
.A(n_760),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_872),
.A2(n_334),
.B(n_321),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_826),
.B(n_19),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_843),
.B(n_612),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_875),
.A2(n_334),
.B(n_321),
.Y(n_1023)
);

NOR2x1_ASAP7_75t_L g1024 ( 
.A(n_816),
.B(n_552),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_882),
.A2(n_334),
.B(n_552),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_868),
.A2(n_552),
.B(n_297),
.Y(n_1026)
);

AO21x1_ASAP7_75t_L g1027 ( 
.A1(n_785),
.A2(n_862),
.B(n_824),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_827),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_886),
.A2(n_552),
.B(n_297),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_842),
.Y(n_1030)
);

NOR2x1p5_ASAP7_75t_L g1031 ( 
.A(n_839),
.B(n_21),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_844),
.A2(n_297),
.B(n_264),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_845),
.A2(n_297),
.B(n_194),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_871),
.Y(n_1034)
);

OAI321xp33_ASAP7_75t_L g1035 ( 
.A1(n_731),
.A2(n_21),
.A3(n_24),
.B1(n_25),
.B2(n_26),
.C(n_27),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_748),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_767),
.B(n_732),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_866),
.B(n_25),
.Y(n_1038)
);

NAND2x1p5_ASAP7_75t_L g1039 ( 
.A(n_774),
.B(n_148),
.Y(n_1039)
);

AOI21xp33_ASAP7_75t_L g1040 ( 
.A1(n_825),
.A2(n_28),
.B(n_29),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_748),
.Y(n_1041)
);

CKINVDCx8_ASAP7_75t_R g1042 ( 
.A(n_879),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_767),
.B(n_29),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_849),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_885),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_828),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_825),
.B(n_31),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_728),
.B(n_297),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_879),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_867),
.A2(n_297),
.B(n_76),
.Y(n_1050)
);

OAI21xp33_ASAP7_75t_L g1051 ( 
.A1(n_864),
.A2(n_33),
.B(n_34),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_737),
.B(n_34),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_L g1053 ( 
.A(n_743),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_827),
.B(n_297),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_745),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_869),
.A2(n_297),
.B(n_97),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_809),
.B(n_42),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_858),
.B(n_43),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_770),
.A2(n_830),
.B(n_785),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_824),
.A2(n_92),
.B(n_188),
.Y(n_1060)
);

INVxp67_ASAP7_75t_L g1061 ( 
.A(n_794),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_858),
.B(n_43),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_873),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_1063)
);

BUFx12f_ASAP7_75t_L g1064 ( 
.A(n_734),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_884),
.B(n_49),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_855),
.A2(n_862),
.B(n_722),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_855),
.A2(n_105),
.B(n_185),
.Y(n_1067)
);

OAI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_874),
.A2(n_768),
.B(n_787),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_848),
.B(n_51),
.Y(n_1069)
);

AOI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_780),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_768),
.A2(n_58),
.B1(n_59),
.B2(n_62),
.Y(n_1071)
);

NOR2xp67_ASAP7_75t_L g1072 ( 
.A(n_840),
.B(n_128),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_773),
.A2(n_122),
.B(n_183),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_937),
.B(n_835),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_937),
.A2(n_811),
.B(n_837),
.C(n_833),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_910),
.A2(n_764),
.B1(n_734),
.B2(n_846),
.Y(n_1076)
);

BUFx2_ASAP7_75t_L g1077 ( 
.A(n_903),
.Y(n_1077)
);

AOI22x1_ASAP7_75t_L g1078 ( 
.A1(n_990),
.A2(n_800),
.B1(n_815),
.B2(n_804),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_998),
.A2(n_786),
.B(n_846),
.C(n_800),
.Y(n_1079)
);

CKINVDCx11_ASAP7_75t_R g1080 ( 
.A(n_918),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_915),
.A2(n_764),
.B(n_62),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_930),
.A2(n_59),
.B1(n_63),
.B2(n_64),
.Y(n_1082)
);

AO32x2_ASAP7_75t_L g1083 ( 
.A1(n_1071),
.A2(n_66),
.A3(n_68),
.B1(n_69),
.B2(n_72),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_1006),
.B(n_66),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_894),
.B(n_68),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1030),
.B(n_101),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_955),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_1037),
.B(n_116),
.Y(n_1088)
);

INVx1_ASAP7_75t_SL g1089 ( 
.A(n_973),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_933),
.A2(n_135),
.B(n_139),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_936),
.B(n_191),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1044),
.B(n_154),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_1037),
.B(n_157),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_901),
.A2(n_161),
.B1(n_165),
.B2(n_172),
.Y(n_1094)
);

O2A1O1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_1040),
.A2(n_177),
.B(n_1047),
.C(n_1043),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_892),
.B(n_925),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_892),
.B(n_925),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_R g1098 ( 
.A(n_1041),
.B(n_1042),
.Y(n_1098)
);

OR2x2_ASAP7_75t_L g1099 ( 
.A(n_936),
.B(n_904),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_1049),
.Y(n_1100)
);

AOI21x1_ASAP7_75t_L g1101 ( 
.A1(n_900),
.A2(n_913),
.B(n_1027),
.Y(n_1101)
);

O2A1O1Ixp5_ASAP7_75t_SL g1102 ( 
.A1(n_953),
.A2(n_1008),
.B(n_1058),
.C(n_1048),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_889),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_945),
.A2(n_960),
.B1(n_957),
.B2(n_928),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_914),
.B(n_1001),
.Y(n_1105)
);

A2O1A1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_946),
.A2(n_1021),
.B(n_982),
.C(n_992),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_926),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_1019),
.B(n_923),
.Y(n_1108)
);

CKINVDCx20_ASAP7_75t_R g1109 ( 
.A(n_1007),
.Y(n_1109)
);

O2A1O1Ixp33_ASAP7_75t_SL g1110 ( 
.A1(n_1058),
.A2(n_942),
.B(n_954),
.C(n_1062),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_939),
.A2(n_890),
.B(n_943),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_948),
.B(n_928),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_923),
.B(n_996),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_898),
.B(n_916),
.Y(n_1114)
);

AOI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_945),
.A2(n_1001),
.B1(n_1038),
.B2(n_964),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_SL g1116 ( 
.A(n_968),
.B(n_1010),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_969),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_938),
.B(n_958),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_899),
.A2(n_895),
.B(n_912),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_949),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_962),
.B(n_976),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_938),
.B(n_964),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_932),
.A2(n_911),
.B(n_921),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_989),
.Y(n_1124)
);

AO21x1_ASAP7_75t_L g1125 ( 
.A1(n_1056),
.A2(n_900),
.B(n_913),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_926),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_993),
.B(n_972),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_995),
.B(n_961),
.Y(n_1128)
);

CKINVDCx20_ASAP7_75t_R g1129 ( 
.A(n_1036),
.Y(n_1129)
);

INVx2_ASAP7_75t_SL g1130 ( 
.A(n_1036),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_963),
.A2(n_992),
.B1(n_982),
.B2(n_1021),
.Y(n_1131)
);

OAI21xp33_ASAP7_75t_SL g1132 ( 
.A1(n_965),
.A2(n_986),
.B(n_966),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_970),
.B(n_1016),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_926),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_987),
.Y(n_1135)
);

O2A1O1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_940),
.A2(n_1035),
.B(n_1046),
.C(n_1051),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_1028),
.B(n_987),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1053),
.B(n_922),
.Y(n_1138)
);

A2O1A1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_956),
.A2(n_931),
.B(n_1069),
.C(n_924),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_1053),
.B(n_920),
.Y(n_1140)
);

NAND2x1p5_ASAP7_75t_L g1141 ( 
.A(n_1028),
.B(n_987),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_1022),
.B(n_971),
.Y(n_1142)
);

O2A1O1Ixp33_ASAP7_75t_SL g1143 ( 
.A1(n_1054),
.A2(n_1063),
.B(n_1017),
.C(n_909),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_944),
.A2(n_907),
.B(n_905),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_891),
.A2(n_906),
.B(n_897),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_951),
.B(n_1024),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1059),
.A2(n_1066),
.B(n_1057),
.C(n_1061),
.Y(n_1147)
);

INVxp67_ASAP7_75t_SL g1148 ( 
.A(n_1002),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_984),
.A2(n_951),
.B1(n_1070),
.B2(n_934),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1061),
.B(n_980),
.Y(n_1150)
);

OR2x6_ASAP7_75t_L g1151 ( 
.A(n_1064),
.B(n_987),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_908),
.A2(n_887),
.B1(n_888),
.B2(n_1045),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_980),
.B(n_983),
.Y(n_1153)
);

INVx4_ASAP7_75t_L g1154 ( 
.A(n_981),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_926),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1031),
.B(n_1034),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_981),
.A2(n_983),
.B1(n_919),
.B2(n_1005),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_L g1158 ( 
.A(n_952),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1055),
.B(n_952),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1065),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1052),
.Y(n_1161)
);

AO21x1_ASAP7_75t_L g1162 ( 
.A1(n_919),
.A2(n_1033),
.B(n_1054),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_941),
.Y(n_1163)
);

O2A1O1Ixp33_ASAP7_75t_SL g1164 ( 
.A1(n_947),
.A2(n_950),
.B(n_994),
.C(n_935),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_941),
.B(n_979),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_959),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_952),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_979),
.B(n_994),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1013),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1068),
.B(n_979),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_979),
.B(n_967),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_977),
.B(n_988),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_985),
.A2(n_974),
.B1(n_1000),
.B2(n_1004),
.Y(n_1173)
);

AOI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1029),
.A2(n_902),
.B(n_1025),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1015),
.A2(n_893),
.B(n_896),
.Y(n_1175)
);

INVx2_ASAP7_75t_SL g1176 ( 
.A(n_1039),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_1072),
.A2(n_917),
.B1(n_975),
.B2(n_1012),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_1009),
.B(n_1003),
.Y(n_1178)
);

O2A1O1Ixp5_ASAP7_75t_SL g1179 ( 
.A1(n_929),
.A2(n_1026),
.B(n_999),
.C(n_1032),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1011),
.B(n_997),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_991),
.B(n_1039),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1050),
.A2(n_1067),
.B(n_1060),
.C(n_1073),
.Y(n_1182)
);

INVx2_ASAP7_75t_SL g1183 ( 
.A(n_1014),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_978),
.A2(n_1018),
.B(n_1020),
.C(n_1023),
.Y(n_1184)
);

INVx2_ASAP7_75t_SL g1185 ( 
.A(n_927),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_910),
.B(n_618),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_937),
.B(n_790),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_955),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_990),
.A2(n_915),
.B(n_930),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_910),
.B(n_618),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_910),
.B(n_618),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_926),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_910),
.B(n_618),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_937),
.B(n_790),
.Y(n_1194)
);

O2A1O1Ixp5_ASAP7_75t_L g1195 ( 
.A1(n_1047),
.A2(n_1027),
.B(n_1043),
.C(n_1058),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_973),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_990),
.A2(n_915),
.B(n_930),
.Y(n_1197)
);

NAND2xp33_ASAP7_75t_L g1198 ( 
.A(n_937),
.B(n_930),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_918),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_910),
.B(n_930),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_937),
.B(n_790),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_910),
.B(n_618),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_SL g1203 ( 
.A1(n_1001),
.A2(n_618),
.B1(n_669),
.B2(n_517),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_937),
.B(n_790),
.Y(n_1204)
);

AO21x1_ASAP7_75t_L g1205 ( 
.A1(n_937),
.A2(n_1006),
.B(n_998),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_937),
.A2(n_795),
.B1(n_661),
.B2(n_649),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_990),
.A2(n_915),
.B(n_930),
.Y(n_1207)
);

OR2x2_ASAP7_75t_L g1208 ( 
.A(n_910),
.B(n_817),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_990),
.A2(n_915),
.B(n_930),
.Y(n_1209)
);

CKINVDCx6p67_ASAP7_75t_R g1210 ( 
.A(n_918),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_937),
.B(n_790),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_910),
.B(n_930),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_903),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_990),
.A2(n_915),
.B(n_930),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_937),
.A2(n_998),
.B(n_1006),
.C(n_1037),
.Y(n_1215)
);

AND3x2_ASAP7_75t_L g1216 ( 
.A(n_937),
.B(n_621),
.C(n_669),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_910),
.B(n_618),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_955),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_R g1219 ( 
.A(n_1041),
.B(n_618),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_937),
.B(n_790),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_955),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_910),
.B(n_930),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_910),
.B(n_930),
.Y(n_1223)
);

A2O1A1Ixp33_ASAP7_75t_SL g1224 ( 
.A1(n_937),
.A2(n_631),
.B(n_637),
.C(n_841),
.Y(n_1224)
);

O2A1O1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_937),
.A2(n_998),
.B(n_1006),
.C(n_726),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_910),
.B(n_618),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_937),
.B(n_790),
.Y(n_1227)
);

AO31x2_ASAP7_75t_L g1228 ( 
.A1(n_1125),
.A2(n_1162),
.A3(n_1147),
.B(n_1205),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1186),
.A2(n_1191),
.B(n_1190),
.Y(n_1229)
);

BUFx10_ASAP7_75t_L g1230 ( 
.A(n_1199),
.Y(n_1230)
);

BUFx12f_ASAP7_75t_L g1231 ( 
.A(n_1080),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1078),
.A2(n_1144),
.B(n_1145),
.Y(n_1232)
);

BUFx8_ASAP7_75t_L g1233 ( 
.A(n_1077),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1206),
.A2(n_1131),
.B1(n_1200),
.B2(n_1212),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1087),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1193),
.B(n_1202),
.Y(n_1236)
);

AO32x2_ASAP7_75t_L g1237 ( 
.A1(n_1152),
.A2(n_1082),
.A3(n_1076),
.B1(n_1157),
.B2(n_1185),
.Y(n_1237)
);

AOI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1203),
.A2(n_1226),
.B1(n_1217),
.B2(n_1115),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1103),
.Y(n_1239)
);

NAND3x1_ASAP7_75t_L g1240 ( 
.A(n_1142),
.B(n_1127),
.C(n_1122),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1111),
.A2(n_1209),
.A3(n_1189),
.B(n_1197),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1189),
.A2(n_1207),
.B(n_1197),
.Y(n_1242)
);

BUFx3_ASAP7_75t_L g1243 ( 
.A(n_1213),
.Y(n_1243)
);

OAI22x1_ASAP7_75t_L g1244 ( 
.A1(n_1149),
.A2(n_1074),
.B1(n_1118),
.B2(n_1227),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1207),
.A2(n_1209),
.B(n_1214),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1196),
.B(n_1105),
.Y(n_1246)
);

OAI22x1_ASAP7_75t_L g1247 ( 
.A1(n_1118),
.A2(n_1201),
.B1(n_1220),
.B2(n_1211),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1222),
.B(n_1223),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1120),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1188),
.Y(n_1250)
);

O2A1O1Ixp33_ASAP7_75t_SL g1251 ( 
.A1(n_1224),
.A2(n_1215),
.B(n_1133),
.C(n_1225),
.Y(n_1251)
);

AO31x2_ASAP7_75t_L g1252 ( 
.A1(n_1111),
.A2(n_1214),
.A3(n_1119),
.B(n_1144),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1196),
.B(n_1089),
.Y(n_1253)
);

AO21x2_ASAP7_75t_L g1254 ( 
.A1(n_1079),
.A2(n_1123),
.B(n_1119),
.Y(n_1254)
);

A2O1A1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1106),
.A2(n_1225),
.B(n_1093),
.C(n_1136),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1208),
.B(n_1187),
.Y(n_1256)
);

INVx2_ASAP7_75t_SL g1257 ( 
.A(n_1098),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1148),
.A2(n_1182),
.B(n_1110),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1198),
.B(n_1138),
.Y(n_1259)
);

A2O1A1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1136),
.A2(n_1114),
.B(n_1095),
.C(n_1075),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1148),
.A2(n_1175),
.B(n_1123),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1096),
.B(n_1097),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1175),
.A2(n_1145),
.B(n_1104),
.Y(n_1263)
);

INVx3_ASAP7_75t_L g1264 ( 
.A(n_1137),
.Y(n_1264)
);

INVx3_ASAP7_75t_SL g1265 ( 
.A(n_1210),
.Y(n_1265)
);

INVx8_ASAP7_75t_L g1266 ( 
.A(n_1109),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1100),
.B(n_1099),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_1151),
.Y(n_1268)
);

AOI221x1_ASAP7_75t_L g1269 ( 
.A1(n_1081),
.A2(n_1139),
.B1(n_1090),
.B2(n_1094),
.C(n_1112),
.Y(n_1269)
);

NAND2x1_ASAP7_75t_L g1270 ( 
.A(n_1154),
.B(n_1155),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1195),
.A2(n_1095),
.B(n_1121),
.Y(n_1271)
);

OAI21xp33_ASAP7_75t_L g1272 ( 
.A1(n_1084),
.A2(n_1085),
.B(n_1081),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_SL g1273 ( 
.A1(n_1091),
.A2(n_1146),
.B1(n_1150),
.B2(n_1140),
.Y(n_1273)
);

INVx1_ASAP7_75t_SL g1274 ( 
.A(n_1219),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1174),
.A2(n_1179),
.B(n_1184),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1128),
.B(n_1108),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1181),
.A2(n_1172),
.B(n_1143),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1184),
.A2(n_1079),
.B(n_1101),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1132),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1178),
.A2(n_1180),
.B(n_1173),
.Y(n_1280)
);

INVx3_ASAP7_75t_SL g1281 ( 
.A(n_1129),
.Y(n_1281)
);

NAND3x1_ASAP7_75t_L g1282 ( 
.A(n_1113),
.B(n_1156),
.C(n_1216),
.Y(n_1282)
);

AOI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1116),
.A2(n_1204),
.B1(n_1194),
.B2(n_1216),
.Y(n_1283)
);

A2O1A1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1075),
.A2(n_1195),
.B(n_1160),
.C(n_1161),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1130),
.Y(n_1285)
);

O2A1O1Ixp5_ASAP7_75t_SL g1286 ( 
.A1(n_1159),
.A2(n_1088),
.B(n_1166),
.C(n_1221),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1218),
.B(n_1169),
.Y(n_1287)
);

O2A1O1Ixp33_ASAP7_75t_SL g1288 ( 
.A1(n_1171),
.A2(n_1086),
.B(n_1092),
.C(n_1176),
.Y(n_1288)
);

O2A1O1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1164),
.A2(n_1153),
.B(n_1177),
.C(n_1163),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1168),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1117),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1124),
.A2(n_1168),
.B1(n_1183),
.B2(n_1151),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1177),
.A2(n_1165),
.B(n_1155),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1165),
.A2(n_1192),
.B(n_1167),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1107),
.A2(n_1192),
.B(n_1167),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1083),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1107),
.A2(n_1192),
.B(n_1167),
.Y(n_1297)
);

AND2x2_ASAP7_75t_SL g1298 ( 
.A(n_1083),
.B(n_1158),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1107),
.Y(n_1299)
);

AO32x2_ASAP7_75t_L g1300 ( 
.A1(n_1083),
.A2(n_1102),
.A3(n_1126),
.B1(n_1134),
.B2(n_1158),
.Y(n_1300)
);

OAI222xp33_ASAP7_75t_L g1301 ( 
.A1(n_1083),
.A2(n_1141),
.B1(n_1135),
.B2(n_1158),
.C1(n_1126),
.C2(n_1134),
.Y(n_1301)
);

NAND3x1_ASAP7_75t_L g1302 ( 
.A(n_1135),
.B(n_937),
.C(n_1131),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1134),
.Y(n_1303)
);

O2A1O1Ixp33_ASAP7_75t_SL g1304 ( 
.A1(n_1224),
.A2(n_1215),
.B(n_1133),
.C(n_1212),
.Y(n_1304)
);

A2O1A1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1131),
.A2(n_937),
.B(n_1006),
.C(n_998),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1078),
.A2(n_1144),
.B(n_1145),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1151),
.B(n_923),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1078),
.A2(n_1144),
.B(n_1145),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_SL g1309 ( 
.A(n_1116),
.B(n_618),
.Y(n_1309)
);

AO21x1_ASAP7_75t_L g1310 ( 
.A1(n_1133),
.A2(n_937),
.B(n_998),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1087),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1089),
.B(n_1196),
.Y(n_1312)
);

AOI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1131),
.A2(n_937),
.B1(n_795),
.B2(n_618),
.Y(n_1313)
);

NAND3xp33_ASAP7_75t_L g1314 ( 
.A(n_1106),
.B(n_937),
.C(n_1131),
.Y(n_1314)
);

A2O1A1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1131),
.A2(n_937),
.B(n_1006),
.C(n_998),
.Y(n_1315)
);

OA21x2_ASAP7_75t_L g1316 ( 
.A1(n_1123),
.A2(n_1119),
.B(n_1195),
.Y(n_1316)
);

O2A1O1Ixp33_ASAP7_75t_SL g1317 ( 
.A1(n_1224),
.A2(n_1215),
.B(n_1133),
.C(n_1212),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1189),
.A2(n_1207),
.B(n_1197),
.Y(n_1318)
);

AOI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1131),
.A2(n_937),
.B1(n_795),
.B2(n_618),
.Y(n_1319)
);

OAI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1131),
.A2(n_998),
.B1(n_1006),
.B2(n_1115),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1189),
.A2(n_1207),
.B(n_1197),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1206),
.A2(n_1131),
.B1(n_1212),
.B2(n_1200),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_1186),
.B(n_1190),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1219),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1078),
.A2(n_1144),
.B(n_1145),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1087),
.Y(n_1326)
);

AOI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1131),
.A2(n_937),
.B1(n_795),
.B2(n_618),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1078),
.A2(n_1144),
.B(n_1145),
.Y(n_1328)
);

A2O1A1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1131),
.A2(n_937),
.B(n_1006),
.C(n_998),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_1219),
.Y(n_1330)
);

INVx5_ASAP7_75t_L g1331 ( 
.A(n_1151),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1087),
.Y(n_1332)
);

INVx2_ASAP7_75t_SL g1333 ( 
.A(n_1098),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1078),
.A2(n_1144),
.B(n_1145),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1137),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1131),
.B(n_937),
.Y(n_1336)
);

AO31x2_ASAP7_75t_L g1337 ( 
.A1(n_1125),
.A2(n_1162),
.A3(n_1027),
.B(n_1147),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1189),
.A2(n_1207),
.B(n_1197),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1186),
.B(n_1217),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1186),
.B(n_1190),
.Y(n_1340)
);

NAND3xp33_ASAP7_75t_L g1341 ( 
.A(n_1106),
.B(n_937),
.C(n_1131),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1189),
.A2(n_1207),
.B(n_1197),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1186),
.B(n_1190),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1078),
.A2(n_1144),
.B(n_1145),
.Y(n_1344)
);

AO21x2_ASAP7_75t_L g1345 ( 
.A1(n_1111),
.A2(n_890),
.B(n_1056),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1189),
.A2(n_1207),
.B(n_1197),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1186),
.B(n_1217),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1186),
.B(n_1217),
.Y(n_1348)
);

AO31x2_ASAP7_75t_L g1349 ( 
.A1(n_1125),
.A2(n_1162),
.A3(n_1027),
.B(n_1147),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1186),
.A2(n_1191),
.B(n_1190),
.Y(n_1350)
);

OAI21xp33_ASAP7_75t_L g1351 ( 
.A1(n_1206),
.A2(n_937),
.B(n_1131),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1186),
.B(n_1217),
.Y(n_1352)
);

BUFx6f_ASAP7_75t_L g1353 ( 
.A(n_1151),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1151),
.B(n_923),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1189),
.A2(n_1207),
.B(n_1197),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_SL g1356 ( 
.A(n_1131),
.B(n_937),
.Y(n_1356)
);

AOI221xp5_ASAP7_75t_SL g1357 ( 
.A1(n_1215),
.A2(n_1225),
.B1(n_1198),
.B2(n_1106),
.C(n_946),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1186),
.B(n_1190),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1189),
.A2(n_1207),
.B(n_1197),
.Y(n_1359)
);

BUFx12f_ASAP7_75t_L g1360 ( 
.A(n_1080),
.Y(n_1360)
);

A2O1A1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1131),
.A2(n_937),
.B(n_1006),
.C(n_998),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1170),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1186),
.B(n_1217),
.Y(n_1363)
);

NAND3xp33_ASAP7_75t_L g1364 ( 
.A(n_1106),
.B(n_937),
.C(n_1131),
.Y(n_1364)
);

BUFx8_ASAP7_75t_L g1365 ( 
.A(n_1077),
.Y(n_1365)
);

O2A1O1Ixp33_ASAP7_75t_L g1366 ( 
.A1(n_1224),
.A2(n_937),
.B(n_1215),
.C(n_1006),
.Y(n_1366)
);

CKINVDCx20_ASAP7_75t_R g1367 ( 
.A(n_1219),
.Y(n_1367)
);

A2O1A1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1131),
.A2(n_937),
.B(n_1006),
.C(n_998),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1189),
.A2(n_1207),
.B(n_1197),
.Y(n_1369)
);

NOR2xp67_ASAP7_75t_L g1370 ( 
.A(n_1208),
.B(n_996),
.Y(n_1370)
);

OAI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1186),
.A2(n_1191),
.B(n_1190),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1206),
.A2(n_1131),
.B1(n_1212),
.B2(n_1200),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1087),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1078),
.A2(n_1144),
.B(n_1145),
.Y(n_1374)
);

AO21x1_ASAP7_75t_L g1375 ( 
.A1(n_1133),
.A2(n_937),
.B(n_998),
.Y(n_1375)
);

OR2x6_ASAP7_75t_L g1376 ( 
.A(n_1151),
.B(n_904),
.Y(n_1376)
);

AO31x2_ASAP7_75t_L g1377 ( 
.A1(n_1125),
.A2(n_1162),
.A3(n_1027),
.B(n_1147),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1087),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1170),
.Y(n_1379)
);

AO32x2_ASAP7_75t_L g1380 ( 
.A1(n_1152),
.A2(n_1071),
.A3(n_1082),
.B1(n_1076),
.B2(n_1157),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1186),
.B(n_1217),
.Y(n_1381)
);

NAND3xp33_ASAP7_75t_L g1382 ( 
.A(n_1106),
.B(n_937),
.C(n_1131),
.Y(n_1382)
);

NOR2xp67_ASAP7_75t_L g1383 ( 
.A(n_1208),
.B(n_996),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1238),
.A2(n_1327),
.B1(n_1319),
.B2(n_1313),
.Y(n_1384)
);

INVx6_ASAP7_75t_L g1385 ( 
.A(n_1331),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1351),
.A2(n_1336),
.B1(n_1356),
.B2(n_1382),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1248),
.B(n_1276),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1243),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1264),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1235),
.Y(n_1390)
);

BUFx10_ASAP7_75t_L g1391 ( 
.A(n_1330),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_SL g1392 ( 
.A1(n_1314),
.A2(n_1341),
.B1(n_1364),
.B2(n_1298),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_1367),
.Y(n_1393)
);

INVx4_ASAP7_75t_L g1394 ( 
.A(n_1266),
.Y(n_1394)
);

CKINVDCx14_ASAP7_75t_R g1395 ( 
.A(n_1324),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1320),
.A2(n_1234),
.B1(n_1372),
.B2(n_1322),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1239),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1335),
.Y(n_1398)
);

INVx8_ASAP7_75t_L g1399 ( 
.A(n_1266),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1246),
.B(n_1253),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1249),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1250),
.Y(n_1402)
);

INVx3_ASAP7_75t_L g1403 ( 
.A(n_1335),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1312),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1311),
.Y(n_1405)
);

BUFx2_ASAP7_75t_L g1406 ( 
.A(n_1233),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1273),
.A2(n_1358),
.B1(n_1343),
.B2(n_1323),
.Y(n_1407)
);

INVx5_ASAP7_75t_L g1408 ( 
.A(n_1376),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_SL g1409 ( 
.A1(n_1229),
.A2(n_1350),
.B1(n_1371),
.B2(n_1340),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1310),
.A2(n_1375),
.B1(n_1381),
.B2(n_1352),
.Y(n_1410)
);

INVx4_ASAP7_75t_SL g1411 ( 
.A(n_1268),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1326),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1332),
.Y(n_1413)
);

INVxp67_ASAP7_75t_SL g1414 ( 
.A(n_1287),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_SL g1415 ( 
.A1(n_1236),
.A2(n_1347),
.B1(n_1363),
.B2(n_1348),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1339),
.A2(n_1244),
.B1(n_1272),
.B2(n_1271),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_SL g1417 ( 
.A1(n_1309),
.A2(n_1296),
.B1(n_1353),
.B2(n_1268),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_1233),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_SL g1419 ( 
.A1(n_1296),
.A2(n_1268),
.B1(n_1353),
.B2(n_1279),
.Y(n_1419)
);

INVx4_ASAP7_75t_L g1420 ( 
.A(n_1265),
.Y(n_1420)
);

INVx1_ASAP7_75t_SL g1421 ( 
.A(n_1274),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1262),
.A2(n_1259),
.B1(n_1256),
.B2(n_1247),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1373),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1378),
.A2(n_1283),
.B1(n_1279),
.B2(n_1291),
.Y(n_1424)
);

BUFx8_ASAP7_75t_L g1425 ( 
.A(n_1231),
.Y(n_1425)
);

BUFx3_ASAP7_75t_L g1426 ( 
.A(n_1303),
.Y(n_1426)
);

INVx4_ASAP7_75t_L g1427 ( 
.A(n_1230),
.Y(n_1427)
);

BUFx12f_ASAP7_75t_L g1428 ( 
.A(n_1360),
.Y(n_1428)
);

INVx2_ASAP7_75t_SL g1429 ( 
.A(n_1230),
.Y(n_1429)
);

INVx6_ASAP7_75t_L g1430 ( 
.A(n_1365),
.Y(n_1430)
);

BUFx2_ASAP7_75t_SL g1431 ( 
.A(n_1257),
.Y(n_1431)
);

CKINVDCx11_ASAP7_75t_R g1432 ( 
.A(n_1281),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1305),
.A2(n_1329),
.B1(n_1368),
.B2(n_1315),
.Y(n_1433)
);

BUFx8_ASAP7_75t_SL g1434 ( 
.A(n_1285),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1290),
.A2(n_1292),
.B1(n_1362),
.B2(n_1379),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1290),
.A2(n_1379),
.B1(n_1362),
.B2(n_1267),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1361),
.B(n_1240),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1345),
.A2(n_1353),
.B1(n_1307),
.B2(n_1354),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1299),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1357),
.B(n_1255),
.Y(n_1440)
);

INVx8_ASAP7_75t_L g1441 ( 
.A(n_1307),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1354),
.A2(n_1383),
.B1(n_1370),
.B2(n_1365),
.Y(n_1442)
);

CKINVDCx11_ASAP7_75t_R g1443 ( 
.A(n_1333),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1270),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1277),
.A2(n_1293),
.B1(n_1260),
.B2(n_1254),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_1294),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1302),
.A2(n_1366),
.B1(n_1284),
.B2(n_1263),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1282),
.A2(n_1258),
.B1(n_1280),
.B2(n_1261),
.Y(n_1448)
);

BUFx6f_ASAP7_75t_L g1449 ( 
.A(n_1237),
.Y(n_1449)
);

INVx6_ASAP7_75t_L g1450 ( 
.A(n_1295),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1251),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1316),
.A2(n_1289),
.B1(n_1369),
.B2(n_1359),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1316),
.A2(n_1338),
.B1(n_1355),
.B2(n_1318),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1300),
.B(n_1380),
.Y(n_1454)
);

CKINVDCx6p67_ASAP7_75t_R g1455 ( 
.A(n_1304),
.Y(n_1455)
);

INVx4_ASAP7_75t_L g1456 ( 
.A(n_1297),
.Y(n_1456)
);

BUFx12f_ASAP7_75t_L g1457 ( 
.A(n_1317),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1228),
.Y(n_1458)
);

CKINVDCx14_ASAP7_75t_R g1459 ( 
.A(n_1301),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1300),
.A2(n_1380),
.B1(n_1278),
.B2(n_1346),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1300),
.B(n_1380),
.Y(n_1461)
);

BUFx8_ASAP7_75t_L g1462 ( 
.A(n_1237),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1242),
.A2(n_1342),
.B1(n_1321),
.B2(n_1245),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1269),
.A2(n_1237),
.B1(n_1275),
.B2(n_1286),
.Y(n_1464)
);

BUFx3_ASAP7_75t_L g1465 ( 
.A(n_1337),
.Y(n_1465)
);

CKINVDCx12_ASAP7_75t_R g1466 ( 
.A(n_1288),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_SL g1467 ( 
.A1(n_1337),
.A2(n_1377),
.B1(n_1349),
.B2(n_1252),
.Y(n_1467)
);

AOI22xp5_ASAP7_75t_SL g1468 ( 
.A1(n_1349),
.A2(n_1377),
.B1(n_1241),
.B2(n_1252),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1377),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1232),
.A2(n_1325),
.B1(n_1344),
.B2(n_1306),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1241),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1308),
.A2(n_1328),
.B1(n_1334),
.B2(n_1374),
.Y(n_1472)
);

AOI22xp5_ASAP7_75t_SL g1473 ( 
.A1(n_1252),
.A2(n_1343),
.B1(n_1358),
.B2(n_1323),
.Y(n_1473)
);

INVx1_ASAP7_75t_SL g1474 ( 
.A(n_1266),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1235),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1351),
.A2(n_937),
.B1(n_795),
.B2(n_1336),
.Y(n_1476)
);

OAI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1323),
.A2(n_937),
.B(n_998),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1235),
.Y(n_1478)
);

CKINVDCx6p67_ASAP7_75t_R g1479 ( 
.A(n_1265),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1351),
.A2(n_937),
.B1(n_795),
.B2(n_1336),
.Y(n_1480)
);

OAI21xp33_ASAP7_75t_L g1481 ( 
.A1(n_1351),
.A2(n_937),
.B(n_1206),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1351),
.A2(n_937),
.B1(n_795),
.B2(n_1336),
.Y(n_1482)
);

CKINVDCx11_ASAP7_75t_R g1483 ( 
.A(n_1231),
.Y(n_1483)
);

CKINVDCx20_ASAP7_75t_R g1484 ( 
.A(n_1367),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_1330),
.Y(n_1485)
);

INVx3_ASAP7_75t_SL g1486 ( 
.A(n_1330),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1351),
.A2(n_937),
.B1(n_795),
.B2(n_1336),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1248),
.B(n_1276),
.Y(n_1488)
);

BUFx12f_ASAP7_75t_L g1489 ( 
.A(n_1330),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1351),
.A2(n_937),
.B1(n_795),
.B2(n_1336),
.Y(n_1490)
);

INVx6_ASAP7_75t_L g1491 ( 
.A(n_1331),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1312),
.Y(n_1492)
);

INVx8_ASAP7_75t_L g1493 ( 
.A(n_1266),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1248),
.B(n_1276),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1235),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1235),
.Y(n_1496)
);

BUFx3_ASAP7_75t_L g1497 ( 
.A(n_1243),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1351),
.A2(n_937),
.B1(n_795),
.B2(n_1336),
.Y(n_1498)
);

BUFx2_ASAP7_75t_SL g1499 ( 
.A(n_1367),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1351),
.A2(n_937),
.B1(n_795),
.B2(n_1336),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1330),
.Y(n_1501)
);

INVx6_ASAP7_75t_L g1502 ( 
.A(n_1331),
.Y(n_1502)
);

INVx8_ASAP7_75t_L g1503 ( 
.A(n_1266),
.Y(n_1503)
);

AOI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1323),
.A2(n_1203),
.B1(n_937),
.B2(n_1343),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1351),
.A2(n_937),
.B1(n_795),
.B2(n_1336),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1312),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1351),
.A2(n_937),
.B1(n_795),
.B2(n_1336),
.Y(n_1507)
);

BUFx10_ASAP7_75t_L g1508 ( 
.A(n_1330),
.Y(n_1508)
);

INVx1_ASAP7_75t_SL g1509 ( 
.A(n_1266),
.Y(n_1509)
);

INVxp67_ASAP7_75t_SL g1510 ( 
.A(n_1287),
.Y(n_1510)
);

INVx2_ASAP7_75t_SL g1511 ( 
.A(n_1266),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1243),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1351),
.A2(n_937),
.B1(n_795),
.B2(n_1336),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1351),
.A2(n_937),
.B1(n_795),
.B2(n_1336),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_SL g1515 ( 
.A1(n_1407),
.A2(n_1504),
.B1(n_1409),
.B2(n_1392),
.Y(n_1515)
);

INVx4_ASAP7_75t_L g1516 ( 
.A(n_1457),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1439),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1404),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1449),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1454),
.B(n_1461),
.Y(n_1520)
);

OAI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1396),
.A2(n_1407),
.B(n_1386),
.Y(n_1521)
);

OAI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1396),
.A2(n_1386),
.B(n_1477),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1492),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1465),
.B(n_1449),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1506),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1449),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1459),
.A2(n_1462),
.B1(n_1481),
.B2(n_1384),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1471),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1449),
.B(n_1400),
.Y(n_1529)
);

OAI21x1_ASAP7_75t_L g1530 ( 
.A1(n_1452),
.A2(n_1453),
.B(n_1470),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1465),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1390),
.B(n_1397),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1458),
.Y(n_1533)
);

OA21x2_ASAP7_75t_L g1534 ( 
.A1(n_1463),
.A2(n_1464),
.B(n_1460),
.Y(n_1534)
);

O2A1O1Ixp33_ASAP7_75t_SL g1535 ( 
.A1(n_1440),
.A2(n_1433),
.B(n_1437),
.C(n_1451),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1401),
.B(n_1402),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1405),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1412),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1469),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1413),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1467),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1423),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1475),
.Y(n_1543)
);

INVx4_ASAP7_75t_SL g1544 ( 
.A(n_1385),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1421),
.B(n_1415),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1473),
.B(n_1410),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1478),
.Y(n_1547)
);

OA21x2_ASAP7_75t_L g1548 ( 
.A1(n_1463),
.A2(n_1464),
.B(n_1460),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1495),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1496),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1468),
.B(n_1445),
.Y(n_1551)
);

AOI21x1_ASAP7_75t_L g1552 ( 
.A1(n_1447),
.A2(n_1448),
.B(n_1387),
.Y(n_1552)
);

AOI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1488),
.A2(n_1494),
.B(n_1466),
.Y(n_1553)
);

INVx1_ASAP7_75t_SL g1554 ( 
.A(n_1446),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1414),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1388),
.Y(n_1556)
);

OA21x2_ASAP7_75t_L g1557 ( 
.A1(n_1470),
.A2(n_1472),
.B(n_1445),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1459),
.B(n_1416),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1510),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1497),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1450),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1416),
.B(n_1436),
.Y(n_1562)
);

INVx3_ASAP7_75t_L g1563 ( 
.A(n_1456),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1450),
.Y(n_1564)
);

OAI21x1_ASAP7_75t_L g1565 ( 
.A1(n_1472),
.A2(n_1444),
.B(n_1438),
.Y(n_1565)
);

INVx3_ASAP7_75t_L g1566 ( 
.A(n_1457),
.Y(n_1566)
);

BUFx8_ASAP7_75t_SL g1567 ( 
.A(n_1428),
.Y(n_1567)
);

OAI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1476),
.A2(n_1514),
.B1(n_1513),
.B2(n_1480),
.Y(n_1568)
);

AOI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1410),
.A2(n_1490),
.B(n_1513),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1436),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1424),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1424),
.Y(n_1572)
);

A2O1A1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1476),
.A2(n_1514),
.B(n_1507),
.C(n_1505),
.Y(n_1573)
);

INVx3_ASAP7_75t_L g1574 ( 
.A(n_1455),
.Y(n_1574)
);

INVx1_ASAP7_75t_SL g1575 ( 
.A(n_1512),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1422),
.B(n_1498),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1389),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1389),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1480),
.B(n_1490),
.Y(n_1579)
);

OAI21x1_ASAP7_75t_L g1580 ( 
.A1(n_1422),
.A2(n_1435),
.B(n_1398),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1398),
.Y(n_1581)
);

INVx3_ASAP7_75t_L g1582 ( 
.A(n_1403),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1403),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1482),
.B(n_1500),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1482),
.A2(n_1500),
.B1(n_1507),
.B2(n_1487),
.Y(n_1585)
);

AO31x2_ASAP7_75t_L g1586 ( 
.A1(n_1419),
.A2(n_1435),
.A3(n_1505),
.B(n_1487),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1498),
.B(n_1426),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1484),
.B(n_1474),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1483),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1417),
.B(n_1408),
.Y(n_1590)
);

BUFx2_ASAP7_75t_L g1591 ( 
.A(n_1408),
.Y(n_1591)
);

BUFx2_ASAP7_75t_L g1592 ( 
.A(n_1434),
.Y(n_1592)
);

OAI21x1_ASAP7_75t_L g1593 ( 
.A1(n_1442),
.A2(n_1491),
.B(n_1502),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_L g1594 ( 
.A(n_1484),
.B(n_1509),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1395),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1395),
.Y(n_1596)
);

OAI21xp5_ASAP7_75t_L g1597 ( 
.A1(n_1511),
.A2(n_1429),
.B(n_1394),
.Y(n_1597)
);

OAI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1522),
.A2(n_1420),
.B(n_1406),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1538),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1529),
.B(n_1520),
.Y(n_1600)
);

OA21x2_ASAP7_75t_L g1601 ( 
.A1(n_1530),
.A2(n_1418),
.B(n_1411),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_1524),
.B(n_1519),
.Y(n_1602)
);

NOR2x1_ASAP7_75t_SL g1603 ( 
.A(n_1553),
.B(n_1552),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1515),
.B(n_1535),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1520),
.B(n_1394),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1518),
.B(n_1427),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1524),
.B(n_1519),
.Y(n_1607)
);

OAI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1522),
.A2(n_1420),
.B(n_1427),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1575),
.B(n_1430),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1575),
.B(n_1430),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1542),
.Y(n_1611)
);

OA21x2_ASAP7_75t_L g1612 ( 
.A1(n_1530),
.A2(n_1441),
.B(n_1485),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1556),
.B(n_1430),
.Y(n_1613)
);

AOI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1515),
.A2(n_1431),
.B1(n_1428),
.B2(n_1479),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1523),
.B(n_1503),
.Y(n_1615)
);

OR2x6_ASAP7_75t_L g1616 ( 
.A(n_1593),
.B(n_1503),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1552),
.B(n_1432),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1526),
.B(n_1551),
.Y(n_1618)
);

NAND2xp33_ASAP7_75t_SL g1619 ( 
.A(n_1574),
.B(n_1486),
.Y(n_1619)
);

OAI21xp5_ASAP7_75t_L g1620 ( 
.A1(n_1521),
.A2(n_1393),
.B(n_1501),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1551),
.B(n_1499),
.Y(n_1621)
);

AOI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1521),
.A2(n_1503),
.B(n_1399),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1532),
.B(n_1486),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1560),
.B(n_1443),
.Y(n_1624)
);

OAI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1585),
.A2(n_1399),
.B1(n_1493),
.B2(n_1489),
.Y(n_1625)
);

NOR2x1_ASAP7_75t_SL g1626 ( 
.A(n_1553),
.B(n_1489),
.Y(n_1626)
);

AO32x2_ASAP7_75t_L g1627 ( 
.A1(n_1568),
.A2(n_1399),
.A3(n_1493),
.B1(n_1443),
.B2(n_1483),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1525),
.B(n_1493),
.Y(n_1628)
);

OAI21x1_ASAP7_75t_SL g1629 ( 
.A1(n_1516),
.A2(n_1425),
.B(n_1391),
.Y(n_1629)
);

O2A1O1Ixp33_ASAP7_75t_L g1630 ( 
.A1(n_1546),
.A2(n_1391),
.B(n_1508),
.C(n_1425),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1517),
.B(n_1508),
.Y(n_1631)
);

A2O1A1Ixp33_ASAP7_75t_L g1632 ( 
.A1(n_1569),
.A2(n_1573),
.B(n_1527),
.C(n_1568),
.Y(n_1632)
);

A2O1A1Ixp33_ASAP7_75t_L g1633 ( 
.A1(n_1569),
.A2(n_1579),
.B(n_1584),
.C(n_1576),
.Y(n_1633)
);

OAI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1545),
.A2(n_1576),
.B(n_1584),
.Y(n_1634)
);

O2A1O1Ixp33_ASAP7_75t_L g1635 ( 
.A1(n_1579),
.A2(n_1554),
.B(n_1541),
.C(n_1574),
.Y(n_1635)
);

AOI21x1_ASAP7_75t_L g1636 ( 
.A1(n_1597),
.A2(n_1564),
.B(n_1561),
.Y(n_1636)
);

O2A1O1Ixp33_ASAP7_75t_SL g1637 ( 
.A1(n_1574),
.A2(n_1566),
.B(n_1596),
.C(n_1595),
.Y(n_1637)
);

OA21x2_ASAP7_75t_L g1638 ( 
.A1(n_1565),
.A2(n_1580),
.B(n_1541),
.Y(n_1638)
);

OAI22xp5_ASAP7_75t_SL g1639 ( 
.A1(n_1589),
.A2(n_1592),
.B1(n_1516),
.B2(n_1554),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1537),
.B(n_1540),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1532),
.B(n_1536),
.Y(n_1641)
);

A2O1A1Ixp33_ASAP7_75t_L g1642 ( 
.A1(n_1558),
.A2(n_1562),
.B(n_1587),
.C(n_1580),
.Y(n_1642)
);

A2O1A1Ixp33_ASAP7_75t_L g1643 ( 
.A1(n_1558),
.A2(n_1562),
.B(n_1580),
.C(n_1541),
.Y(n_1643)
);

AO21x2_ASAP7_75t_L g1644 ( 
.A1(n_1571),
.A2(n_1572),
.B(n_1590),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1543),
.B(n_1547),
.Y(n_1645)
);

INVx2_ASAP7_75t_SL g1646 ( 
.A(n_1578),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1574),
.B(n_1566),
.Y(n_1647)
);

O2A1O1Ixp33_ASAP7_75t_L g1648 ( 
.A1(n_1597),
.A2(n_1566),
.B(n_1577),
.C(n_1583),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1531),
.B(n_1544),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1549),
.B(n_1550),
.Y(n_1650)
);

AO32x2_ASAP7_75t_L g1651 ( 
.A1(n_1570),
.A2(n_1559),
.A3(n_1555),
.B1(n_1534),
.B2(n_1548),
.Y(n_1651)
);

BUFx8_ASAP7_75t_L g1652 ( 
.A(n_1567),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1599),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1641),
.B(n_1534),
.Y(n_1654)
);

NAND4xp25_ASAP7_75t_L g1655 ( 
.A(n_1604),
.B(n_1594),
.C(n_1588),
.D(n_1566),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1600),
.B(n_1557),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1611),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1646),
.Y(n_1658)
);

BUFx2_ASAP7_75t_L g1659 ( 
.A(n_1612),
.Y(n_1659)
);

BUFx2_ASAP7_75t_L g1660 ( 
.A(n_1612),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1618),
.B(n_1548),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1640),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1618),
.B(n_1548),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1612),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1650),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1632),
.A2(n_1577),
.B1(n_1581),
.B2(n_1583),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1645),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1617),
.B(n_1582),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1638),
.Y(n_1669)
);

BUFx2_ASAP7_75t_L g1670 ( 
.A(n_1601),
.Y(n_1670)
);

BUFx2_ASAP7_75t_L g1671 ( 
.A(n_1601),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1651),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1642),
.B(n_1528),
.Y(n_1673)
);

INVxp67_ASAP7_75t_SL g1674 ( 
.A(n_1601),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1604),
.A2(n_1539),
.B1(n_1586),
.B2(n_1533),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1649),
.B(n_1563),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1651),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1636),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_SL g1679 ( 
.A1(n_1614),
.A2(n_1539),
.B1(n_1591),
.B2(n_1581),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1642),
.B(n_1528),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1657),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1656),
.B(n_1605),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1669),
.Y(n_1683)
);

INVx3_ASAP7_75t_L g1684 ( 
.A(n_1664),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1672),
.B(n_1654),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1656),
.B(n_1643),
.Y(n_1686)
);

INVx1_ASAP7_75t_SL g1687 ( 
.A(n_1653),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1655),
.B(n_1621),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1656),
.B(n_1643),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1669),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1653),
.Y(n_1691)
);

INVx4_ASAP7_75t_L g1692 ( 
.A(n_1676),
.Y(n_1692)
);

INVxp33_ASAP7_75t_L g1693 ( 
.A(n_1655),
.Y(n_1693)
);

AOI33xp33_ASAP7_75t_L g1694 ( 
.A1(n_1672),
.A2(n_1621),
.A3(n_1635),
.B1(n_1637),
.B2(n_1623),
.B3(n_1630),
.Y(n_1694)
);

BUFx2_ASAP7_75t_L g1695 ( 
.A(n_1664),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1657),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1654),
.B(n_1644),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1656),
.B(n_1623),
.Y(n_1698)
);

NAND4xp25_ASAP7_75t_L g1699 ( 
.A(n_1655),
.B(n_1620),
.C(n_1632),
.D(n_1606),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1654),
.B(n_1633),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1672),
.B(n_1633),
.Y(n_1701)
);

A2O1A1Ixp33_ASAP7_75t_SL g1702 ( 
.A1(n_1668),
.A2(n_1608),
.B(n_1647),
.C(n_1598),
.Y(n_1702)
);

BUFx2_ASAP7_75t_L g1703 ( 
.A(n_1664),
.Y(n_1703)
);

NOR2x1_ASAP7_75t_L g1704 ( 
.A(n_1666),
.B(n_1631),
.Y(n_1704)
);

INVx4_ASAP7_75t_L g1705 ( 
.A(n_1676),
.Y(n_1705)
);

OAI33xp33_ASAP7_75t_L g1706 ( 
.A1(n_1666),
.A2(n_1639),
.A3(n_1625),
.B1(n_1615),
.B2(n_1628),
.B3(n_1648),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1658),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1661),
.B(n_1602),
.Y(n_1708)
);

OR2x2_ASAP7_75t_SL g1709 ( 
.A(n_1677),
.B(n_1678),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1661),
.B(n_1607),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1665),
.B(n_1603),
.Y(n_1711)
);

AND2x2_ASAP7_75t_SL g1712 ( 
.A(n_1673),
.B(n_1649),
.Y(n_1712)
);

INVxp67_ASAP7_75t_L g1713 ( 
.A(n_1711),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1701),
.B(n_1665),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1708),
.B(n_1661),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1708),
.B(n_1661),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1691),
.Y(n_1717)
);

NOR2xp67_ASAP7_75t_L g1718 ( 
.A(n_1692),
.B(n_1705),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1691),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1701),
.B(n_1665),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1696),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1696),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1696),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1701),
.B(n_1677),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1692),
.B(n_1674),
.Y(n_1725)
);

HB1xp67_ASAP7_75t_L g1726 ( 
.A(n_1707),
.Y(n_1726)
);

CKINVDCx20_ASAP7_75t_R g1727 ( 
.A(n_1688),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1685),
.B(n_1677),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1687),
.B(n_1677),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1692),
.B(n_1674),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1683),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1708),
.B(n_1663),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1687),
.B(n_1662),
.Y(n_1733)
);

AOI22xp5_ASAP7_75t_L g1734 ( 
.A1(n_1693),
.A2(n_1675),
.B1(n_1634),
.B2(n_1680),
.Y(n_1734)
);

BUFx3_ASAP7_75t_L g1735 ( 
.A(n_1709),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1685),
.B(n_1662),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1700),
.B(n_1709),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1710),
.B(n_1663),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1704),
.B(n_1667),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1704),
.B(n_1667),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1683),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1683),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1710),
.B(n_1663),
.Y(n_1743)
);

INVxp67_ASAP7_75t_SL g1744 ( 
.A(n_1683),
.Y(n_1744)
);

BUFx3_ASAP7_75t_L g1745 ( 
.A(n_1709),
.Y(n_1745)
);

INVx3_ASAP7_75t_L g1746 ( 
.A(n_1692),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1698),
.B(n_1659),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1690),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1681),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1690),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1714),
.B(n_1693),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1715),
.B(n_1698),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1717),
.Y(n_1753)
);

BUFx2_ASAP7_75t_SL g1754 ( 
.A(n_1735),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1717),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1719),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1715),
.B(n_1698),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1719),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1726),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1726),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1714),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1713),
.Y(n_1762)
);

AND2x4_ASAP7_75t_L g1763 ( 
.A(n_1735),
.B(n_1692),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1737),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1724),
.B(n_1700),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1720),
.Y(n_1766)
);

AND2x4_ASAP7_75t_L g1767 ( 
.A(n_1735),
.B(n_1705),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1715),
.B(n_1705),
.Y(n_1768)
);

AND2x4_ASAP7_75t_L g1769 ( 
.A(n_1745),
.B(n_1705),
.Y(n_1769)
);

INVx2_ASAP7_75t_SL g1770 ( 
.A(n_1745),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1720),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1749),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1737),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1713),
.B(n_1694),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1737),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1716),
.B(n_1705),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1749),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1716),
.B(n_1682),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1721),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1724),
.B(n_1700),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1721),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1739),
.B(n_1694),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1739),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1722),
.Y(n_1784)
);

NAND4xp25_ASAP7_75t_L g1785 ( 
.A(n_1745),
.B(n_1702),
.C(n_1699),
.D(n_1703),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1722),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1731),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1723),
.Y(n_1788)
);

AOI211xp5_ASAP7_75t_L g1789 ( 
.A1(n_1740),
.A2(n_1706),
.B(n_1699),
.C(n_1702),
.Y(n_1789)
);

HB1xp67_ASAP7_75t_L g1790 ( 
.A(n_1740),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1716),
.B(n_1682),
.Y(n_1791)
);

OR2x2_ASAP7_75t_L g1792 ( 
.A(n_1736),
.B(n_1711),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_L g1793 ( 
.A(n_1727),
.B(n_1652),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1732),
.B(n_1682),
.Y(n_1794)
);

OR2x6_ASAP7_75t_L g1795 ( 
.A(n_1729),
.B(n_1616),
.Y(n_1795)
);

OAI211xp5_ASAP7_75t_SL g1796 ( 
.A1(n_1729),
.A2(n_1733),
.B(n_1734),
.C(n_1684),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1778),
.B(n_1732),
.Y(n_1797)
);

INVx1_ASAP7_75t_SL g1798 ( 
.A(n_1793),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1778),
.B(n_1732),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1791),
.B(n_1738),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1789),
.B(n_1686),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1791),
.B(n_1738),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1751),
.B(n_1686),
.Y(n_1803)
);

NAND2x1_ASAP7_75t_L g1804 ( 
.A(n_1769),
.B(n_1746),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1753),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1753),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1764),
.Y(n_1807)
);

AO211x2_ASAP7_75t_L g1808 ( 
.A1(n_1785),
.A2(n_1627),
.B(n_1706),
.C(n_1622),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1755),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1794),
.B(n_1738),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_L g1811 ( 
.A(n_1774),
.B(n_1652),
.Y(n_1811)
);

NOR2xp67_ASAP7_75t_L g1812 ( 
.A(n_1770),
.B(n_1746),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1762),
.B(n_1782),
.Y(n_1813)
);

AOI221xp5_ASAP7_75t_L g1814 ( 
.A1(n_1796),
.A2(n_1689),
.B1(n_1686),
.B2(n_1734),
.C(n_1744),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1755),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1794),
.B(n_1743),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1756),
.Y(n_1817)
);

INVx3_ASAP7_75t_L g1818 ( 
.A(n_1769),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1761),
.B(n_1689),
.Y(n_1819)
);

INVx1_ASAP7_75t_SL g1820 ( 
.A(n_1754),
.Y(n_1820)
);

NOR2xp33_ASAP7_75t_L g1821 ( 
.A(n_1765),
.B(n_1652),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1756),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1752),
.B(n_1743),
.Y(n_1823)
);

INVx1_ASAP7_75t_SL g1824 ( 
.A(n_1754),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1758),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1759),
.Y(n_1826)
);

HB1xp67_ASAP7_75t_L g1827 ( 
.A(n_1783),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1765),
.B(n_1736),
.Y(n_1828)
);

NOR3xp33_ASAP7_75t_L g1829 ( 
.A(n_1770),
.B(n_1744),
.C(n_1688),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1759),
.Y(n_1830)
);

INVxp67_ASAP7_75t_L g1831 ( 
.A(n_1790),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1758),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1760),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1760),
.Y(n_1834)
);

NAND2x1p5_ASAP7_75t_L g1835 ( 
.A(n_1820),
.B(n_1712),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1801),
.B(n_1764),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1813),
.B(n_1773),
.Y(n_1837)
);

OAI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1831),
.A2(n_1727),
.B(n_1773),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_L g1839 ( 
.A(n_1798),
.B(n_1780),
.Y(n_1839)
);

OAI22xp33_ASAP7_75t_L g1840 ( 
.A1(n_1814),
.A2(n_1780),
.B1(n_1775),
.B2(n_1795),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1805),
.Y(n_1841)
);

AND2x4_ASAP7_75t_L g1842 ( 
.A(n_1824),
.B(n_1775),
.Y(n_1842)
);

OAI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1803),
.A2(n_1819),
.B1(n_1795),
.B2(n_1689),
.Y(n_1843)
);

AOI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1808),
.A2(n_1675),
.B1(n_1795),
.B2(n_1659),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1805),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1828),
.B(n_1792),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1827),
.B(n_1761),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1806),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1806),
.Y(n_1849)
);

NOR4xp25_ASAP7_75t_SL g1850 ( 
.A(n_1826),
.B(n_1703),
.C(n_1695),
.D(n_1766),
.Y(n_1850)
);

AOI31xp33_ASAP7_75t_L g1851 ( 
.A1(n_1811),
.A2(n_1769),
.A3(n_1763),
.B(n_1767),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1808),
.B(n_1766),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1809),
.Y(n_1853)
);

XNOR2xp5_ASAP7_75t_L g1854 ( 
.A(n_1829),
.B(n_1712),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1809),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1818),
.Y(n_1856)
);

OAI221xp5_ASAP7_75t_L g1857 ( 
.A1(n_1807),
.A2(n_1795),
.B1(n_1728),
.B2(n_1771),
.C(n_1697),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1807),
.B(n_1771),
.Y(n_1858)
);

INVx1_ASAP7_75t_SL g1859 ( 
.A(n_1821),
.Y(n_1859)
);

AOI21xp33_ASAP7_75t_L g1860 ( 
.A1(n_1833),
.A2(n_1777),
.B(n_1772),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1815),
.Y(n_1861)
);

AOI211xp5_ASAP7_75t_L g1862 ( 
.A1(n_1852),
.A2(n_1817),
.B(n_1822),
.C(n_1815),
.Y(n_1862)
);

OAI221xp5_ASAP7_75t_L g1863 ( 
.A1(n_1844),
.A2(n_1828),
.B1(n_1728),
.B2(n_1818),
.C(n_1812),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1839),
.B(n_1830),
.Y(n_1864)
);

OAI221xp5_ASAP7_75t_L g1865 ( 
.A1(n_1852),
.A2(n_1728),
.B1(n_1818),
.B2(n_1832),
.C(n_1825),
.Y(n_1865)
);

AOI221xp5_ASAP7_75t_L g1866 ( 
.A1(n_1840),
.A2(n_1822),
.B1(n_1817),
.B2(n_1832),
.C(n_1825),
.Y(n_1866)
);

OAI21xp5_ASAP7_75t_SL g1867 ( 
.A1(n_1851),
.A2(n_1769),
.B(n_1767),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1835),
.Y(n_1868)
);

OAI222xp33_ASAP7_75t_L g1869 ( 
.A1(n_1836),
.A2(n_1834),
.B1(n_1833),
.B2(n_1697),
.C1(n_1671),
.C2(n_1670),
.Y(n_1869)
);

AOI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1850),
.A2(n_1804),
.B(n_1834),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1846),
.B(n_1792),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1842),
.B(n_1797),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1841),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1842),
.B(n_1797),
.Y(n_1874)
);

OAI221xp5_ASAP7_75t_L g1875 ( 
.A1(n_1835),
.A2(n_1660),
.B1(n_1659),
.B2(n_1670),
.C(n_1671),
.Y(n_1875)
);

AOI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1838),
.A2(n_1660),
.B1(n_1671),
.B2(n_1670),
.Y(n_1876)
);

OAI31xp33_ASAP7_75t_L g1877 ( 
.A1(n_1857),
.A2(n_1660),
.A3(n_1697),
.B(n_1678),
.Y(n_1877)
);

INVxp33_ASAP7_75t_L g1878 ( 
.A(n_1838),
.Y(n_1878)
);

OAI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1854),
.A2(n_1800),
.B1(n_1802),
.B2(n_1799),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1845),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1848),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1856),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1871),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1872),
.Y(n_1884)
);

NAND2x1_ASAP7_75t_L g1885 ( 
.A(n_1868),
.B(n_1849),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1878),
.B(n_1859),
.Y(n_1886)
);

INVx1_ASAP7_75t_SL g1887 ( 
.A(n_1874),
.Y(n_1887)
);

O2A1O1Ixp33_ASAP7_75t_L g1888 ( 
.A1(n_1878),
.A2(n_1837),
.B(n_1847),
.C(n_1860),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1882),
.Y(n_1889)
);

AOI222xp33_ASAP7_75t_L g1890 ( 
.A1(n_1865),
.A2(n_1863),
.B1(n_1869),
.B2(n_1866),
.C1(n_1864),
.C2(n_1882),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1881),
.Y(n_1891)
);

INVxp67_ASAP7_75t_L g1892 ( 
.A(n_1873),
.Y(n_1892)
);

AOI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1870),
.A2(n_1860),
.B(n_1858),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1867),
.B(n_1799),
.Y(n_1894)
);

NOR2xp33_ASAP7_75t_L g1895 ( 
.A(n_1886),
.B(n_1879),
.Y(n_1895)
);

AOI211x1_ASAP7_75t_L g1896 ( 
.A1(n_1893),
.A2(n_1869),
.B(n_1843),
.C(n_1875),
.Y(n_1896)
);

NOR3xp33_ASAP7_75t_L g1897 ( 
.A(n_1886),
.B(n_1862),
.C(n_1880),
.Y(n_1897)
);

OAI21xp5_ASAP7_75t_SL g1898 ( 
.A1(n_1890),
.A2(n_1876),
.B(n_1877),
.Y(n_1898)
);

AO21x1_ASAP7_75t_L g1899 ( 
.A1(n_1888),
.A2(n_1855),
.B(n_1853),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1889),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1887),
.B(n_1861),
.Y(n_1901)
);

NAND2x1_ASAP7_75t_L g1902 ( 
.A(n_1883),
.B(n_1763),
.Y(n_1902)
);

OAI21xp5_ASAP7_75t_L g1903 ( 
.A1(n_1892),
.A2(n_1885),
.B(n_1894),
.Y(n_1903)
);

NAND3xp33_ASAP7_75t_L g1904 ( 
.A(n_1889),
.B(n_1804),
.C(n_1787),
.Y(n_1904)
);

BUFx2_ASAP7_75t_L g1905 ( 
.A(n_1894),
.Y(n_1905)
);

AOI22xp5_ASAP7_75t_L g1906 ( 
.A1(n_1898),
.A2(n_1884),
.B1(n_1891),
.B2(n_1787),
.Y(n_1906)
);

OAI321xp33_ASAP7_75t_L g1907 ( 
.A1(n_1903),
.A2(n_1891),
.A3(n_1679),
.B1(n_1816),
.B2(n_1810),
.C(n_1802),
.Y(n_1907)
);

OAI221xp5_ASAP7_75t_L g1908 ( 
.A1(n_1897),
.A2(n_1777),
.B1(n_1772),
.B2(n_1695),
.C(n_1703),
.Y(n_1908)
);

OAI222xp33_ASAP7_75t_L g1909 ( 
.A1(n_1905),
.A2(n_1763),
.B1(n_1767),
.B2(n_1810),
.C1(n_1800),
.C2(n_1816),
.Y(n_1909)
);

AOI21xp33_ASAP7_75t_SL g1910 ( 
.A1(n_1895),
.A2(n_1629),
.B(n_1823),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1896),
.B(n_1900),
.Y(n_1911)
);

AOI321xp33_ASAP7_75t_L g1912 ( 
.A1(n_1901),
.A2(n_1823),
.A3(n_1673),
.B1(n_1680),
.B2(n_1664),
.C(n_1730),
.Y(n_1912)
);

NOR2xp33_ASAP7_75t_SL g1913 ( 
.A(n_1909),
.B(n_1904),
.Y(n_1913)
);

AOI211xp5_ASAP7_75t_L g1914 ( 
.A1(n_1911),
.A2(n_1899),
.B(n_1902),
.C(n_1637),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1906),
.Y(n_1915)
);

AOI221xp5_ASAP7_75t_L g1916 ( 
.A1(n_1907),
.A2(n_1908),
.B1(n_1910),
.B2(n_1912),
.C(n_1788),
.Y(n_1916)
);

AOI221xp5_ASAP7_75t_L g1917 ( 
.A1(n_1911),
.A2(n_1788),
.B1(n_1786),
.B2(n_1784),
.C(n_1781),
.Y(n_1917)
);

NAND4xp75_ASAP7_75t_L g1918 ( 
.A(n_1911),
.B(n_1712),
.C(n_1718),
.D(n_1747),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1911),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1915),
.Y(n_1920)
);

NOR2x1_ASAP7_75t_L g1921 ( 
.A(n_1919),
.B(n_1779),
.Y(n_1921)
);

OAI22xp5_ASAP7_75t_L g1922 ( 
.A1(n_1914),
.A2(n_1786),
.B1(n_1784),
.B2(n_1781),
.Y(n_1922)
);

NOR2x1_ASAP7_75t_L g1923 ( 
.A(n_1918),
.B(n_1913),
.Y(n_1923)
);

NAND4xp75_ASAP7_75t_L g1924 ( 
.A(n_1916),
.B(n_1712),
.C(n_1718),
.D(n_1610),
.Y(n_1924)
);

NOR2x1_ASAP7_75t_L g1925 ( 
.A(n_1917),
.B(n_1779),
.Y(n_1925)
);

OR2x6_ASAP7_75t_L g1926 ( 
.A(n_1923),
.B(n_1624),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1921),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1924),
.B(n_1695),
.Y(n_1928)
);

AOI31xp33_ASAP7_75t_L g1929 ( 
.A1(n_1920),
.A2(n_1619),
.A3(n_1768),
.B(n_1776),
.Y(n_1929)
);

XOR2xp5_ASAP7_75t_L g1930 ( 
.A(n_1927),
.B(n_1922),
.Y(n_1930)
);

AO22x2_ASAP7_75t_L g1931 ( 
.A1(n_1930),
.A2(n_1928),
.B1(n_1926),
.B2(n_1925),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1931),
.Y(n_1932)
);

XOR2xp5_ASAP7_75t_L g1933 ( 
.A(n_1931),
.B(n_1626),
.Y(n_1933)
);

OAI22xp5_ASAP7_75t_SL g1934 ( 
.A1(n_1932),
.A2(n_1929),
.B1(n_1725),
.B2(n_1730),
.Y(n_1934)
);

OAI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1933),
.A2(n_1733),
.B1(n_1752),
.B2(n_1757),
.Y(n_1935)
);

XNOR2x1_ASAP7_75t_L g1936 ( 
.A(n_1935),
.B(n_1609),
.Y(n_1936)
);

AOI22xp33_ASAP7_75t_L g1937 ( 
.A1(n_1934),
.A2(n_1741),
.B1(n_1742),
.B2(n_1731),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1936),
.Y(n_1938)
);

OR2x6_ASAP7_75t_L g1939 ( 
.A(n_1938),
.B(n_1937),
.Y(n_1939)
);

AOI21xp5_ASAP7_75t_L g1940 ( 
.A1(n_1939),
.A2(n_1741),
.B(n_1731),
.Y(n_1940)
);

AOI221xp5_ASAP7_75t_L g1941 ( 
.A1(n_1940),
.A2(n_1741),
.B1(n_1750),
.B2(n_1748),
.C(n_1742),
.Y(n_1941)
);

AOI211xp5_ASAP7_75t_L g1942 ( 
.A1(n_1941),
.A2(n_1619),
.B(n_1647),
.C(n_1613),
.Y(n_1942)
);


endmodule