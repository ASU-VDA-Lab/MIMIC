module fake_jpeg_13276_n_316 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_316);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_316;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g131 ( 
.A(n_47),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_49),
.Y(n_117)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_52),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_53),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_57),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_22),
.B(n_10),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_60),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_10),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_59),
.B(n_45),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_17),
.B(n_10),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_22),
.B(n_7),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_61),
.B(n_67),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_24),
.B(n_7),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_19),
.B(n_11),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_68),
.B(n_73),
.Y(n_110)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_39),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_72),
.B(n_76),
.Y(n_127)
);

INVx6_ASAP7_75t_SL g73 ( 
.A(n_39),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

BUFx10_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_24),
.B(n_11),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_78),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_80),
.Y(n_120)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_82),
.Y(n_121)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_30),
.B(n_6),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_84),
.Y(n_126)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_86),
.Y(n_124)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_88),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_39),
.Y(n_88)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_SL g132 ( 
.A1(n_89),
.A2(n_0),
.B(n_2),
.Y(n_132)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_90),
.B(n_5),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_91),
.B(n_106),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_62),
.A2(n_28),
.B1(n_25),
.B2(n_41),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_95),
.A2(n_99),
.B1(n_114),
.B2(n_128),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_48),
.A2(n_25),
.B1(n_28),
.B2(n_34),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_96),
.A2(n_135),
.B1(n_122),
.B2(n_121),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_65),
.A2(n_34),
.B1(n_41),
.B2(n_29),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_97),
.B(n_129),
.C(n_103),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_62),
.A2(n_18),
.B1(n_40),
.B2(n_33),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_101),
.B(n_91),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_60),
.B(n_33),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_20),
.C(n_46),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_122),
.C(n_129),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_40),
.B1(n_45),
.B2(n_30),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_112),
.A2(n_123),
.B1(n_134),
.B2(n_100),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_76),
.A2(n_40),
.B1(n_20),
.B2(n_46),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_63),
.A2(n_23),
.B1(n_38),
.B2(n_27),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_115),
.A2(n_119),
.B1(n_141),
.B2(n_117),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_82),
.A2(n_42),
.B1(n_38),
.B2(n_27),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_75),
.A2(n_42),
.B1(n_12),
.B2(n_3),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_55),
.A2(n_5),
.B1(n_14),
.B2(n_15),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_56),
.A2(n_74),
.B1(n_71),
.B2(n_84),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_89),
.A2(n_5),
.B1(n_14),
.B2(n_15),
.Y(n_129)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_132),
.A2(n_141),
.B1(n_115),
.B2(n_92),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_64),
.A2(n_15),
.B1(n_16),
.B2(n_0),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_51),
.A2(n_0),
.B1(n_2),
.B2(n_53),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_66),
.A2(n_70),
.B1(n_47),
.B2(n_72),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_120),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_142),
.B(n_146),
.Y(n_195)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_124),
.B1(n_97),
.B2(n_119),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_145),
.A2(n_161),
.B1(n_168),
.B2(n_174),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_147),
.B(n_153),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

INVx4_ASAP7_75t_SL g185 ( 
.A(n_148),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_106),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_172),
.C(n_175),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_127),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_150),
.B(n_158),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_93),
.B(n_98),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_154),
.Y(n_204)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_156),
.Y(n_197)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_107),
.Y(n_157)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_157),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_101),
.B(n_104),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_105),
.Y(n_159)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_160),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_118),
.A2(n_126),
.B1(n_109),
.B2(n_110),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_130),
.B(n_94),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_163),
.B(n_167),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_102),
.Y(n_164)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_94),
.Y(n_165)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_165),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_127),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_116),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_169),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_136),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_171),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_108),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_108),
.B(n_139),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_182),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_139),
.A2(n_137),
.B1(n_111),
.B2(n_125),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_113),
.B(n_116),
.C(n_138),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_111),
.A2(n_137),
.B1(n_125),
.B2(n_138),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_176),
.A2(n_178),
.B1(n_180),
.B2(n_169),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_100),
.B(n_117),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_175),
.C(n_171),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_117),
.A2(n_138),
.B1(n_113),
.B2(n_103),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_131),
.B(n_92),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_179),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_103),
.A2(n_121),
.B1(n_96),
.B2(n_124),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_103),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_181),
.Y(n_203)
);

O2A1O1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_145),
.A2(n_131),
.B(n_170),
.C(n_148),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_184),
.A2(n_190),
.B(n_204),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_182),
.A2(n_131),
.B(n_147),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_186),
.A2(n_152),
.B(n_157),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_173),
.A2(n_180),
.B(n_143),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_184),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_199),
.C(n_212),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_149),
.B(n_166),
.C(n_153),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_166),
.B(n_153),
.C(n_143),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_204),
.A2(n_168),
.B1(n_162),
.B2(n_153),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_213),
.A2(n_214),
.B1(n_219),
.B2(n_187),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_201),
.A2(n_172),
.B1(n_177),
.B2(n_156),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_215),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_210),
.B(n_165),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_229),
.Y(n_243)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_155),
.C(n_160),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_220),
.B(n_228),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_221),
.Y(n_240)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_222),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_181),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_224),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_183),
.B(n_164),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_202),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_227),
.Y(n_255)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_189),
.Y(n_226)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_226),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_194),
.Y(n_227)
);

MAJx2_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_188),
.C(n_212),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_188),
.B(n_192),
.C(n_186),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_208),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_232),
.Y(n_250)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_193),
.Y(n_231)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_192),
.B(n_201),
.C(n_190),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_196),
.B(n_193),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_235),
.Y(n_251)
);

OAI21xp33_ASAP7_75t_L g234 ( 
.A1(n_185),
.A2(n_196),
.B(n_209),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_234),
.A2(n_185),
.B(n_209),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_203),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_203),
.B(n_187),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_238),
.A2(n_247),
.B(n_230),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_236),
.A2(n_191),
.B1(n_205),
.B2(n_185),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_241),
.A2(n_249),
.B1(n_219),
.B2(n_214),
.Y(n_256)
);

XOR2x1_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_208),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_220),
.Y(n_257)
);

OA22x2_ASAP7_75t_L g262 ( 
.A1(n_245),
.A2(n_213),
.B1(n_219),
.B2(n_221),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_227),
.A2(n_205),
.B1(n_197),
.B2(n_206),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_206),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_231),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_256),
.A2(n_268),
.B1(n_270),
.B2(n_251),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_243),
.Y(n_278)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_239),
.Y(n_258)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_258),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_229),
.C(n_228),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_260),
.C(n_269),
.Y(n_277)
);

OAI322xp33_ASAP7_75t_L g260 ( 
.A1(n_255),
.A2(n_228),
.A3(n_224),
.B1(n_218),
.B2(n_233),
.C1(n_225),
.C2(n_223),
.Y(n_260)
);

NOR2x1_ASAP7_75t_SL g261 ( 
.A(n_238),
.B(n_218),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_261),
.Y(n_279)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_262),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_237),
.B(n_250),
.Y(n_274)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_264),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_265),
.B(n_266),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_187),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_252),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_271),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_241),
.A2(n_215),
.B1(n_226),
.B2(n_197),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_217),
.C(n_222),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_240),
.A2(n_247),
.B1(n_249),
.B2(n_245),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_207),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_267),
.A2(n_237),
.B1(n_242),
.B2(n_254),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_273),
.A2(n_282),
.B1(n_262),
.B2(n_264),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_274),
.A2(n_263),
.B(n_265),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_278),
.B(n_261),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_250),
.C(n_243),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_257),
.C(n_269),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_284),
.B(n_285),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_271),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_288),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_258),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_287),
.A2(n_291),
.B1(n_272),
.B2(n_276),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_262),
.C(n_270),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_292),
.C(n_280),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_279),
.A2(n_260),
.B(n_256),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_279),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_262),
.C(n_268),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_296),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_289),
.A2(n_272),
.B1(n_274),
.B2(n_281),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_294),
.A2(n_295),
.B1(n_293),
.B2(n_296),
.Y(n_300)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_288),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_248),
.C(n_254),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_304),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_295),
.A2(n_277),
.B(n_284),
.Y(n_301)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_301),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_294),
.A2(n_276),
.B1(n_283),
.B2(n_248),
.Y(n_303)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_303),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_303),
.A2(n_299),
.B1(n_244),
.B2(n_246),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_305),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_306),
.A2(n_302),
.B(n_308),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_311),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_305),
.A2(n_297),
.B(n_301),
.Y(n_311)
);

NAND2xp33_ASAP7_75t_R g313 ( 
.A(n_310),
.B(n_299),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_307),
.C(n_304),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_312),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_244),
.Y(n_316)
);


endmodule