module fake_jpeg_26216_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_4),
.B(n_5),
.Y(n_31)
);

BUFx4f_ASAP7_75t_SL g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_8),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_21),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_48),
.B(n_34),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_49),
.B(n_24),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_54),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

BUFx4f_ASAP7_75t_SL g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_61),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_31),
.B(n_33),
.Y(n_62)
);

NAND3xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_9),
.C(n_15),
.Y(n_86)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_67),
.Y(n_87)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_21),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_32),
.Y(n_116)
);

AO22x1_ASAP7_75t_SL g73 ( 
.A1(n_52),
.A2(n_47),
.B1(n_20),
.B2(n_17),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_73),
.A2(n_78),
.B1(n_95),
.B2(n_96),
.Y(n_106)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_75),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_66),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_81),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_50),
.A2(n_47),
.B1(n_43),
.B2(n_42),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_57),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_22),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_83),
.B(n_86),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_60),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_93),
.Y(n_121)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g93 ( 
.A(n_59),
.Y(n_93)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_50),
.A2(n_20),
.B1(n_29),
.B2(n_28),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_45),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_68),
.A2(n_20),
.B1(n_45),
.B2(n_40),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_54),
.A2(n_28),
.B1(n_23),
.B2(n_22),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_97),
.Y(n_120)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_99),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_72),
.A2(n_34),
.B(n_69),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_117),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_67),
.B1(n_64),
.B2(n_65),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_110),
.A2(n_114),
.B1(n_92),
.B2(n_76),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_111),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_73),
.A2(n_28),
.B1(n_23),
.B2(n_17),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_113),
.A2(n_123),
.B1(n_80),
.B2(n_92),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_73),
.A2(n_23),
.B1(n_69),
.B2(n_17),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_116),
.B(n_125),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_99),
.Y(n_117)
);

BUFx10_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_18),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_124),
.C(n_26),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_46),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_122),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_74),
.A2(n_24),
.B1(n_33),
.B2(n_19),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_78),
.B(n_95),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_126),
.B(n_76),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_83),
.B(n_32),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_107),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_112),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_128),
.B(n_129),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_108),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_130),
.Y(n_179)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_133),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_93),
.Y(n_133)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_138),
.Y(n_176)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

FAx1_ASAP7_75t_SL g140 ( 
.A(n_116),
.B(n_94),
.CI(n_98),
.CON(n_140),
.SN(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_122),
.B(n_106),
.C(n_100),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_143),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_85),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_99),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_146),
.A2(n_126),
.B1(n_125),
.B2(n_105),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_94),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_147),
.A2(n_27),
.B(n_30),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_112),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_148),
.B(n_152),
.Y(n_160)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_151),
.A2(n_156),
.B1(n_46),
.B2(n_71),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_85),
.Y(n_152)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_153),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_82),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_79),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_117),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_155),
.B(n_105),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_111),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_157),
.A2(n_162),
.B1(n_182),
.B2(n_188),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_119),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_159),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_106),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_161),
.A2(n_171),
.B(n_186),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_136),
.A2(n_122),
.B1(n_110),
.B2(n_100),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_172),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_147),
.A2(n_80),
.B1(n_104),
.B2(n_101),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_164),
.A2(n_167),
.B1(n_185),
.B2(n_187),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_104),
.B1(n_101),
.B2(n_79),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_134),
.C(n_136),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_180),
.C(n_184),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_35),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_137),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_134),
.B(n_145),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_175),
.B(n_178),
.Y(n_194)
);

AO21x1_ASAP7_75t_L g177 ( 
.A1(n_140),
.A2(n_26),
.B(n_36),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_181),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_145),
.B(n_19),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_35),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_71),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_131),
.A2(n_156),
.B1(n_140),
.B2(n_151),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_35),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_131),
.A2(n_46),
.B1(n_36),
.B2(n_18),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_128),
.A2(n_30),
.B1(n_102),
.B2(n_10),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_148),
.A2(n_155),
.B1(n_137),
.B2(n_144),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_160),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_191),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_163),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_193),
.Y(n_227)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_176),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_196),
.B(n_197),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_144),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_167),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_198),
.B(n_202),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_139),
.C(n_135),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_169),
.C(n_184),
.Y(n_232)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_164),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_203),
.B(n_209),
.Y(n_235)
);

AOI32xp33_ASAP7_75t_L g205 ( 
.A1(n_186),
.A2(n_161),
.A3(n_180),
.B1(n_168),
.B2(n_182),
.Y(n_205)
);

XNOR2x2_ASAP7_75t_SL g237 ( 
.A(n_205),
.B(n_207),
.Y(n_237)
);

INVxp33_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_211),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_144),
.Y(n_208)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_208),
.Y(n_222)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_175),
.Y(n_209)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_138),
.Y(n_212)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_212),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_149),
.Y(n_213)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_173),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_215),
.Y(n_240)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_217),
.Y(n_244)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_171),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_165),
.A2(n_132),
.B1(n_149),
.B2(n_30),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_219),
.A2(n_183),
.B1(n_132),
.B2(n_189),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_223),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_198),
.A2(n_159),
.B1(n_189),
.B2(n_170),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_SL g266 ( 
.A(n_226),
.B(n_237),
.C(n_238),
.Y(n_266)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_211),
.Y(n_228)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_231),
.Y(n_250)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_200),
.C(n_193),
.Y(n_262)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_208),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_243),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_242),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_218),
.A2(n_168),
.B1(n_177),
.B2(n_158),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_201),
.B(n_30),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_245),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_202),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_214),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_201),
.B(n_199),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_210),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_246)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_246),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_207),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_247),
.A2(n_226),
.B(n_206),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_245),
.B(n_204),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_254),
.Y(n_274)
);

FAx1_ASAP7_75t_SL g252 ( 
.A(n_223),
.B(n_199),
.CI(n_190),
.CON(n_252),
.SN(n_252)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_252),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_241),
.B(n_204),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_256),
.Y(n_279)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_239),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_235),
.Y(n_257)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_257),
.Y(n_275)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_236),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_260),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_210),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_2),
.Y(n_284)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_221),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_268),
.C(n_228),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_229),
.B(n_203),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_265),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_224),
.B(n_194),
.Y(n_267)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_267),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_196),
.C(n_218),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_268),
.A2(n_225),
.B1(n_234),
.B2(n_220),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_272),
.A2(n_278),
.B1(n_254),
.B2(n_259),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_266),
.A2(n_247),
.B1(n_246),
.B2(n_222),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_273),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_243),
.Y(n_276)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_276),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_266),
.A2(n_237),
.B1(n_244),
.B2(n_242),
.Y(n_278)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_280),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_248),
.Y(n_295)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_250),
.Y(n_282)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_282),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_1),
.Y(n_283)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_261),
.Y(n_290)
);

NAND3xp33_ASAP7_75t_L g285 ( 
.A(n_252),
.B(n_3),
.C(n_5),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_285),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_262),
.C(n_261),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_299),
.C(n_274),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_271),
.A2(n_253),
.B1(n_263),
.B2(n_251),
.Y(n_287)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

AO21x1_ASAP7_75t_L g289 ( 
.A1(n_280),
.A2(n_251),
.B(n_252),
.Y(n_289)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_294),
.Y(n_306)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_293),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_249),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_300),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_273),
.A2(n_6),
.B(n_7),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_296),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_278),
.C(n_276),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_269),
.Y(n_301)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_301),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_275),
.Y(n_303)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_303),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_274),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_7),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_292),
.A2(n_277),
.B1(n_279),
.B2(n_270),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_313),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_311),
.C(n_295),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_270),
.C(n_283),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_290),
.B(n_6),
.Y(n_313)
);

FAx1_ASAP7_75t_SL g314 ( 
.A(n_311),
.B(n_289),
.CI(n_294),
.CON(n_314),
.SN(n_314)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_314),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_317),
.B(n_318),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_312),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_307),
.A2(n_288),
.B1(n_10),
.B2(n_11),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_319),
.B(n_320),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_302),
.B(n_10),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_322),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_310),
.A2(n_11),
.B(n_12),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_304),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_324),
.B(n_329),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_304),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_309),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_330),
.A2(n_320),
.B(n_314),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_333),
.Y(n_334)
);

AOI322xp5_ASAP7_75t_L g333 ( 
.A1(n_327),
.A2(n_323),
.A3(n_319),
.B1(n_305),
.B2(n_306),
.C1(n_15),
.C2(n_16),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_324),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_326),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_325),
.B(n_332),
.Y(n_338)
);

A2O1A1Ixp33_ASAP7_75t_SL g339 ( 
.A1(n_338),
.A2(n_328),
.B(n_12),
.C(n_14),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_12),
.Y(n_340)
);


endmodule