module fake_jpeg_16391_n_231 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_231);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_36),
.Y(n_54)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_23),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_SL g43 ( 
.A1(n_38),
.A2(n_16),
.B(n_28),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_55),
.B(n_58),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_38),
.A2(n_24),
.B1(n_16),
.B2(n_21),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_44),
.A2(n_49),
.B1(n_50),
.B2(n_56),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_24),
.B1(n_16),
.B2(n_23),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_24),
.B1(n_29),
.B2(n_15),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_34),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_15),
.B1(n_29),
.B2(n_18),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_61),
.B1(n_42),
.B2(n_35),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_33),
.A2(n_30),
.B1(n_21),
.B2(n_26),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_32),
.A2(n_30),
.B1(n_26),
.B2(n_22),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_33),
.A2(n_30),
.B1(n_19),
.B2(n_18),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_32),
.A2(n_19),
.B1(n_31),
.B2(n_28),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_0),
.B(n_2),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_31),
.B1(n_28),
.B2(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_84),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_52),
.B(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_65),
.B(n_69),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_36),
.B1(n_42),
.B2(n_35),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_70),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_68),
.A2(n_76),
.B1(n_82),
.B2(n_46),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_17),
.Y(n_69)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

OR2x2_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_17),
.Y(n_72)
);

NOR2xp67_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_31),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_54),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_62),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_74),
.A2(n_77),
.B(n_50),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_47),
.A2(n_11),
.B1(n_3),
.B2(n_4),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_34),
.B1(n_41),
.B2(n_37),
.Y(n_76)
);

AND2x4_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_34),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_80),
.Y(n_100)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_47),
.A2(n_11),
.B1(n_3),
.B2(n_4),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_41),
.Y(n_84)
);

CKINVDCx11_ASAP7_75t_R g85 ( 
.A(n_80),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_85),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_63),
.A2(n_49),
.B1(n_56),
.B2(n_55),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_86),
.A2(n_88),
.B1(n_94),
.B2(n_98),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_63),
.A2(n_58),
.B1(n_48),
.B2(n_59),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_89),
.B(n_73),
.Y(n_112)
);

NAND2xp33_ASAP7_75t_SL g90 ( 
.A(n_77),
.B(n_72),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_84),
.Y(n_119)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_95),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_92),
.A2(n_0),
.B(n_39),
.Y(n_129)
);

NOR3xp33_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_74),
.C(n_76),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_77),
.A2(n_48),
.B1(n_59),
.B2(n_61),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_77),
.A2(n_59),
.B1(n_46),
.B2(n_47),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_53),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_78),
.Y(n_113)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_12),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_104),
.B(n_78),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_83),
.B1(n_71),
.B2(n_68),
.Y(n_124)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_107),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_110),
.Y(n_132)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_112),
.A2(n_119),
.B(n_129),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_123),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_116),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_115),
.A2(n_124),
.B(n_97),
.Y(n_136)
);

INVxp33_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_118),
.Y(n_135)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_120),
.Y(n_139)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_69),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_98),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_125),
.B(n_100),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_64),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_127),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_79),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_87),
.B(n_45),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_94),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_93),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_136),
.B(n_137),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_90),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_110),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_145),
.Y(n_157)
);

AOI322xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_104),
.A3(n_92),
.B1(n_103),
.B2(n_88),
.C1(n_86),
.C2(n_102),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_142),
.B(n_143),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_103),
.B(n_99),
.Y(n_143)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_117),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_104),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_129),
.C(n_128),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_100),
.B1(n_81),
.B2(n_96),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_147),
.A2(n_148),
.B1(n_108),
.B2(n_109),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_81),
.Y(n_150)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_150),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_132),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_151),
.B(n_166),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_149),
.Y(n_181)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_159),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_126),
.C(n_113),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_162),
.C(n_143),
.Y(n_172)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_118),
.Y(n_160)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_137),
.A2(n_114),
.B1(n_124),
.B2(n_112),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_161),
.A2(n_163),
.B1(n_133),
.B2(n_138),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_123),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_120),
.Y(n_164)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_164),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_111),
.Y(n_165)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_132),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_131),
.Y(n_167)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_131),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_151),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_181),
.C(n_169),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_137),
.B1(n_130),
.B2(n_144),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_174),
.A2(n_177),
.B1(n_155),
.B2(n_163),
.Y(n_194)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_176),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_161),
.A2(n_136),
.B1(n_133),
.B2(n_138),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_158),
.B(n_140),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_162),
.Y(n_187)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_183),
.B(n_166),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_179),
.A2(n_153),
.B1(n_130),
.B2(n_154),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_193),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_186),
.B(n_192),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_194),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_152),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_189),
.C(n_196),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_195),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_175),
.B(n_165),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

AOI322xp5_ASAP7_75t_SL g195 ( 
.A1(n_177),
.A2(n_169),
.A3(n_155),
.B1(n_167),
.B2(n_168),
.C1(n_156),
.C2(n_135),
.Y(n_195)
);

OAI31xp33_ASAP7_75t_L g196 ( 
.A1(n_174),
.A2(n_150),
.A3(n_145),
.B(n_141),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_182),
.C(n_178),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_200),
.C(n_204),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_181),
.C(n_171),
.Y(n_200)
);

FAx1_ASAP7_75t_SL g202 ( 
.A(n_187),
.B(n_184),
.CI(n_135),
.CON(n_202),
.SN(n_202)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_202),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_180),
.C(n_170),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_111),
.C(n_159),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_206),
.B(n_193),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_203),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_201),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_196),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_208),
.B(n_213),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_209),
.C(n_207),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_91),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_203),
.Y(n_218)
);

A2O1A1O1Ixp25_ASAP7_75t_L g213 ( 
.A1(n_202),
.A2(n_91),
.B(n_25),
.C(n_6),
.D(n_7),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_216),
.C(n_218),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_219),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_205),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_210),
.A2(n_122),
.B1(n_70),
.B2(n_7),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_215),
.A2(n_70),
.B1(n_5),
.B2(n_7),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_221),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_217),
.A2(n_101),
.B(n_8),
.Y(n_221)
);

AOI322xp5_ASAP7_75t_L g225 ( 
.A1(n_223),
.A2(n_101),
.A3(n_41),
.B1(n_39),
.B2(n_37),
.C1(n_25),
.C2(n_13),
.Y(n_225)
);

AOI332xp33_ASAP7_75t_L g227 ( 
.A1(n_225),
.A2(n_101),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.B3(n_8),
.C1(n_14),
.C2(n_13),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_3),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_25),
.C(n_13),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_227),
.A2(n_228),
.B(n_224),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_9),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_9),
.Y(n_231)
);


endmodule