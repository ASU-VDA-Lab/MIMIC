module fake_jpeg_11751_n_63 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_63);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_63;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_28),
.B(n_31),
.Y(n_35)
);

INVxp33_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_30),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_26),
.Y(n_31)
);

FAx1_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_26),
.CI(n_24),
.CON(n_32),
.SN(n_32)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_33),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_0),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_32),
.A2(n_25),
.B1(n_21),
.B2(n_10),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_40),
.B1(n_2),
.B2(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_39),
.Y(n_44)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_41),
.B(n_1),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_45),
.C(n_46),
.Y(n_51)
);

INVxp67_ASAP7_75t_SL g54 ( 
.A(n_43),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_2),
.B(n_4),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_34),
.B(n_36),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_39),
.B1(n_13),
.B2(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

AND2x6_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_55),
.Y(n_58)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_48),
.C(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_57),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_11),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_54),
.B(n_58),
.Y(n_60)
);

AOI322xp5_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_57),
.A3(n_50),
.B1(n_54),
.B2(n_17),
.C1(n_19),
.C2(n_15),
.Y(n_61)
);

NAND3xp33_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_18),
.C(n_5),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_4),
.B(n_5),
.Y(n_63)
);


endmodule