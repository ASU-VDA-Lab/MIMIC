module fake_netlist_6_4068_n_1909 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1909);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1909;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1892;
wire n_1459;
wire n_1614;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_171;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g171 ( 
.A(n_2),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_34),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_142),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_52),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_1),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_61),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_14),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_36),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_95),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_122),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_27),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_42),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_78),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_70),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_22),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_33),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_35),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

BUFx10_ASAP7_75t_L g190 ( 
.A(n_133),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_147),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_137),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_116),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_107),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_146),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_62),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_43),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_125),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_85),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_111),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_18),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_77),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_84),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_1),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_13),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_121),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_93),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_63),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_91),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_156),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_97),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_117),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_72),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_94),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_73),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g216 ( 
.A(n_168),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_154),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_150),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_31),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_51),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_112),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_101),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_53),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_68),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_141),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_109),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_148),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_29),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_114),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_162),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_129),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_48),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_139),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_165),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_27),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_8),
.Y(n_236)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_4),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_115),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_6),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_12),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_39),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_103),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_0),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_38),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_149),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_124),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_6),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_12),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_9),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_71),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_30),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_25),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_96),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_82),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_24),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_166),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_161),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_118),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_44),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_140),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_62),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_152),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_87),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_29),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_11),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_49),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_53),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_61),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_60),
.Y(n_269)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_92),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_104),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_39),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_79),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_83),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_48),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_151),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_110),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_20),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_67),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_52),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_36),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_2),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_24),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_153),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_25),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_66),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_14),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_13),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_45),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_132),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_65),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_42),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_43),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_134),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_32),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_76),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_126),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_163),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_20),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_37),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_145),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_74),
.Y(n_302)
);

BUFx10_ASAP7_75t_L g303 ( 
.A(n_54),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_100),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_56),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_106),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_80),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_35),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_38),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_41),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_86),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_130),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_3),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_31),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_45),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_90),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_17),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_54),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_123),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_9),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_60),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_75),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_56),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_169),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_41),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_105),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_158),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_30),
.Y(n_328)
);

BUFx8_ASAP7_75t_SL g329 ( 
.A(n_69),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_23),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_11),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_49),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_50),
.Y(n_333)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_157),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_120),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_159),
.Y(n_336)
);

BUFx2_ASAP7_75t_SL g337 ( 
.A(n_51),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_102),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_46),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_34),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_237),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_200),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_329),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_246),
.B(n_0),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_207),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_237),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_208),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_237),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_209),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_247),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_237),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_290),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_237),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_237),
.Y(n_354)
);

NOR2xp67_ASAP7_75t_L g355 ( 
.A(n_247),
.B(n_3),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_247),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_210),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_237),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_237),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_212),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_297),
.Y(n_361)
);

INVxp33_ASAP7_75t_SL g362 ( 
.A(n_174),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_223),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_173),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_325),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_334),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_213),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_325),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_325),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_246),
.B(n_4),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_193),
.B(n_5),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_325),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_221),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_175),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_303),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_303),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_303),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_222),
.Y(n_378)
);

NOR2xp67_ASAP7_75t_L g379 ( 
.A(n_334),
.B(n_5),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_224),
.Y(n_380)
);

INVxp67_ASAP7_75t_SL g381 ( 
.A(n_334),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_225),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_325),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_171),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_229),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_176),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_171),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_260),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_230),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_231),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_299),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_233),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_190),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_234),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_238),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_253),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_178),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_243),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_243),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_257),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_258),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_263),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_337),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_333),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_271),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_333),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_178),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_172),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_277),
.Y(n_409)
);

NOR2xp67_ASAP7_75t_L g410 ( 
.A(n_241),
.B(n_7),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_186),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_279),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_196),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_284),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_205),
.Y(n_415)
);

INVxp33_ASAP7_75t_L g416 ( 
.A(n_228),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_300),
.B(n_7),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_270),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_294),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_236),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_214),
.B(n_8),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_240),
.Y(n_422)
);

INVxp67_ASAP7_75t_SL g423 ( 
.A(n_184),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_365),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_350),
.B(n_214),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_346),
.Y(n_426)
);

OA21x2_ASAP7_75t_L g427 ( 
.A1(n_341),
.A2(n_249),
.B(n_248),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_365),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_346),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_368),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_368),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_369),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_346),
.Y(n_433)
);

BUFx8_ASAP7_75t_L g434 ( 
.A(n_407),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_351),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_369),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_351),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_379),
.B(n_250),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_351),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_341),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_379),
.B(n_388),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_372),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_410),
.B(n_190),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_366),
.B(n_180),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_356),
.B(n_423),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_418),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_381),
.B(n_180),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_378),
.Y(n_448)
);

OAI21x1_ASAP7_75t_L g449 ( 
.A1(n_388),
.A2(n_276),
.B(n_250),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_372),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_386),
.Y(n_451)
);

AND2x6_ASAP7_75t_L g452 ( 
.A(n_388),
.B(n_276),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_348),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_383),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_383),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_348),
.Y(n_456)
);

NAND3xp33_ASAP7_75t_L g457 ( 
.A(n_344),
.B(n_255),
.C(n_241),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_370),
.B(n_181),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_388),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_353),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_386),
.B(n_353),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_418),
.Y(n_462)
);

INVx5_ASAP7_75t_L g463 ( 
.A(n_418),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_354),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_354),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_358),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_358),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_359),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_359),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_408),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_384),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_384),
.Y(n_472)
);

AND2x6_ASAP7_75t_L g473 ( 
.A(n_421),
.B(n_260),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_386),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_355),
.B(n_181),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_375),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_355),
.B(n_260),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_407),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_408),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_387),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_387),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_398),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_413),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_397),
.B(n_185),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_398),
.Y(n_485)
);

INVx6_ASAP7_75t_L g486 ( 
.A(n_393),
.Y(n_486)
);

AND2x6_ASAP7_75t_L g487 ( 
.A(n_371),
.B(n_260),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_399),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_399),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_404),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_404),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_410),
.B(n_260),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_406),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_406),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_413),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_393),
.B(n_190),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_415),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_415),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_420),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_446),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_446),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_446),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_468),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_451),
.B(n_345),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_451),
.B(n_347),
.Y(n_505)
);

CKINVDCx6p67_ASAP7_75t_R g506 ( 
.A(n_496),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_425),
.B(n_374),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_429),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_444),
.B(n_349),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_484),
.B(n_357),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_484),
.B(n_360),
.Y(n_511)
);

NAND2xp33_ASAP7_75t_SL g512 ( 
.A(n_496),
.B(n_364),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_425),
.B(n_445),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_468),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_451),
.B(n_367),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_429),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_425),
.B(n_373),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_476),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_476),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_444),
.Y(n_520)
);

AND2x6_ASAP7_75t_L g521 ( 
.A(n_477),
.B(n_273),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_447),
.B(n_380),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_447),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_445),
.B(n_374),
.Y(n_524)
);

BUFx10_ASAP7_75t_L g525 ( 
.A(n_486),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_465),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_475),
.B(n_385),
.Y(n_527)
);

NAND2xp33_ASAP7_75t_L g528 ( 
.A(n_487),
.B(n_389),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_465),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_429),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_475),
.B(n_394),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_429),
.Y(n_532)
);

INVx1_ASAP7_75t_SL g533 ( 
.A(n_476),
.Y(n_533)
);

AOI21x1_ASAP7_75t_L g534 ( 
.A1(n_461),
.A2(n_191),
.B(n_189),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_446),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_433),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_433),
.Y(n_537)
);

INVx4_ASAP7_75t_SL g538 ( 
.A(n_473),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_465),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_465),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_446),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_465),
.Y(n_542)
);

INVx2_ASAP7_75t_SL g543 ( 
.A(n_438),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_440),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_446),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_445),
.B(n_395),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_446),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_440),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_492),
.B(n_396),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_478),
.B(n_403),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_433),
.Y(n_551)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_458),
.B(n_391),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_474),
.Y(n_553)
);

OR2x6_ASAP7_75t_L g554 ( 
.A(n_486),
.B(n_255),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_443),
.B(n_401),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_478),
.B(n_420),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_433),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_439),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_439),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_446),
.Y(n_560)
);

INVx1_ASAP7_75t_SL g561 ( 
.A(n_448),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_439),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_458),
.B(n_405),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_439),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_474),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_443),
.B(n_414),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_457),
.B(n_362),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_440),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_440),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_457),
.B(n_382),
.Y(n_570)
);

OR2x6_ASAP7_75t_L g571 ( 
.A(n_486),
.B(n_192),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_453),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_492),
.B(n_202),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_478),
.B(n_390),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_478),
.B(n_195),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g576 ( 
.A(n_461),
.B(n_363),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_435),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_426),
.Y(n_578)
);

BUFx10_ASAP7_75t_L g579 ( 
.A(n_486),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_435),
.Y(n_580)
);

OR2x2_ASAP7_75t_L g581 ( 
.A(n_427),
.B(n_376),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_453),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_471),
.B(n_422),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_435),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_435),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_435),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_486),
.B(n_392),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_453),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_453),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_486),
.B(n_400),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_456),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_456),
.Y(n_592)
);

OAI22xp33_ASAP7_75t_SL g593 ( 
.A1(n_438),
.A2(n_377),
.B1(n_411),
.B2(n_275),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_492),
.B(n_274),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_456),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_486),
.B(n_402),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_426),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_492),
.B(n_296),
.Y(n_598)
);

OR2x6_ASAP7_75t_L g599 ( 
.A(n_438),
.B(n_198),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_438),
.A2(n_487),
.B1(n_473),
.B2(n_427),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_456),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_438),
.A2(n_252),
.B1(n_269),
.B2(n_330),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_460),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_460),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_426),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_438),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_495),
.B(n_409),
.Y(n_607)
);

INVxp67_ASAP7_75t_SL g608 ( 
.A(n_474),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_495),
.B(n_412),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_463),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_460),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_426),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_492),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_492),
.B(n_419),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_460),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_467),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_467),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_487),
.A2(n_280),
.B1(n_305),
.B2(n_295),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_434),
.B(n_343),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_467),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_467),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_434),
.B(n_216),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_495),
.B(n_416),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_469),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_426),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_469),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_469),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_477),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_474),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_474),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_469),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_424),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_427),
.Y(n_633)
);

INVx6_ASAP7_75t_L g634 ( 
.A(n_474),
.Y(n_634)
);

OR2x6_ASAP7_75t_L g635 ( 
.A(n_427),
.B(n_211),
.Y(n_635)
);

INVx1_ASAP7_75t_SL g636 ( 
.A(n_448),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_471),
.B(n_422),
.Y(n_637)
);

INVx1_ASAP7_75t_SL g638 ( 
.A(n_427),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_434),
.B(n_216),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_495),
.B(n_342),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_424),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_424),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_427),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_477),
.B(n_215),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_441),
.B(n_298),
.Y(n_645)
);

AND3x2_ASAP7_75t_L g646 ( 
.A(n_477),
.B(n_218),
.C(n_217),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_495),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_487),
.A2(n_293),
.B1(n_320),
.B2(n_287),
.Y(n_648)
);

OR2x2_ASAP7_75t_L g649 ( 
.A(n_470),
.B(n_264),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_428),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_474),
.B(n_352),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_436),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_632),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_520),
.B(n_487),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_507),
.B(n_524),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_543),
.B(n_474),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_543),
.B(n_441),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_647),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_632),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_520),
.A2(n_487),
.B1(n_361),
.B2(n_473),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_641),
.Y(n_661)
);

BUFx6f_ASAP7_75t_SL g662 ( 
.A(n_523),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_507),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_606),
.A2(n_628),
.B(n_613),
.Y(n_664)
);

O2A1O1Ixp33_ASAP7_75t_L g665 ( 
.A1(n_581),
.A2(n_498),
.B(n_497),
.C(n_470),
.Y(n_665)
);

INVx8_ASAP7_75t_L g666 ( 
.A(n_554),
.Y(n_666)
);

INVx6_ASAP7_75t_L g667 ( 
.A(n_644),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_523),
.B(n_487),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_552),
.B(n_292),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_556),
.Y(n_670)
);

NOR2xp67_ASAP7_75t_L g671 ( 
.A(n_552),
.B(n_477),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_563),
.B(n_487),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_580),
.Y(n_673)
);

AND2x6_ASAP7_75t_SL g674 ( 
.A(n_570),
.B(n_281),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_509),
.B(n_487),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_546),
.B(n_185),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_524),
.Y(n_677)
);

INVxp67_ASAP7_75t_L g678 ( 
.A(n_518),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_522),
.B(n_487),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_641),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_513),
.B(n_479),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_642),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_513),
.B(n_487),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_623),
.B(n_441),
.Y(n_684)
);

BUFx5_ASAP7_75t_L g685 ( 
.A(n_633),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_633),
.A2(n_473),
.B1(n_477),
.B2(n_449),
.Y(n_686)
);

AND2x6_ASAP7_75t_SL g687 ( 
.A(n_574),
.B(n_417),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_613),
.B(n_441),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_518),
.B(n_417),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_517),
.B(n_441),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_628),
.B(n_434),
.Y(n_691)
);

OAI21xp5_ASAP7_75t_L g692 ( 
.A1(n_643),
.A2(n_449),
.B(n_473),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_583),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_642),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_503),
.B(n_464),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_533),
.B(n_576),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_503),
.B(n_464),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_583),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_514),
.B(n_464),
.Y(n_699)
);

NAND2xp33_ASAP7_75t_L g700 ( 
.A(n_638),
.B(n_473),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_581),
.B(n_194),
.Y(n_701)
);

NAND2x1p5_ASAP7_75t_L g702 ( 
.A(n_638),
.B(n_643),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_514),
.B(n_464),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_576),
.B(n_194),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_580),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_573),
.B(n_594),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_550),
.B(n_464),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_600),
.B(n_607),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_637),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_637),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_609),
.B(n_644),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_533),
.B(n_479),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_650),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_550),
.B(n_464),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_652),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_650),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_644),
.B(n_434),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_549),
.B(n_464),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_652),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_556),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_526),
.B(n_464),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_526),
.B(n_529),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_539),
.B(n_466),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_539),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_575),
.B(n_483),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_540),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_540),
.B(n_542),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_589),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_542),
.B(n_466),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_589),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_591),
.Y(n_731)
);

INVx4_ASAP7_75t_L g732 ( 
.A(n_502),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_519),
.B(n_199),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_504),
.B(n_466),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_505),
.B(n_515),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_510),
.B(n_199),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_644),
.B(n_466),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_575),
.Y(n_738)
);

NAND2xp33_ASAP7_75t_L g739 ( 
.A(n_521),
.B(n_473),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_575),
.B(n_466),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_649),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_591),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_595),
.Y(n_743)
);

OAI221xp5_ASAP7_75t_L g744 ( 
.A1(n_602),
.A2(n_483),
.B1(n_498),
.B2(n_497),
.C(n_327),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_SL g745 ( 
.A(n_506),
.B(n_340),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_525),
.B(n_434),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_511),
.B(n_203),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_649),
.B(n_497),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_575),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_645),
.B(n_466),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_651),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_595),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_527),
.B(n_203),
.Y(n_753)
);

NOR2x1p5_ASAP7_75t_L g754 ( 
.A(n_506),
.B(n_174),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_640),
.B(n_498),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_598),
.B(n_466),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_567),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_500),
.B(n_466),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_577),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_601),
.Y(n_760)
);

NAND2xp33_ASAP7_75t_L g761 ( 
.A(n_521),
.B(n_473),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_500),
.B(n_473),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_531),
.B(n_206),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_577),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_555),
.B(n_206),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_525),
.B(n_273),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_646),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_566),
.B(n_256),
.Y(n_768)
);

NAND2x1_ASAP7_75t_L g769 ( 
.A(n_634),
.B(n_473),
.Y(n_769)
);

NAND3xp33_ASAP7_75t_L g770 ( 
.A(n_614),
.B(n_220),
.C(n_219),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_553),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_500),
.B(n_473),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_553),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_553),
.Y(n_774)
);

BUFx5_ASAP7_75t_L g775 ( 
.A(n_525),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_593),
.B(n_256),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_500),
.B(n_426),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_587),
.A2(n_322),
.B1(n_326),
.B2(n_335),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_501),
.B(n_426),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_635),
.A2(n_449),
.B1(n_273),
.B2(n_270),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_635),
.Y(n_781)
);

NOR3xp33_ASAP7_75t_L g782 ( 
.A(n_512),
.B(n_235),
.C(n_232),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_584),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_501),
.B(n_426),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_593),
.B(n_301),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_601),
.Y(n_786)
);

INVx2_ASAP7_75t_SL g787 ( 
.A(n_635),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_501),
.B(n_437),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_590),
.A2(n_596),
.B1(n_528),
.B2(n_599),
.Y(n_789)
);

OAI22xp5_ASAP7_75t_L g790 ( 
.A1(n_554),
.A2(n_226),
.B1(n_227),
.B2(n_242),
.Y(n_790)
);

OR2x2_ASAP7_75t_L g791 ( 
.A(n_561),
.B(n_177),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_525),
.B(n_273),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_501),
.B(n_535),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_584),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_599),
.A2(n_336),
.B1(n_338),
.B2(n_306),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_615),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_535),
.B(n_437),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_579),
.B(n_273),
.Y(n_798)
);

NOR2xp67_ASAP7_75t_L g799 ( 
.A(n_622),
.B(n_480),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_535),
.B(n_437),
.Y(n_800)
);

BUFx6f_ASAP7_75t_SL g801 ( 
.A(n_635),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_635),
.A2(n_270),
.B1(n_307),
.B2(n_254),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_535),
.B(n_437),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_599),
.A2(n_306),
.B1(n_319),
.B2(n_312),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_580),
.Y(n_805)
);

AOI221xp5_ASAP7_75t_L g806 ( 
.A1(n_639),
.A2(n_177),
.B1(n_339),
.B2(n_179),
.C(n_182),
.Y(n_806)
);

O2A1O1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_544),
.A2(n_604),
.B(n_588),
.C(n_592),
.Y(n_807)
);

INVxp67_ASAP7_75t_L g808 ( 
.A(n_561),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_547),
.B(n_597),
.Y(n_809)
);

NAND2xp33_ASAP7_75t_L g810 ( 
.A(n_521),
.B(n_270),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_585),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_547),
.B(n_437),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_547),
.B(n_437),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_547),
.B(n_437),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_619),
.B(n_301),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_599),
.B(n_471),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_579),
.B(n_538),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_585),
.Y(n_818)
);

BUFx8_ASAP7_75t_L g819 ( 
.A(n_636),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_615),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_586),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_597),
.B(n_437),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_586),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_755),
.B(n_597),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_670),
.Y(n_825)
);

INVx5_ASAP7_75t_L g826 ( 
.A(n_666),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_706),
.B(n_597),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_775),
.B(n_579),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_670),
.Y(n_829)
);

O2A1O1Ixp33_ASAP7_75t_L g830 ( 
.A1(n_708),
.A2(n_599),
.B(n_554),
.C(n_617),
.Y(n_830)
);

OAI21xp5_ASAP7_75t_L g831 ( 
.A1(n_683),
.A2(n_608),
.B(n_548),
.Y(n_831)
);

OAI21xp33_ASAP7_75t_L g832 ( 
.A1(n_669),
.A2(n_182),
.B(n_179),
.Y(n_832)
);

INVx4_ASAP7_75t_L g833 ( 
.A(n_667),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_775),
.B(n_579),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_693),
.B(n_554),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_692),
.A2(n_548),
.B(n_544),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_671),
.B(n_605),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_655),
.B(n_636),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_771),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_696),
.B(n_554),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_653),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_709),
.B(n_605),
.Y(n_842)
);

BUFx12f_ASAP7_75t_L g843 ( 
.A(n_819),
.Y(n_843)
);

O2A1O1Ixp5_ASAP7_75t_L g844 ( 
.A1(n_708),
.A2(n_534),
.B(n_605),
.C(n_631),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_775),
.B(n_538),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_657),
.A2(n_629),
.B(n_565),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_657),
.A2(n_629),
.B(n_565),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_709),
.B(n_605),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_688),
.A2(n_629),
.B(n_565),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_718),
.A2(n_630),
.B(n_541),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_653),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_684),
.A2(n_630),
.B(n_541),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_676),
.A2(n_648),
.B(n_618),
.C(n_316),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_756),
.A2(n_630),
.B(n_541),
.Y(n_854)
);

AOI22x1_ASAP7_75t_SL g855 ( 
.A1(n_658),
.A2(n_314),
.B1(n_204),
.B2(n_201),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_773),
.A2(n_541),
.B(n_502),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_712),
.B(n_571),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_771),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_735),
.B(n_568),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_659),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_681),
.B(n_568),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_676),
.B(n_569),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_690),
.B(n_685),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_663),
.B(n_538),
.Y(n_864)
);

OAI21xp5_ASAP7_75t_L g865 ( 
.A1(n_700),
.A2(n_672),
.B(n_675),
.Y(n_865)
);

AOI211xp5_ASAP7_75t_L g866 ( 
.A1(n_669),
.A2(n_314),
.B(n_204),
.C(n_339),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_819),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_789),
.A2(n_571),
.B1(n_634),
.B2(n_291),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_711),
.A2(n_677),
.B1(n_660),
.B2(n_781),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_659),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_698),
.B(n_571),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_724),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_741),
.B(n_571),
.Y(n_873)
);

NOR3xp33_ASAP7_75t_L g874 ( 
.A(n_806),
.B(n_304),
.C(n_302),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_685),
.B(n_569),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_685),
.B(n_572),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_773),
.A2(n_541),
.B(n_502),
.Y(n_877)
);

OAI22x1_ASAP7_75t_L g878 ( 
.A1(n_678),
.A2(n_313),
.B1(n_187),
.B2(n_188),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_741),
.B(n_571),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_704),
.B(n_572),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_685),
.B(n_582),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_L g882 ( 
.A1(n_679),
.A2(n_588),
.B(n_582),
.Y(n_882)
);

NOR2xp67_ASAP7_75t_L g883 ( 
.A(n_808),
.B(n_534),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_661),
.Y(n_884)
);

AOI21x1_ASAP7_75t_L g885 ( 
.A1(n_656),
.A2(n_603),
.B(n_592),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_775),
.B(n_538),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_685),
.B(n_603),
.Y(n_887)
);

CKINVDCx11_ASAP7_75t_R g888 ( 
.A(n_674),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_748),
.B(n_499),
.Y(n_889)
);

A2O1A1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_815),
.A2(n_245),
.B(n_324),
.C(n_286),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_774),
.A2(n_545),
.B(n_502),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_702),
.Y(n_892)
);

AO21x1_ASAP7_75t_L g893 ( 
.A1(n_711),
.A2(n_262),
.B(n_604),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_685),
.B(n_611),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_774),
.A2(n_545),
.B(n_502),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_750),
.A2(n_560),
.B(n_545),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_734),
.A2(n_664),
.B(n_707),
.Y(n_897)
);

AO21x2_ASAP7_75t_L g898 ( 
.A1(n_691),
.A2(n_616),
.B(n_611),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_726),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_704),
.B(n_662),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_701),
.B(n_616),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_710),
.B(n_499),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_662),
.B(n_617),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_816),
.B(n_488),
.Y(n_904)
);

OAI22xp5_ASAP7_75t_L g905 ( 
.A1(n_702),
.A2(n_634),
.B1(n_612),
.B2(n_625),
.Y(n_905)
);

BUFx3_ASAP7_75t_L g906 ( 
.A(n_757),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_667),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_701),
.B(n_620),
.Y(n_908)
);

OAI21xp33_ASAP7_75t_L g909 ( 
.A1(n_733),
.A2(n_187),
.B(n_183),
.Y(n_909)
);

NOR2xp67_ASAP7_75t_L g910 ( 
.A(n_778),
.B(n_620),
.Y(n_910)
);

O2A1O1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_665),
.A2(n_626),
.B(n_631),
.C(n_627),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_715),
.B(n_626),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_719),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_738),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_720),
.B(n_621),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_714),
.A2(n_560),
.B(n_545),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_667),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_787),
.A2(n_521),
.B1(n_634),
.B2(n_627),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_656),
.A2(n_625),
.B(n_560),
.Y(n_919)
);

NOR2x1_ASAP7_75t_L g920 ( 
.A(n_751),
.B(n_436),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_661),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_775),
.B(n_545),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_749),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_680),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_680),
.Y(n_925)
);

A2O1A1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_815),
.A2(n_621),
.B(n_624),
.C(n_537),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_791),
.B(n_624),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_775),
.B(n_560),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_801),
.A2(n_521),
.B1(n_612),
.B2(n_578),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_654),
.A2(n_668),
.B(n_686),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_817),
.A2(n_625),
.B(n_612),
.Y(n_931)
);

OAI21x1_ASAP7_75t_L g932 ( 
.A1(n_762),
.A2(n_557),
.B(n_508),
.Y(n_932)
);

NOR2xp67_ASAP7_75t_L g933 ( 
.A(n_770),
.B(n_736),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_751),
.B(n_560),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_817),
.A2(n_625),
.B(n_612),
.Y(n_935)
);

BUFx8_ASAP7_75t_L g936 ( 
.A(n_689),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_816),
.B(n_578),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_771),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_733),
.B(n_499),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_737),
.A2(n_625),
.B(n_612),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_SL g941 ( 
.A(n_745),
.B(n_216),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_682),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_736),
.A2(n_551),
.B(n_516),
.C(n_564),
.Y(n_943)
);

A2O1A1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_747),
.A2(n_551),
.B(n_516),
.C(n_564),
.Y(n_944)
);

O2A1O1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_744),
.A2(n_557),
.B(n_562),
.C(n_559),
.Y(n_945)
);

O2A1O1Ixp5_ASAP7_75t_L g946 ( 
.A1(n_766),
.A2(n_537),
.B(n_530),
.C(n_562),
.Y(n_946)
);

INVxp67_ASAP7_75t_L g947 ( 
.A(n_725),
.Y(n_947)
);

OAI321xp33_ASAP7_75t_L g948 ( 
.A1(n_747),
.A2(n_488),
.A3(n_491),
.B1(n_494),
.B2(n_428),
.C(n_432),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_725),
.B(n_578),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_740),
.A2(n_578),
.B(n_610),
.Y(n_950)
);

NOR3xp33_ASAP7_75t_L g951 ( 
.A(n_753),
.B(n_302),
.C(n_304),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_682),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_753),
.B(n_578),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_763),
.B(n_532),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_694),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_767),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_763),
.B(n_499),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_694),
.Y(n_958)
);

INVx4_ASAP7_75t_L g959 ( 
.A(n_771),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_766),
.A2(n_610),
.B(n_462),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_792),
.A2(n_610),
.B(n_462),
.Y(n_961)
);

CKINVDCx10_ASAP7_75t_R g962 ( 
.A(n_687),
.Y(n_962)
);

BUFx12f_ASAP7_75t_L g963 ( 
.A(n_754),
.Y(n_963)
);

NAND3xp33_ASAP7_75t_L g964 ( 
.A(n_765),
.B(n_268),
.C(n_288),
.Y(n_964)
);

NOR2x2_ASAP7_75t_L g965 ( 
.A(n_776),
.B(n_183),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_713),
.B(n_532),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_776),
.B(n_239),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_713),
.B(n_536),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_666),
.Y(n_969)
);

OR2x6_ASAP7_75t_L g970 ( 
.A(n_666),
.B(n_488),
.Y(n_970)
);

A2O1A1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_765),
.A2(n_536),
.B(n_559),
.C(n_558),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_792),
.A2(n_610),
.B(n_462),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_716),
.B(n_521),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_798),
.A2(n_462),
.B(n_463),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_732),
.A2(n_462),
.B(n_463),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_769),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_716),
.B(n_521),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_732),
.A2(n_809),
.B(n_793),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_785),
.B(n_244),
.Y(n_979)
);

OAI21xp33_ASAP7_75t_L g980 ( 
.A1(n_768),
.A2(n_309),
.B(n_197),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_801),
.Y(n_981)
);

AOI33xp33_ASAP7_75t_L g982 ( 
.A1(n_802),
.A2(n_494),
.A3(n_491),
.B1(n_188),
.B2(n_318),
.B3(n_197),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_728),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_722),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_785),
.B(n_251),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_686),
.B(n_802),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_768),
.A2(n_482),
.B(n_480),
.C(n_490),
.Y(n_987)
);

NOR3xp33_ASAP7_75t_L g988 ( 
.A(n_782),
.B(n_790),
.C(n_804),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_727),
.Y(n_989)
);

BUFx12f_ASAP7_75t_L g990 ( 
.A(n_795),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_799),
.B(n_311),
.Y(n_991)
);

AOI22xp33_ASAP7_75t_L g992 ( 
.A1(n_780),
.A2(n_270),
.B1(n_201),
.B2(n_309),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_728),
.B(n_480),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_777),
.A2(n_463),
.B(n_459),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_759),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_695),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_780),
.A2(n_311),
.B1(n_319),
.B2(n_312),
.Y(n_997)
);

AND2x2_ASAP7_75t_SL g998 ( 
.A(n_739),
.B(n_428),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_779),
.A2(n_463),
.B(n_459),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_697),
.B(n_259),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_730),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_807),
.A2(n_459),
.B(n_430),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_699),
.A2(n_480),
.B(n_482),
.C(n_490),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_764),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_703),
.A2(n_480),
.B(n_482),
.C(n_490),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_784),
.A2(n_463),
.B(n_430),
.Y(n_1006)
);

AOI21x1_ASAP7_75t_L g1007 ( 
.A1(n_772),
.A2(n_455),
.B(n_430),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_788),
.A2(n_463),
.B(n_432),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_730),
.B(n_482),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_673),
.B(n_705),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_731),
.B(n_482),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_721),
.A2(n_432),
.B(n_442),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_805),
.B(n_270),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_986),
.A2(n_717),
.B1(n_691),
.B2(n_746),
.Y(n_1014)
);

AOI33xp33_ASAP7_75t_L g1015 ( 
.A1(n_866),
.A2(n_491),
.A3(n_494),
.B1(n_818),
.B2(n_811),
.B3(n_823),
.Y(n_1015)
);

BUFx2_ASAP7_75t_L g1016 ( 
.A(n_936),
.Y(n_1016)
);

A2O1A1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_967),
.A2(n_985),
.B(n_979),
.C(n_933),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_828),
.A2(n_746),
.B(n_717),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_986),
.A2(n_743),
.B1(n_796),
.B2(n_820),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_989),
.B(n_731),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_913),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_947),
.B(n_783),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_967),
.A2(n_794),
.B(n_821),
.C(n_729),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_983),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_838),
.B(n_723),
.Y(n_1025)
);

NOR3xp33_ASAP7_75t_L g1026 ( 
.A(n_979),
.B(n_272),
.C(n_265),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_936),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_989),
.B(n_742),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_985),
.A2(n_761),
.B1(n_810),
.B2(n_338),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_857),
.B(n_742),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_839),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_951),
.A2(n_796),
.B(n_820),
.C(n_743),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_828),
.A2(n_803),
.B(n_814),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_840),
.B(n_752),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_900),
.B(n_947),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_872),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_956),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_834),
.A2(n_813),
.B(n_812),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_992),
.A2(n_752),
.B1(n_760),
.B2(n_786),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_984),
.B(n_760),
.Y(n_1040)
);

OR2x6_ASAP7_75t_L g1041 ( 
.A(n_969),
.B(n_797),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_874),
.A2(n_786),
.B(n_758),
.C(n_822),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_839),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_899),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_927),
.B(n_800),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_951),
.A2(n_485),
.B(n_490),
.C(n_266),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_1001),
.Y(n_1047)
);

BUFx4_ASAP7_75t_SL g1048 ( 
.A(n_867),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_942),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_874),
.A2(n_455),
.B(n_454),
.C(n_450),
.Y(n_1050)
);

BUFx5_ASAP7_75t_L g1051 ( 
.A(n_998),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_840),
.B(n_900),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_927),
.B(n_261),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_906),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_890),
.A2(n_455),
.B(n_454),
.C(n_450),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_992),
.A2(n_308),
.B1(n_310),
.B2(n_313),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_880),
.B(n_485),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_902),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_969),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_843),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_841),
.Y(n_1061)
);

INVxp67_ASAP7_75t_L g1062 ( 
.A(n_878),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_988),
.A2(n_490),
.B1(n_485),
.B2(n_431),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_880),
.B(n_485),
.Y(n_1064)
);

NOR2xp67_ASAP7_75t_SL g1065 ( 
.A(n_826),
.B(n_308),
.Y(n_1065)
);

AOI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_988),
.A2(n_485),
.B1(n_431),
.B2(n_450),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_851),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_SL g1068 ( 
.A1(n_903),
.A2(n_454),
.B(n_442),
.C(n_431),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_860),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_834),
.A2(n_463),
.B(n_481),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_863),
.A2(n_481),
.B(n_472),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_941),
.B(n_267),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_859),
.A2(n_869),
.B1(n_908),
.B2(n_901),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_922),
.A2(n_481),
.B(n_472),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_932),
.A2(n_442),
.B(n_481),
.Y(n_1075)
);

AOI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_873),
.A2(n_879),
.B1(n_835),
.B2(n_964),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_889),
.B(n_939),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_914),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_996),
.B(n_957),
.Y(n_1079)
);

INVx4_ASAP7_75t_L g1080 ( 
.A(n_969),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_922),
.A2(n_472),
.B(n_489),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_969),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_996),
.B(n_472),
.Y(n_1083)
);

INVx3_ASAP7_75t_L g1084 ( 
.A(n_839),
.Y(n_1084)
);

INVxp67_ASAP7_75t_L g1085 ( 
.A(n_981),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_904),
.B(n_283),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_928),
.A2(n_493),
.B(n_489),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_833),
.B(n_285),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_833),
.B(n_289),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_826),
.B(n_108),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_861),
.A2(n_321),
.B1(n_310),
.B2(n_315),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_832),
.B(n_278),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_980),
.B(n_282),
.Y(n_1093)
);

O2A1O1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_909),
.A2(n_323),
.B(n_331),
.C(n_328),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_923),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_997),
.A2(n_332),
.B(n_317),
.C(n_318),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_825),
.B(n_315),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_928),
.A2(n_493),
.B(n_489),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1000),
.B(n_824),
.Y(n_1099)
);

NAND3xp33_ASAP7_75t_L g1100 ( 
.A(n_1000),
.B(n_321),
.C(n_317),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_835),
.B(n_270),
.Y(n_1101)
);

BUFx8_ASAP7_75t_L g1102 ( 
.A(n_963),
.Y(n_1102)
);

INVx2_ASAP7_75t_SL g1103 ( 
.A(n_981),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_870),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_884),
.Y(n_1105)
);

AOI21x1_ASAP7_75t_L g1106 ( 
.A1(n_934),
.A2(n_270),
.B(n_489),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_990),
.Y(n_1107)
);

O2A1O1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_853),
.A2(n_10),
.B(n_15),
.C(n_16),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_830),
.A2(n_493),
.B(n_489),
.C(n_16),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_921),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_904),
.Y(n_1111)
);

BUFx12f_ASAP7_75t_L g1112 ( 
.A(n_888),
.Y(n_1112)
);

OR2x2_ASAP7_75t_L g1113 ( 
.A(n_829),
.B(n_493),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_924),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_873),
.B(n_879),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_839),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_871),
.B(n_493),
.Y(n_1117)
);

NOR3xp33_ASAP7_75t_SL g1118 ( 
.A(n_903),
.B(n_10),
.C(n_15),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_862),
.B(n_493),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_965),
.Y(n_1120)
);

AOI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_871),
.A2(n_452),
.B1(n_493),
.B2(n_489),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_892),
.B(n_17),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_R g1123 ( 
.A(n_826),
.B(n_81),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_925),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_952),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_955),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_L g1127 ( 
.A1(n_892),
.A2(n_452),
.B1(n_493),
.B2(n_489),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_865),
.A2(n_452),
.B(n_489),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_991),
.A2(n_18),
.B(n_19),
.C(n_21),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_958),
.Y(n_1130)
);

INVx4_ASAP7_75t_L g1131 ( 
.A(n_826),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_827),
.B(n_19),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_970),
.B(n_907),
.Y(n_1133)
);

INVx4_ASAP7_75t_L g1134 ( 
.A(n_858),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_995),
.B(n_21),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_915),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_930),
.A2(n_844),
.B(n_836),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_858),
.Y(n_1138)
);

AOI211xp5_ASAP7_75t_SL g1139 ( 
.A1(n_948),
.A2(n_22),
.B(n_23),
.C(n_26),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_837),
.A2(n_452),
.B(n_89),
.Y(n_1140)
);

O2A1O1Ixp33_ASAP7_75t_SL g1141 ( 
.A1(n_987),
.A2(n_864),
.B(n_1003),
.C(n_1005),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_982),
.B(n_26),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_858),
.Y(n_1143)
);

O2A1O1Ixp5_ASAP7_75t_L g1144 ( 
.A1(n_893),
.A2(n_98),
.B(n_170),
.C(n_167),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_953),
.A2(n_452),
.B(n_88),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_910),
.A2(n_831),
.B(n_954),
.C(n_883),
.Y(n_1146)
);

INVx5_ASAP7_75t_L g1147 ( 
.A(n_858),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_938),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_934),
.A2(n_28),
.B(n_32),
.C(n_33),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_938),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1004),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_846),
.A2(n_28),
.B(n_37),
.C(n_40),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_897),
.A2(n_452),
.B(n_113),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_920),
.B(n_40),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_907),
.B(n_44),
.Y(n_1155)
);

OA21x2_ASAP7_75t_L g1156 ( 
.A1(n_882),
.A2(n_452),
.B(n_127),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_847),
.A2(n_46),
.B(n_47),
.C(n_50),
.Y(n_1157)
);

OAI221xp5_ASAP7_75t_L g1158 ( 
.A1(n_917),
.A2(n_47),
.B1(n_55),
.B2(n_57),
.C(n_58),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_917),
.B(n_55),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_938),
.Y(n_1160)
);

NOR2x1_ASAP7_75t_L g1161 ( 
.A(n_959),
.B(n_970),
.Y(n_1161)
);

INVx1_ASAP7_75t_SL g1162 ( 
.A(n_938),
.Y(n_1162)
);

A2O1A1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_849),
.A2(n_57),
.B(n_58),
.C(n_59),
.Y(n_1163)
);

AOI21x1_ASAP7_75t_L g1164 ( 
.A1(n_852),
.A2(n_452),
.B(n_64),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_875),
.A2(n_452),
.B(n_99),
.Y(n_1165)
);

NAND2xp33_ASAP7_75t_L g1166 ( 
.A(n_976),
.B(n_452),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_937),
.A2(n_452),
.B1(n_59),
.B2(n_128),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_912),
.B(n_119),
.Y(n_1168)
);

AOI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_937),
.A2(n_949),
.B1(n_998),
.B2(n_970),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_842),
.A2(n_131),
.B(n_136),
.C(n_138),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_848),
.A2(n_911),
.B(n_978),
.C(n_850),
.Y(n_1171)
);

BUFx4f_ASAP7_75t_L g1172 ( 
.A(n_976),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_876),
.B(n_894),
.Y(n_1173)
);

INVx5_ASAP7_75t_L g1174 ( 
.A(n_1116),
.Y(n_1174)
);

INVxp67_ASAP7_75t_SL g1175 ( 
.A(n_1172),
.Y(n_1175)
);

A2O1A1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1017),
.A2(n_868),
.B(n_918),
.C(n_854),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1052),
.B(n_1035),
.Y(n_1177)
);

NAND3xp33_ASAP7_75t_L g1178 ( 
.A(n_1026),
.B(n_855),
.C(n_926),
.Y(n_1178)
);

INVxp67_ASAP7_75t_L g1179 ( 
.A(n_1054),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1115),
.B(n_959),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1136),
.B(n_976),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1021),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1053),
.B(n_976),
.Y(n_1183)
);

CKINVDCx11_ASAP7_75t_R g1184 ( 
.A(n_1112),
.Y(n_1184)
);

AO31x2_ASAP7_75t_L g1185 ( 
.A1(n_1014),
.A2(n_971),
.A3(n_944),
.B(n_943),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1075),
.A2(n_1038),
.B(n_1033),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1036),
.Y(n_1187)
);

INVx5_ASAP7_75t_L g1188 ( 
.A(n_1116),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1076),
.A2(n_929),
.B1(n_881),
.B2(n_887),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1100),
.A2(n_1002),
.B(n_945),
.C(n_916),
.Y(n_1190)
);

HB1xp67_ASAP7_75t_L g1191 ( 
.A(n_1111),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_1037),
.Y(n_1192)
);

INVx1_ASAP7_75t_SL g1193 ( 
.A(n_1086),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1044),
.Y(n_1194)
);

OAI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1139),
.A2(n_977),
.B1(n_973),
.B2(n_968),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1106),
.A2(n_896),
.B(n_885),
.Y(n_1196)
);

BUFx2_ASAP7_75t_L g1197 ( 
.A(n_1085),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1078),
.Y(n_1198)
);

AO32x2_ASAP7_75t_L g1199 ( 
.A1(n_1014),
.A2(n_905),
.A3(n_898),
.B1(n_1007),
.B2(n_1012),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1079),
.B(n_966),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_SL g1201 ( 
.A(n_1107),
.B(n_962),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1058),
.B(n_1077),
.Y(n_1202)
);

NAND3xp33_ASAP7_75t_L g1203 ( 
.A(n_1093),
.B(n_1013),
.C(n_940),
.Y(n_1203)
);

AOI221x1_ASAP7_75t_L g1204 ( 
.A1(n_1109),
.A2(n_919),
.B1(n_931),
.B2(n_935),
.C(n_877),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1025),
.B(n_898),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_1100),
.B(n_1010),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1092),
.B(n_1010),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1099),
.B(n_1011),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1071),
.A2(n_895),
.B(n_891),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_1059),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1019),
.A2(n_856),
.B(n_946),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1146),
.A2(n_1073),
.B(n_1171),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1073),
.A2(n_845),
.B(n_886),
.Y(n_1213)
);

O2A1O1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1096),
.A2(n_1013),
.B(n_1009),
.C(n_993),
.Y(n_1214)
);

AO31x2_ASAP7_75t_L g1215 ( 
.A1(n_1023),
.A2(n_1008),
.A3(n_1006),
.B(n_999),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1173),
.A2(n_845),
.B(n_886),
.Y(n_1216)
);

AOI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1122),
.A2(n_994),
.B1(n_950),
.B2(n_974),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1020),
.B(n_960),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_1059),
.Y(n_1219)
);

CKINVDCx11_ASAP7_75t_R g1220 ( 
.A(n_1016),
.Y(n_1220)
);

BUFx2_ASAP7_75t_L g1221 ( 
.A(n_1103),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_1102),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1172),
.A2(n_961),
.B(n_972),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1046),
.A2(n_975),
.A3(n_155),
.B(n_160),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1028),
.B(n_143),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1019),
.A2(n_164),
.B(n_1164),
.Y(n_1226)
);

AO31x2_ASAP7_75t_L g1227 ( 
.A1(n_1032),
.A2(n_1039),
.A3(n_1153),
.B(n_1152),
.Y(n_1227)
);

INVx1_ASAP7_75t_SL g1228 ( 
.A(n_1048),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1137),
.A2(n_1045),
.B(n_1119),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_SL g1230 ( 
.A1(n_1108),
.A2(n_1149),
.B(n_1169),
.Y(n_1230)
);

O2A1O1Ixp33_ASAP7_75t_SL g1231 ( 
.A1(n_1139),
.A2(n_1157),
.B(n_1170),
.C(n_1163),
.Y(n_1231)
);

AO31x2_ASAP7_75t_L g1232 ( 
.A1(n_1039),
.A2(n_1064),
.A3(n_1057),
.B(n_1132),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_SL g1233 ( 
.A1(n_1142),
.A2(n_1168),
.B(n_1068),
.C(n_1101),
.Y(n_1233)
);

AO31x2_ASAP7_75t_L g1234 ( 
.A1(n_1081),
.A2(n_1074),
.A3(n_1098),
.B(n_1087),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1095),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_1059),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1022),
.B(n_1040),
.Y(n_1237)
);

HB1xp67_ASAP7_75t_L g1238 ( 
.A(n_1022),
.Y(n_1238)
);

NAND3xp33_ASAP7_75t_L g1239 ( 
.A(n_1118),
.B(n_1094),
.C(n_1072),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1070),
.A2(n_1128),
.B(n_1042),
.Y(n_1240)
);

INVx8_ASAP7_75t_L g1241 ( 
.A(n_1147),
.Y(n_1241)
);

OR2x2_ASAP7_75t_L g1242 ( 
.A(n_1151),
.B(n_1091),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1137),
.A2(n_1015),
.B(n_1029),
.C(n_1129),
.Y(n_1243)
);

NAND3xp33_ASAP7_75t_L g1244 ( 
.A(n_1062),
.B(n_1056),
.C(n_1097),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1049),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1133),
.B(n_1051),
.Y(n_1246)
);

OAI22x1_ASAP7_75t_L g1247 ( 
.A1(n_1120),
.A2(n_1135),
.B1(n_1154),
.B2(n_1027),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_1131),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1030),
.A2(n_1158),
.B1(n_1056),
.B2(n_1155),
.Y(n_1249)
);

BUFx6f_ASAP7_75t_L g1250 ( 
.A(n_1082),
.Y(n_1250)
);

AOI21xp33_ASAP7_75t_L g1251 ( 
.A1(n_1091),
.A2(n_1159),
.B(n_1088),
.Y(n_1251)
);

NOR2x1_ASAP7_75t_SL g1252 ( 
.A(n_1147),
.B(n_1131),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1141),
.A2(n_1034),
.B(n_1128),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1105),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1083),
.A2(n_1161),
.B(n_1145),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1133),
.B(n_1024),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1156),
.A2(n_1117),
.B(n_1147),
.Y(n_1257)
);

A2O1A1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1144),
.A2(n_1066),
.B(n_1050),
.C(n_1063),
.Y(n_1258)
);

O2A1O1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1089),
.A2(n_1055),
.B(n_1124),
.C(n_1126),
.Y(n_1259)
);

AO31x2_ASAP7_75t_L g1260 ( 
.A1(n_1165),
.A2(n_1140),
.A3(n_1110),
.B(n_1125),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1047),
.B(n_1114),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1080),
.B(n_1082),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1061),
.B(n_1130),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1082),
.Y(n_1264)
);

AO31x2_ASAP7_75t_L g1265 ( 
.A1(n_1067),
.A2(n_1104),
.A3(n_1069),
.B(n_1134),
.Y(n_1265)
);

INVx3_ASAP7_75t_L g1266 ( 
.A(n_1080),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1162),
.B(n_1113),
.Y(n_1267)
);

NAND2x1_ASAP7_75t_L g1268 ( 
.A(n_1134),
.B(n_1031),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1051),
.B(n_1162),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_1065),
.B(n_1031),
.Y(n_1270)
);

AO21x2_ASAP7_75t_L g1271 ( 
.A1(n_1121),
.A2(n_1166),
.B(n_1123),
.Y(n_1271)
);

A2O1A1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1090),
.A2(n_1167),
.B(n_1043),
.C(n_1160),
.Y(n_1272)
);

NOR2xp67_ASAP7_75t_L g1273 ( 
.A(n_1043),
.B(n_1160),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1156),
.A2(n_1041),
.B(n_1090),
.Y(n_1274)
);

NOR2x1_ASAP7_75t_SL g1275 ( 
.A(n_1041),
.B(n_1148),
.Y(n_1275)
);

AOI221x1_ASAP7_75t_L g1276 ( 
.A1(n_1084),
.A2(n_1150),
.B1(n_1148),
.B2(n_1143),
.C(n_1116),
.Y(n_1276)
);

BUFx10_ASAP7_75t_L g1277 ( 
.A(n_1060),
.Y(n_1277)
);

A2O1A1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1084),
.A2(n_1150),
.B(n_1127),
.C(n_1138),
.Y(n_1278)
);

A2O1A1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1138),
.A2(n_1143),
.B(n_1148),
.C(n_1051),
.Y(n_1279)
);

INVx1_ASAP7_75t_SL g1280 ( 
.A(n_1138),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1041),
.A2(n_1051),
.B(n_1143),
.Y(n_1281)
);

INVx2_ASAP7_75t_SL g1282 ( 
.A(n_1102),
.Y(n_1282)
);

O2A1O1Ixp33_ASAP7_75t_SL g1283 ( 
.A1(n_1051),
.A2(n_1017),
.B(n_986),
.C(n_1139),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1021),
.Y(n_1284)
);

O2A1O1Ixp33_ASAP7_75t_SL g1285 ( 
.A1(n_1017),
.A2(n_986),
.B(n_1139),
.C(n_1046),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1099),
.A2(n_834),
.B(n_828),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1099),
.A2(n_834),
.B(n_828),
.Y(n_1287)
);

AOI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1115),
.A2(n_979),
.B1(n_985),
.B2(n_967),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1099),
.A2(n_834),
.B(n_828),
.Y(n_1289)
);

AO31x2_ASAP7_75t_L g1290 ( 
.A1(n_1014),
.A2(n_1146),
.A3(n_1171),
.B(n_1109),
.Y(n_1290)
);

BUFx2_ASAP7_75t_R g1291 ( 
.A(n_1060),
.Y(n_1291)
);

NOR2xp67_ASAP7_75t_L g1292 ( 
.A(n_1131),
.B(n_520),
.Y(n_1292)
);

O2A1O1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1017),
.A2(n_979),
.B(n_985),
.C(n_967),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1099),
.A2(n_834),
.B(n_828),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1054),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1054),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1054),
.Y(n_1297)
);

O2A1O1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1017),
.A2(n_979),
.B(n_985),
.C(n_967),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1099),
.A2(n_834),
.B(n_828),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1075),
.A2(n_932),
.B(n_1033),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1021),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1021),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1115),
.B(n_655),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1021),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1021),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1021),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1021),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_1048),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1021),
.Y(n_1309)
);

BUFx5_ASAP7_75t_L g1310 ( 
.A(n_1090),
.Y(n_1310)
);

NAND3xp33_ASAP7_75t_SL g1311 ( 
.A(n_1017),
.B(n_941),
.C(n_1026),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1099),
.A2(n_834),
.B(n_828),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1053),
.B(n_524),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1099),
.A2(n_834),
.B(n_828),
.Y(n_1314)
);

O2A1O1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1017),
.A2(n_979),
.B(n_985),
.C(n_967),
.Y(n_1315)
);

AO21x2_ASAP7_75t_L g1316 ( 
.A1(n_1137),
.A2(n_1017),
.B(n_1018),
.Y(n_1316)
);

AOI211x1_ASAP7_75t_L g1317 ( 
.A1(n_1142),
.A2(n_1158),
.B(n_1056),
.C(n_1136),
.Y(n_1317)
);

A2O1A1Ixp33_ASAP7_75t_L g1318 ( 
.A1(n_1017),
.A2(n_967),
.B(n_985),
.C(n_979),
.Y(n_1318)
);

AOI221x1_ASAP7_75t_L g1319 ( 
.A1(n_1017),
.A2(n_1014),
.B1(n_951),
.B2(n_979),
.C(n_985),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1075),
.A2(n_932),
.B(n_1033),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1115),
.B(n_655),
.Y(n_1321)
);

AOI221x1_ASAP7_75t_L g1322 ( 
.A1(n_1017),
.A2(n_1014),
.B1(n_951),
.B2(n_979),
.C(n_985),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1099),
.A2(n_834),
.B(n_828),
.Y(n_1323)
);

AO31x2_ASAP7_75t_L g1324 ( 
.A1(n_1014),
.A2(n_1146),
.A3(n_1171),
.B(n_1109),
.Y(n_1324)
);

INVx4_ASAP7_75t_L g1325 ( 
.A(n_1172),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1075),
.A2(n_932),
.B(n_1033),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1052),
.B(n_342),
.Y(n_1327)
);

INVx1_ASAP7_75t_SL g1328 ( 
.A(n_1054),
.Y(n_1328)
);

A2O1A1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1017),
.A2(n_967),
.B(n_985),
.C(n_979),
.Y(n_1329)
);

AO31x2_ASAP7_75t_L g1330 ( 
.A1(n_1014),
.A2(n_1146),
.A3(n_1171),
.B(n_1109),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_SL g1331 ( 
.A1(n_1108),
.A2(n_893),
.B(n_830),
.Y(n_1331)
);

NOR2xp67_ASAP7_75t_SL g1332 ( 
.A(n_1131),
.B(n_826),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1075),
.A2(n_932),
.B(n_1033),
.Y(n_1333)
);

A2O1A1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1017),
.A2(n_967),
.B(n_985),
.C(n_979),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1288),
.A2(n_1244),
.B1(n_1177),
.B2(n_1321),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1313),
.B(n_1327),
.Y(n_1336)
);

INVx4_ASAP7_75t_L g1337 ( 
.A(n_1241),
.Y(n_1337)
);

BUFx2_ASAP7_75t_SL g1338 ( 
.A(n_1192),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1303),
.B(n_1288),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_SL g1340 ( 
.A1(n_1222),
.A2(n_1193),
.B1(n_1239),
.B2(n_1247),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_1191),
.Y(n_1341)
);

INVx11_ASAP7_75t_L g1342 ( 
.A(n_1241),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1301),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1305),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_1295),
.Y(n_1345)
);

INVx3_ASAP7_75t_SL g1346 ( 
.A(n_1308),
.Y(n_1346)
);

BUFx8_ASAP7_75t_SL g1347 ( 
.A(n_1296),
.Y(n_1347)
);

CKINVDCx20_ASAP7_75t_R g1348 ( 
.A(n_1184),
.Y(n_1348)
);

OAI22xp33_ASAP7_75t_SL g1349 ( 
.A1(n_1207),
.A2(n_1242),
.B1(n_1180),
.B2(n_1249),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1311),
.A2(n_1230),
.B1(n_1251),
.B2(n_1178),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1318),
.A2(n_1334),
.B1(n_1329),
.B2(n_1298),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1182),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_1297),
.Y(n_1353)
);

CKINVDCx11_ASAP7_75t_R g1354 ( 
.A(n_1277),
.Y(n_1354)
);

INVx11_ASAP7_75t_L g1355 ( 
.A(n_1291),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1325),
.B(n_1175),
.Y(n_1356)
);

BUFx8_ASAP7_75t_SL g1357 ( 
.A(n_1197),
.Y(n_1357)
);

CKINVDCx11_ASAP7_75t_R g1358 ( 
.A(n_1277),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_1221),
.Y(n_1359)
);

INVx8_ASAP7_75t_L g1360 ( 
.A(n_1174),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1187),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1194),
.Y(n_1362)
);

INVx6_ASAP7_75t_L g1363 ( 
.A(n_1325),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1198),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1293),
.A2(n_1315),
.B1(n_1183),
.B2(n_1237),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1261),
.Y(n_1366)
);

BUFx2_ASAP7_75t_L g1367 ( 
.A(n_1179),
.Y(n_1367)
);

BUFx12f_ASAP7_75t_L g1368 ( 
.A(n_1220),
.Y(n_1368)
);

INVx6_ASAP7_75t_L g1369 ( 
.A(n_1174),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1235),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1249),
.A2(n_1212),
.B1(n_1206),
.B2(n_1202),
.Y(n_1371)
);

OAI22xp33_ASAP7_75t_R g1372 ( 
.A1(n_1228),
.A2(n_1282),
.B1(n_1328),
.B2(n_1302),
.Y(n_1372)
);

INVxp67_ASAP7_75t_SL g1373 ( 
.A(n_1269),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1238),
.B(n_1200),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1284),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1304),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_SL g1377 ( 
.A1(n_1310),
.A2(n_1322),
.B1(n_1319),
.B2(n_1331),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1210),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_1210),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1306),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1307),
.Y(n_1381)
);

AOI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1270),
.A2(n_1246),
.B1(n_1201),
.B2(n_1310),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1316),
.A2(n_1208),
.B1(n_1254),
.B2(n_1309),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1245),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_SL g1385 ( 
.A1(n_1310),
.A2(n_1316),
.B1(n_1271),
.B2(n_1283),
.Y(n_1385)
);

AOI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1310),
.A2(n_1271),
.B1(n_1292),
.B2(n_1189),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1181),
.B(n_1256),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1263),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_SL g1389 ( 
.A1(n_1310),
.A2(n_1253),
.B1(n_1275),
.B2(n_1285),
.Y(n_1389)
);

NAND2x1p5_ASAP7_75t_L g1390 ( 
.A(n_1332),
.B(n_1281),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1265),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1262),
.B(n_1280),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1265),
.Y(n_1393)
);

INVx4_ASAP7_75t_L g1394 ( 
.A(n_1188),
.Y(n_1394)
);

BUFx3_ASAP7_75t_L g1395 ( 
.A(n_1188),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1267),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1205),
.B(n_1225),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1276),
.Y(n_1398)
);

BUFx3_ASAP7_75t_L g1399 ( 
.A(n_1188),
.Y(n_1399)
);

BUFx3_ASAP7_75t_L g1400 ( 
.A(n_1262),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1218),
.A2(n_1203),
.B1(n_1229),
.B2(n_1195),
.Y(n_1401)
);

CKINVDCx11_ASAP7_75t_R g1402 ( 
.A(n_1210),
.Y(n_1402)
);

CKINVDCx11_ASAP7_75t_R g1403 ( 
.A(n_1219),
.Y(n_1403)
);

INVx6_ASAP7_75t_L g1404 ( 
.A(n_1219),
.Y(n_1404)
);

BUFx12f_ASAP7_75t_L g1405 ( 
.A(n_1219),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_1236),
.Y(n_1406)
);

BUFx2_ASAP7_75t_L g1407 ( 
.A(n_1236),
.Y(n_1407)
);

INVx1_ASAP7_75t_SL g1408 ( 
.A(n_1236),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1250),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1250),
.B(n_1264),
.Y(n_1410)
);

CKINVDCx8_ASAP7_75t_R g1411 ( 
.A(n_1250),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1317),
.B(n_1292),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1274),
.A2(n_1213),
.B1(n_1317),
.B2(n_1287),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1286),
.A2(n_1294),
.B1(n_1312),
.B2(n_1289),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1258),
.A2(n_1272),
.B1(n_1243),
.B2(n_1278),
.Y(n_1415)
);

AOI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1231),
.A2(n_1233),
.B1(n_1217),
.B2(n_1266),
.Y(n_1416)
);

INVx4_ASAP7_75t_L g1417 ( 
.A(n_1264),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_SL g1418 ( 
.A1(n_1252),
.A2(n_1290),
.B1(n_1330),
.B2(n_1324),
.Y(n_1418)
);

INVx4_ASAP7_75t_L g1419 ( 
.A(n_1264),
.Y(n_1419)
);

AOI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1217),
.A2(n_1273),
.B1(n_1176),
.B2(n_1248),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_SL g1421 ( 
.A1(n_1290),
.A2(n_1330),
.B1(n_1324),
.B2(n_1240),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_SL g1422 ( 
.A1(n_1290),
.A2(n_1330),
.B1(n_1324),
.B2(n_1257),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1259),
.B(n_1232),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1232),
.B(n_1190),
.Y(n_1424)
);

OAI21xp33_ASAP7_75t_L g1425 ( 
.A1(n_1279),
.A2(n_1299),
.B(n_1314),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1248),
.B(n_1268),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1260),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1323),
.A2(n_1216),
.B1(n_1255),
.B2(n_1223),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_SL g1429 ( 
.A1(n_1226),
.A2(n_1199),
.B1(n_1227),
.B2(n_1211),
.Y(n_1429)
);

BUFx2_ASAP7_75t_SL g1430 ( 
.A(n_1224),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1196),
.A2(n_1186),
.B1(n_1209),
.B2(n_1326),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1185),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1214),
.A2(n_1199),
.B1(n_1232),
.B2(n_1227),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1199),
.A2(n_1227),
.B1(n_1204),
.B2(n_1185),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1185),
.A2(n_1215),
.B1(n_1234),
.B2(n_1333),
.Y(n_1435)
);

BUFx2_ASAP7_75t_L g1436 ( 
.A(n_1215),
.Y(n_1436)
);

BUFx10_ASAP7_75t_L g1437 ( 
.A(n_1234),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1234),
.B(n_1300),
.Y(n_1438)
);

BUFx3_ASAP7_75t_L g1439 ( 
.A(n_1320),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1192),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1318),
.A2(n_1334),
.B(n_1329),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1301),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1301),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1269),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1303),
.B(n_1321),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_SL g1446 ( 
.A(n_1291),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1301),
.Y(n_1447)
);

INVx1_ASAP7_75t_SL g1448 ( 
.A(n_1328),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1288),
.A2(n_967),
.B1(n_985),
.B2(n_979),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1288),
.A2(n_967),
.B1(n_985),
.B2(n_979),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_SL g1451 ( 
.A1(n_1244),
.A2(n_745),
.B1(n_941),
.B2(n_669),
.Y(n_1451)
);

INVx1_ASAP7_75t_SL g1452 ( 
.A(n_1328),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1301),
.Y(n_1453)
);

INVx4_ASAP7_75t_L g1454 ( 
.A(n_1241),
.Y(n_1454)
);

INVx1_ASAP7_75t_SL g1455 ( 
.A(n_1328),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1288),
.A2(n_967),
.B1(n_985),
.B2(n_979),
.Y(n_1456)
);

AOI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1318),
.A2(n_1334),
.B(n_1329),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1288),
.A2(n_1318),
.B1(n_1334),
.B2(n_1329),
.Y(n_1458)
);

INVx6_ASAP7_75t_L g1459 ( 
.A(n_1325),
.Y(n_1459)
);

CKINVDCx6p67_ASAP7_75t_R g1460 ( 
.A(n_1184),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1301),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1301),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1303),
.B(n_1321),
.Y(n_1463)
);

CKINVDCx11_ASAP7_75t_R g1464 ( 
.A(n_1184),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1313),
.B(n_1177),
.Y(n_1465)
);

AOI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1288),
.A2(n_448),
.B1(n_352),
.B2(n_361),
.Y(n_1466)
);

INVx5_ASAP7_75t_L g1467 ( 
.A(n_1241),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1301),
.Y(n_1468)
);

BUFx4f_ASAP7_75t_L g1469 ( 
.A(n_1241),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1192),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_SL g1471 ( 
.A1(n_1244),
.A2(n_745),
.B1(n_941),
.B2(n_669),
.Y(n_1471)
);

BUFx8_ASAP7_75t_L g1472 ( 
.A(n_1282),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1424),
.B(n_1444),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1391),
.Y(n_1474)
);

OAI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1449),
.A2(n_1456),
.B1(n_1450),
.B2(n_1451),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1393),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1427),
.Y(n_1477)
);

INVxp67_ASAP7_75t_SL g1478 ( 
.A(n_1444),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1373),
.B(n_1432),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1386),
.B(n_1373),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1449),
.A2(n_1450),
.B1(n_1456),
.B2(n_1471),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1439),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1458),
.A2(n_1457),
.B(n_1441),
.Y(n_1483)
);

OA21x2_ASAP7_75t_L g1484 ( 
.A1(n_1423),
.A2(n_1413),
.B(n_1414),
.Y(n_1484)
);

OAI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1351),
.A2(n_1471),
.B(n_1451),
.Y(n_1485)
);

BUFx3_ASAP7_75t_L g1486 ( 
.A(n_1390),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1436),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1421),
.B(n_1397),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1434),
.Y(n_1489)
);

CKINVDCx20_ASAP7_75t_R g1490 ( 
.A(n_1464),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1433),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1421),
.B(n_1422),
.Y(n_1492)
);

OAI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1466),
.A2(n_1339),
.B1(n_1382),
.B2(n_1463),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_SL g1494 ( 
.A1(n_1340),
.A2(n_1415),
.B1(n_1349),
.B2(n_1365),
.Y(n_1494)
);

OA21x2_ASAP7_75t_L g1495 ( 
.A1(n_1413),
.A2(n_1414),
.B(n_1438),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1422),
.B(n_1371),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1352),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1361),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1362),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1341),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1341),
.Y(n_1501)
);

AOI222xp33_ASAP7_75t_L g1502 ( 
.A1(n_1335),
.A2(n_1445),
.B1(n_1371),
.B2(n_1465),
.C1(n_1372),
.C2(n_1350),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1364),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1428),
.A2(n_1425),
.B(n_1401),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1437),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1370),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1383),
.B(n_1462),
.Y(n_1507)
);

NAND4xp25_ASAP7_75t_L g1508 ( 
.A(n_1335),
.B(n_1350),
.C(n_1388),
.D(n_1374),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1376),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1431),
.A2(n_1428),
.B(n_1435),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1381),
.Y(n_1511)
);

OA21x2_ASAP7_75t_L g1512 ( 
.A1(n_1383),
.A2(n_1401),
.B(n_1431),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1396),
.B(n_1387),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1390),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1377),
.B(n_1418),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1384),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1375),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1430),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1398),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1380),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1377),
.B(n_1418),
.Y(n_1521)
);

AO21x2_ASAP7_75t_L g1522 ( 
.A1(n_1416),
.A2(n_1420),
.B(n_1412),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1366),
.B(n_1385),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1343),
.Y(n_1524)
);

OAI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1448),
.A2(n_1452),
.B1(n_1455),
.B2(n_1470),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1447),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1453),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1394),
.Y(n_1528)
);

AOI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1389),
.A2(n_1385),
.B(n_1429),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1394),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1461),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_L g1532 ( 
.A1(n_1468),
.A2(n_1442),
.B(n_1443),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1429),
.Y(n_1533)
);

BUFx2_ASAP7_75t_L g1534 ( 
.A(n_1359),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1400),
.B(n_1344),
.Y(n_1535)
);

BUFx3_ASAP7_75t_L g1536 ( 
.A(n_1360),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1389),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1426),
.Y(n_1538)
);

OAI21x1_ASAP7_75t_L g1539 ( 
.A1(n_1410),
.A2(n_1336),
.B(n_1360),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1356),
.B(n_1392),
.Y(n_1540)
);

OA21x2_ASAP7_75t_L g1541 ( 
.A1(n_1407),
.A2(n_1392),
.B(n_1408),
.Y(n_1541)
);

OAI21x1_ASAP7_75t_L g1542 ( 
.A1(n_1360),
.A2(n_1467),
.B(n_1369),
.Y(n_1542)
);

AOI21x1_ASAP7_75t_L g1543 ( 
.A1(n_1356),
.A2(n_1353),
.B(n_1440),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_SL g1544 ( 
.A1(n_1338),
.A2(n_1363),
.B1(n_1459),
.B2(n_1345),
.Y(n_1544)
);

OAI21x1_ASAP7_75t_L g1545 ( 
.A1(n_1467),
.A2(n_1369),
.B(n_1399),
.Y(n_1545)
);

AO21x1_ASAP7_75t_L g1546 ( 
.A1(n_1417),
.A2(n_1419),
.B(n_1337),
.Y(n_1546)
);

INVxp67_ASAP7_75t_L g1547 ( 
.A(n_1367),
.Y(n_1547)
);

BUFx2_ASAP7_75t_L g1548 ( 
.A(n_1395),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1395),
.Y(n_1549)
);

AOI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1399),
.A2(n_1411),
.B(n_1404),
.Y(n_1550)
);

BUFx3_ASAP7_75t_L g1551 ( 
.A(n_1345),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1409),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1467),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_L g1554 ( 
.A(n_1357),
.B(n_1346),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1419),
.B(n_1467),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1363),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1357),
.Y(n_1557)
);

OAI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1446),
.A2(n_1469),
.B1(n_1379),
.B2(n_1406),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1363),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1459),
.A2(n_1469),
.B(n_1403),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1378),
.B(n_1402),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_SL g1562 ( 
.A(n_1446),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1459),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1402),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1403),
.Y(n_1565)
);

AOI221xp5_ASAP7_75t_L g1566 ( 
.A1(n_1475),
.A2(n_1337),
.B1(n_1454),
.B2(n_1346),
.C(n_1348),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1483),
.A2(n_1405),
.B(n_1342),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1493),
.B(n_1347),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1538),
.B(n_1354),
.Y(n_1569)
);

AND2x4_ASAP7_75t_SL g1570 ( 
.A(n_1561),
.B(n_1460),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1538),
.B(n_1354),
.Y(n_1571)
);

OAI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1475),
.A2(n_1358),
.B(n_1347),
.Y(n_1572)
);

A2O1A1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1485),
.A2(n_1358),
.B(n_1355),
.C(n_1472),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1486),
.B(n_1472),
.Y(n_1574)
);

BUFx4f_ASAP7_75t_L g1575 ( 
.A(n_1561),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1497),
.Y(n_1576)
);

OAI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1485),
.A2(n_1368),
.B(n_1464),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1523),
.B(n_1488),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1478),
.B(n_1473),
.Y(n_1579)
);

BUFx2_ASAP7_75t_R g1580 ( 
.A(n_1540),
.Y(n_1580)
);

O2A1O1Ixp33_ASAP7_75t_L g1581 ( 
.A1(n_1502),
.A2(n_1481),
.B(n_1508),
.C(n_1504),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1473),
.B(n_1488),
.Y(n_1582)
);

OAI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1494),
.A2(n_1515),
.B1(n_1513),
.B2(n_1496),
.Y(n_1583)
);

AOI21xp5_ASAP7_75t_SL g1584 ( 
.A1(n_1558),
.A2(n_1555),
.B(n_1536),
.Y(n_1584)
);

O2A1O1Ixp33_ASAP7_75t_L g1585 ( 
.A1(n_1502),
.A2(n_1508),
.B(n_1525),
.C(n_1513),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1523),
.B(n_1517),
.Y(n_1586)
);

A2O1A1Ixp33_ASAP7_75t_L g1587 ( 
.A1(n_1529),
.A2(n_1496),
.B(n_1537),
.C(n_1515),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1498),
.B(n_1499),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1540),
.B(n_1541),
.Y(n_1589)
);

OAI21xp33_ASAP7_75t_L g1590 ( 
.A1(n_1521),
.A2(n_1492),
.B(n_1491),
.Y(n_1590)
);

NAND2xp33_ASAP7_75t_R g1591 ( 
.A(n_1554),
.B(n_1534),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1541),
.B(n_1526),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1541),
.B(n_1552),
.Y(n_1593)
);

OAI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1480),
.A2(n_1510),
.B(n_1537),
.Y(n_1594)
);

NOR2x1_ASAP7_75t_SL g1595 ( 
.A(n_1543),
.B(n_1522),
.Y(n_1595)
);

CKINVDCx20_ASAP7_75t_R g1596 ( 
.A(n_1490),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1541),
.B(n_1552),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1479),
.B(n_1519),
.Y(n_1598)
);

OAI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1480),
.A2(n_1510),
.B(n_1543),
.Y(n_1599)
);

AOI22xp5_ASAP7_75t_SL g1600 ( 
.A1(n_1558),
.A2(n_1557),
.B1(n_1564),
.B2(n_1565),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1547),
.B(n_1562),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1498),
.Y(n_1602)
);

O2A1O1Ixp33_ASAP7_75t_SL g1603 ( 
.A1(n_1555),
.A2(n_1549),
.B(n_1564),
.C(n_1565),
.Y(n_1603)
);

OAI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1480),
.A2(n_1512),
.B(n_1484),
.Y(n_1604)
);

OA21x2_ASAP7_75t_L g1605 ( 
.A1(n_1489),
.A2(n_1518),
.B(n_1491),
.Y(n_1605)
);

OA21x2_ASAP7_75t_L g1606 ( 
.A1(n_1489),
.A2(n_1518),
.B(n_1533),
.Y(n_1606)
);

OAI211xp5_ASAP7_75t_L g1607 ( 
.A1(n_1521),
.A2(n_1500),
.B(n_1501),
.C(n_1544),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_SL g1608 ( 
.A1(n_1564),
.A2(n_1565),
.B1(n_1551),
.B2(n_1534),
.Y(n_1608)
);

A2O1A1Ixp33_ASAP7_75t_L g1609 ( 
.A1(n_1480),
.A2(n_1560),
.B(n_1539),
.C(n_1545),
.Y(n_1609)
);

NAND3xp33_ASAP7_75t_L g1610 ( 
.A(n_1520),
.B(n_1531),
.C(n_1527),
.Y(n_1610)
);

A2O1A1Ixp33_ASAP7_75t_L g1611 ( 
.A1(n_1560),
.A2(n_1539),
.B(n_1545),
.C(n_1542),
.Y(n_1611)
);

NOR2x1_ASAP7_75t_SL g1612 ( 
.A(n_1522),
.B(n_1550),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1503),
.B(n_1506),
.Y(n_1613)
);

A2O1A1Ixp33_ASAP7_75t_SL g1614 ( 
.A1(n_1553),
.A2(n_1528),
.B(n_1530),
.C(n_1556),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1503),
.B(n_1506),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1535),
.B(n_1520),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1535),
.B(n_1524),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1509),
.B(n_1511),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1486),
.B(n_1514),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_SL g1620 ( 
.A1(n_1522),
.A2(n_1512),
.B1(n_1484),
.B2(n_1514),
.Y(n_1620)
);

OA21x2_ASAP7_75t_L g1621 ( 
.A1(n_1474),
.A2(n_1476),
.B(n_1477),
.Y(n_1621)
);

OAI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1512),
.A2(n_1484),
.B(n_1532),
.Y(n_1622)
);

OR2x6_ASAP7_75t_L g1623 ( 
.A(n_1542),
.B(n_1505),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1516),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_SL g1625 ( 
.A(n_1585),
.B(n_1563),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1606),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1579),
.B(n_1507),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1606),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1604),
.B(n_1495),
.Y(n_1629)
);

INVx3_ASAP7_75t_L g1630 ( 
.A(n_1621),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1621),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1623),
.B(n_1482),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1579),
.B(n_1507),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1583),
.A2(n_1522),
.B1(n_1484),
.B2(n_1512),
.Y(n_1634)
);

OAI221xp5_ASAP7_75t_L g1635 ( 
.A1(n_1572),
.A2(n_1563),
.B1(n_1559),
.B2(n_1556),
.C(n_1495),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1582),
.B(n_1487),
.Y(n_1636)
);

BUFx2_ASAP7_75t_L g1637 ( 
.A(n_1592),
.Y(n_1637)
);

INVx2_ASAP7_75t_SL g1638 ( 
.A(n_1593),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1576),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1583),
.B(n_1581),
.Y(n_1640)
);

BUFx6f_ASAP7_75t_L g1641 ( 
.A(n_1623),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1611),
.B(n_1609),
.Y(n_1642)
);

INVx3_ASAP7_75t_L g1643 ( 
.A(n_1605),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1602),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1604),
.B(n_1495),
.Y(n_1645)
);

BUFx2_ASAP7_75t_L g1646 ( 
.A(n_1597),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1594),
.B(n_1589),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1624),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1610),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1605),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1613),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1613),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1615),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1615),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1618),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1607),
.B(n_1590),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1647),
.B(n_1599),
.Y(n_1657)
);

OAI21xp5_ASAP7_75t_SL g1658 ( 
.A1(n_1640),
.A2(n_1577),
.B(n_1572),
.Y(n_1658)
);

AOI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1640),
.A2(n_1587),
.B1(n_1577),
.B2(n_1568),
.C(n_1566),
.Y(n_1659)
);

AOI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1656),
.A2(n_1566),
.B1(n_1591),
.B2(n_1569),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1630),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1647),
.B(n_1599),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1647),
.B(n_1638),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1630),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1626),
.B(n_1628),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1649),
.B(n_1627),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1638),
.B(n_1620),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1649),
.B(n_1578),
.Y(n_1668)
);

AND2x4_ASAP7_75t_L g1669 ( 
.A(n_1632),
.B(n_1619),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1627),
.B(n_1598),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1644),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1634),
.A2(n_1622),
.B(n_1595),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1646),
.B(n_1586),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1644),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1648),
.Y(n_1675)
);

BUFx3_ASAP7_75t_L g1676 ( 
.A(n_1641),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1633),
.B(n_1651),
.Y(n_1677)
);

INVx2_ASAP7_75t_SL g1678 ( 
.A(n_1641),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1630),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1656),
.A2(n_1569),
.B1(n_1571),
.B2(n_1575),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1626),
.B(n_1588),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1629),
.B(n_1617),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1629),
.B(n_1612),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1629),
.B(n_1616),
.Y(n_1684)
);

INVx4_ASAP7_75t_L g1685 ( 
.A(n_1641),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1630),
.Y(n_1686)
);

NOR2x1_ASAP7_75t_L g1687 ( 
.A(n_1643),
.B(n_1584),
.Y(n_1687)
);

CKINVDCx16_ASAP7_75t_R g1688 ( 
.A(n_1642),
.Y(n_1688)
);

INVx2_ASAP7_75t_SL g1689 ( 
.A(n_1641),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1631),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1639),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1685),
.B(n_1641),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1657),
.B(n_1637),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1666),
.B(n_1652),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1691),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1691),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1671),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1657),
.B(n_1637),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1657),
.B(n_1645),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1671),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1666),
.B(n_1652),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1668),
.B(n_1653),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1662),
.B(n_1645),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1668),
.B(n_1653),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1677),
.B(n_1636),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1677),
.B(n_1654),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1690),
.Y(n_1707)
);

INVx2_ASAP7_75t_SL g1708 ( 
.A(n_1676),
.Y(n_1708)
);

BUFx3_ASAP7_75t_L g1709 ( 
.A(n_1676),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1665),
.Y(n_1710)
);

NOR4xp25_ASAP7_75t_SL g1711 ( 
.A(n_1658),
.B(n_1603),
.C(n_1635),
.D(n_1625),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_SL g1712 ( 
.A(n_1688),
.B(n_1575),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1662),
.B(n_1642),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1660),
.A2(n_1634),
.B1(n_1580),
.B2(n_1600),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1662),
.B(n_1642),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_SL g1716 ( 
.A(n_1688),
.B(n_1642),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1674),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1690),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1663),
.B(n_1683),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1670),
.B(n_1654),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1681),
.B(n_1636),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1685),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1674),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1675),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1670),
.B(n_1655),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1663),
.B(n_1642),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1663),
.B(n_1641),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1665),
.B(n_1650),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1713),
.B(n_1683),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1702),
.B(n_1684),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1702),
.B(n_1684),
.Y(n_1731)
);

NAND3xp33_ASAP7_75t_L g1732 ( 
.A(n_1711),
.B(n_1659),
.C(n_1658),
.Y(n_1732)
);

NOR2x1p5_ASAP7_75t_L g1733 ( 
.A(n_1709),
.B(n_1676),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1695),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1713),
.B(n_1683),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1704),
.B(n_1684),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1713),
.B(n_1715),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1719),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1721),
.B(n_1705),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1704),
.B(n_1682),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1721),
.B(n_1665),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1719),
.Y(n_1742)
);

O2A1O1Ixp5_ASAP7_75t_SL g1743 ( 
.A1(n_1722),
.A2(n_1714),
.B(n_1710),
.C(n_1716),
.Y(n_1743)
);

NAND4xp25_ASAP7_75t_SL g1744 ( 
.A(n_1715),
.B(n_1659),
.C(n_1660),
.D(n_1687),
.Y(n_1744)
);

OAI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1714),
.A2(n_1635),
.B1(n_1672),
.B2(n_1685),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1715),
.B(n_1669),
.Y(n_1746)
);

HB1xp67_ASAP7_75t_L g1747 ( 
.A(n_1710),
.Y(n_1747)
);

INVxp67_ASAP7_75t_L g1748 ( 
.A(n_1694),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1726),
.B(n_1687),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1695),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1720),
.B(n_1682),
.Y(n_1751)
);

INVx1_ASAP7_75t_SL g1752 ( 
.A(n_1709),
.Y(n_1752)
);

INVx2_ASAP7_75t_SL g1753 ( 
.A(n_1722),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1696),
.Y(n_1754)
);

OAI21xp33_ASAP7_75t_L g1755 ( 
.A1(n_1726),
.A2(n_1672),
.B(n_1667),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1726),
.B(n_1669),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1696),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1697),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1697),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1693),
.B(n_1669),
.Y(n_1760)
);

NAND3xp33_ASAP7_75t_SL g1761 ( 
.A(n_1711),
.B(n_1680),
.C(n_1685),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1720),
.B(n_1682),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1725),
.B(n_1705),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1725),
.B(n_1667),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1694),
.B(n_1667),
.Y(n_1765)
);

AND2x4_ASAP7_75t_L g1766 ( 
.A(n_1709),
.B(n_1685),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1693),
.B(n_1669),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1701),
.B(n_1706),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1693),
.B(n_1698),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1701),
.B(n_1681),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1698),
.B(n_1669),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1737),
.B(n_1719),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1747),
.B(n_1748),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_L g1774 ( 
.A(n_1769),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1738),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1768),
.B(n_1765),
.Y(n_1776)
);

AND2x4_ASAP7_75t_L g1777 ( 
.A(n_1733),
.B(n_1722),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_SL g1778 ( 
.A(n_1732),
.B(n_1580),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1737),
.B(n_1708),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1769),
.B(n_1708),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1752),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1744),
.B(n_1596),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1734),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1746),
.B(n_1708),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1746),
.B(n_1722),
.Y(n_1785)
);

NAND2x1p5_ASAP7_75t_L g1786 ( 
.A(n_1733),
.B(n_1712),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1764),
.B(n_1706),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1734),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1768),
.B(n_1763),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1756),
.B(n_1727),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1745),
.A2(n_1692),
.B1(n_1680),
.B2(n_1727),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1750),
.Y(n_1792)
);

INVx1_ASAP7_75t_SL g1793 ( 
.A(n_1766),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1756),
.B(n_1727),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1750),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1749),
.B(n_1692),
.Y(n_1796)
);

AND2x4_ASAP7_75t_L g1797 ( 
.A(n_1749),
.B(n_1692),
.Y(n_1797)
);

NAND2xp33_ASAP7_75t_L g1798 ( 
.A(n_1755),
.B(n_1608),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1754),
.B(n_1699),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1754),
.B(n_1699),
.Y(n_1800)
);

AOI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1761),
.A2(n_1573),
.B(n_1567),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1739),
.B(n_1728),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1739),
.B(n_1728),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1757),
.B(n_1699),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1738),
.Y(n_1805)
);

INVx1_ASAP7_75t_SL g1806 ( 
.A(n_1766),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1751),
.B(n_1728),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_SL g1808 ( 
.A1(n_1801),
.A2(n_1743),
.B(n_1749),
.Y(n_1808)
);

INVxp67_ASAP7_75t_SL g1809 ( 
.A(n_1781),
.Y(n_1809)
);

AOI221xp5_ASAP7_75t_L g1810 ( 
.A1(n_1798),
.A2(n_1743),
.B1(n_1742),
.B2(n_1757),
.C(n_1759),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1779),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1793),
.B(n_1729),
.Y(n_1812)
);

NOR4xp25_ASAP7_75t_SL g1813 ( 
.A(n_1783),
.B(n_1758),
.C(n_1759),
.D(n_1766),
.Y(n_1813)
);

NAND4xp75_ASAP7_75t_L g1814 ( 
.A(n_1782),
.B(n_1753),
.C(n_1567),
.D(n_1546),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1786),
.B(n_1780),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1783),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1788),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1793),
.B(n_1729),
.Y(n_1818)
);

INVx1_ASAP7_75t_SL g1819 ( 
.A(n_1806),
.Y(n_1819)
);

AOI222xp33_ASAP7_75t_L g1820 ( 
.A1(n_1778),
.A2(n_1742),
.B1(n_1703),
.B2(n_1771),
.C1(n_1760),
.C2(n_1767),
.Y(n_1820)
);

NAND2x1_ASAP7_75t_L g1821 ( 
.A(n_1777),
.B(n_1753),
.Y(n_1821)
);

NAND3xp33_ASAP7_75t_L g1822 ( 
.A(n_1778),
.B(n_1741),
.C(n_1758),
.Y(n_1822)
);

OA21x2_ASAP7_75t_L g1823 ( 
.A1(n_1791),
.A2(n_1805),
.B(n_1775),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1806),
.B(n_1735),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1774),
.B(n_1735),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1788),
.Y(n_1826)
);

AOI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1786),
.A2(n_1796),
.B1(n_1797),
.B2(n_1777),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1792),
.Y(n_1828)
);

AOI22xp5_ASAP7_75t_SL g1829 ( 
.A1(n_1777),
.A2(n_1692),
.B1(n_1601),
.B2(n_1676),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1773),
.B(n_1760),
.Y(n_1830)
);

BUFx2_ASAP7_75t_L g1831 ( 
.A(n_1777),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1792),
.Y(n_1832)
);

OAI22xp5_ASAP7_75t_L g1833 ( 
.A1(n_1786),
.A2(n_1771),
.B1(n_1767),
.B2(n_1730),
.Y(n_1833)
);

INVxp67_ASAP7_75t_L g1834 ( 
.A(n_1809),
.Y(n_1834)
);

HB1xp67_ASAP7_75t_L g1835 ( 
.A(n_1831),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1816),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_SL g1837 ( 
.A(n_1829),
.B(n_1797),
.Y(n_1837)
);

OAI21x1_ASAP7_75t_SL g1838 ( 
.A1(n_1827),
.A2(n_1773),
.B(n_1775),
.Y(n_1838)
);

AOI22xp5_ASAP7_75t_L g1839 ( 
.A1(n_1822),
.A2(n_1796),
.B1(n_1797),
.B2(n_1780),
.Y(n_1839)
);

INVx1_ASAP7_75t_SL g1840 ( 
.A(n_1831),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1819),
.B(n_1790),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1830),
.B(n_1789),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1815),
.B(n_1790),
.Y(n_1843)
);

AOI322xp5_ASAP7_75t_L g1844 ( 
.A1(n_1810),
.A2(n_1789),
.A3(n_1772),
.B1(n_1787),
.B2(n_1703),
.C1(n_1794),
.C2(n_1800),
.Y(n_1844)
);

AOI32xp33_ASAP7_75t_L g1845 ( 
.A1(n_1815),
.A2(n_1797),
.A3(n_1779),
.B1(n_1784),
.B2(n_1794),
.Y(n_1845)
);

AOI21xp33_ASAP7_75t_L g1846 ( 
.A1(n_1823),
.A2(n_1776),
.B(n_1787),
.Y(n_1846)
);

AOI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1820),
.A2(n_1784),
.B1(n_1785),
.B2(n_1692),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1811),
.B(n_1772),
.Y(n_1848)
);

AOI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1823),
.A2(n_1785),
.B1(n_1776),
.B2(n_1804),
.Y(n_1849)
);

OAI21xp33_ASAP7_75t_L g1850 ( 
.A1(n_1808),
.A2(n_1799),
.B(n_1804),
.Y(n_1850)
);

INVx1_ASAP7_75t_SL g1851 ( 
.A(n_1811),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1823),
.B(n_1812),
.Y(n_1852)
);

AOI21xp33_ASAP7_75t_L g1853 ( 
.A1(n_1821),
.A2(n_1775),
.B(n_1805),
.Y(n_1853)
);

AOI221xp5_ASAP7_75t_L g1854 ( 
.A1(n_1846),
.A2(n_1808),
.B1(n_1833),
.B2(n_1824),
.C(n_1818),
.Y(n_1854)
);

NOR3xp33_ASAP7_75t_SL g1855 ( 
.A(n_1850),
.B(n_1814),
.C(n_1825),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1843),
.B(n_1813),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1841),
.B(n_1802),
.Y(n_1857)
);

XNOR2x1_ASAP7_75t_L g1858 ( 
.A(n_1842),
.B(n_1814),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1834),
.B(n_1817),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1848),
.B(n_1802),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1835),
.Y(n_1861)
);

OAI321xp33_ASAP7_75t_L g1862 ( 
.A1(n_1852),
.A2(n_1837),
.A3(n_1839),
.B1(n_1845),
.B2(n_1849),
.C(n_1847),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1851),
.B(n_1840),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1840),
.Y(n_1864)
);

AOI21xp33_ASAP7_75t_L g1865 ( 
.A1(n_1838),
.A2(n_1832),
.B(n_1828),
.Y(n_1865)
);

OAI22x1_ASAP7_75t_L g1866 ( 
.A1(n_1836),
.A2(n_1826),
.B1(n_1805),
.B2(n_1795),
.Y(n_1866)
);

AOI31xp33_ASAP7_75t_L g1867 ( 
.A1(n_1864),
.A2(n_1853),
.A3(n_1803),
.B(n_1795),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1863),
.B(n_1844),
.Y(n_1868)
);

NAND3xp33_ASAP7_75t_SL g1869 ( 
.A(n_1854),
.B(n_1803),
.C(n_1800),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_SL g1870 ( 
.A(n_1862),
.B(n_1799),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1861),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1856),
.B(n_1703),
.Y(n_1872)
);

AOI211x1_ASAP7_75t_L g1873 ( 
.A1(n_1865),
.A2(n_1859),
.B(n_1862),
.C(n_1855),
.Y(n_1873)
);

NOR3xp33_ASAP7_75t_SL g1874 ( 
.A(n_1865),
.B(n_1762),
.C(n_1731),
.Y(n_1874)
);

NOR2x1_ASAP7_75t_L g1875 ( 
.A(n_1858),
.B(n_1741),
.Y(n_1875)
);

OAI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1857),
.A2(n_1807),
.B(n_1770),
.Y(n_1876)
);

OAI21xp33_ASAP7_75t_SL g1877 ( 
.A1(n_1860),
.A2(n_1807),
.B(n_1736),
.Y(n_1877)
);

AOI211xp5_ASAP7_75t_L g1878 ( 
.A1(n_1870),
.A2(n_1868),
.B(n_1869),
.C(n_1871),
.Y(n_1878)
);

AOI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1867),
.A2(n_1866),
.B(n_1570),
.Y(n_1879)
);

AOI221xp5_ASAP7_75t_L g1880 ( 
.A1(n_1873),
.A2(n_1689),
.B1(n_1678),
.B2(n_1740),
.C(n_1770),
.Y(n_1880)
);

AOI311xp33_ASAP7_75t_L g1881 ( 
.A1(n_1872),
.A2(n_1724),
.A3(n_1723),
.B(n_1700),
.C(n_1717),
.Y(n_1881)
);

AOI221xp5_ASAP7_75t_L g1882 ( 
.A1(n_1867),
.A2(n_1678),
.B1(n_1689),
.B2(n_1698),
.C(n_1679),
.Y(n_1882)
);

NOR3xp33_ASAP7_75t_L g1883 ( 
.A(n_1878),
.B(n_1875),
.C(n_1877),
.Y(n_1883)
);

AOI221xp5_ASAP7_75t_L g1884 ( 
.A1(n_1879),
.A2(n_1874),
.B1(n_1876),
.B2(n_1678),
.C(n_1689),
.Y(n_1884)
);

NAND4xp25_ASAP7_75t_L g1885 ( 
.A(n_1880),
.B(n_1574),
.C(n_1571),
.D(n_1536),
.Y(n_1885)
);

NOR3xp33_ASAP7_75t_L g1886 ( 
.A(n_1882),
.B(n_1574),
.C(n_1553),
.Y(n_1886)
);

AOI21xp5_ASAP7_75t_L g1887 ( 
.A1(n_1881),
.A2(n_1718),
.B(n_1707),
.Y(n_1887)
);

AOI221x1_ASAP7_75t_L g1888 ( 
.A1(n_1879),
.A2(n_1707),
.B1(n_1718),
.B2(n_1679),
.C(n_1664),
.Y(n_1888)
);

XNOR2x1_ASAP7_75t_L g1889 ( 
.A(n_1883),
.B(n_1536),
.Y(n_1889)
);

NOR2x1_ASAP7_75t_L g1890 ( 
.A(n_1885),
.B(n_1707),
.Y(n_1890)
);

NOR2x1_ASAP7_75t_L g1891 ( 
.A(n_1887),
.B(n_1718),
.Y(n_1891)
);

NAND4xp75_ASAP7_75t_L g1892 ( 
.A(n_1888),
.B(n_1884),
.C(n_1886),
.D(n_1546),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1883),
.Y(n_1893)
);

AOI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1893),
.A2(n_1679),
.B(n_1661),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1889),
.B(n_1673),
.Y(n_1895)
);

OR2x2_ASAP7_75t_L g1896 ( 
.A(n_1892),
.B(n_1679),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1895),
.Y(n_1897)
);

INVxp67_ASAP7_75t_SL g1898 ( 
.A(n_1897),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1898),
.Y(n_1899)
);

INVx3_ASAP7_75t_SL g1900 ( 
.A(n_1898),
.Y(n_1900)
);

AO22x2_ASAP7_75t_L g1901 ( 
.A1(n_1899),
.A2(n_1896),
.B1(n_1894),
.B2(n_1891),
.Y(n_1901)
);

OAI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1900),
.A2(n_1890),
.B1(n_1686),
.B2(n_1661),
.Y(n_1902)
);

AO21x2_ASAP7_75t_L g1903 ( 
.A1(n_1902),
.A2(n_1686),
.B(n_1664),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1901),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1904),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1905),
.B(n_1903),
.Y(n_1906)
);

XNOR2xp5_ASAP7_75t_L g1907 ( 
.A(n_1906),
.B(n_1903),
.Y(n_1907)
);

AOI22xp33_ASAP7_75t_L g1908 ( 
.A1(n_1907),
.A2(n_1686),
.B1(n_1664),
.B2(n_1661),
.Y(n_1908)
);

AOI211xp5_ASAP7_75t_L g1909 ( 
.A1(n_1908),
.A2(n_1548),
.B(n_1553),
.C(n_1614),
.Y(n_1909)
);


endmodule