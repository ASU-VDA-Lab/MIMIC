module fake_jpeg_30204_n_538 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_538);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_538;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_8),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_18),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_54),
.B(n_56),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_17),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_55),
.B(n_69),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_24),
.B(n_15),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_59),
.Y(n_142)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_61),
.Y(n_165)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_24),
.B(n_15),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_64),
.B(n_79),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_32),
.B(n_17),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_65),
.B(n_76),
.Y(n_123)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_68),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_32),
.B(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_72),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_75),
.Y(n_149)
);

BUFx4f_ASAP7_75t_SL g76 ( 
.A(n_43),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_99),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_17),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_0),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_80),
.B(n_81),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_0),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_26),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_22),
.B(n_0),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_22),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_93),
.Y(n_161)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_19),
.Y(n_95)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_19),
.Y(n_98)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

BUFx12_ASAP7_75t_L g99 ( 
.A(n_19),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_35),
.Y(n_100)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_101),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_38),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_58),
.A2(n_21),
.B1(n_38),
.B2(n_28),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_114),
.A2(n_127),
.B1(n_157),
.B2(n_145),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_117),
.B(n_125),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_80),
.A2(n_21),
.B1(n_36),
.B2(n_49),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_122),
.A2(n_140),
.B1(n_3),
.B2(n_4),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_54),
.B(n_49),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_81),
.A2(n_21),
.B1(n_36),
.B2(n_39),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_56),
.A2(n_36),
.B1(n_34),
.B2(n_37),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_144),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_88),
.A2(n_30),
.B1(n_35),
.B2(n_28),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_145),
.A2(n_155),
.B1(n_159),
.B2(n_83),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_64),
.B(n_41),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_146),
.B(n_150),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_79),
.B(n_39),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_91),
.Y(n_151)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_151),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_57),
.A2(n_30),
.B1(n_35),
.B2(n_28),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_78),
.B(n_41),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_164),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_67),
.A2(n_28),
.B1(n_38),
.B2(n_42),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_102),
.A2(n_30),
.B1(n_38),
.B2(n_28),
.Y(n_159)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_70),
.Y(n_162)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_162),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_76),
.B(n_37),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_166),
.A2(n_191),
.B1(n_188),
.B2(n_222),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_108),
.B(n_34),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_167),
.B(n_179),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_153),
.A2(n_48),
.B1(n_47),
.B2(n_38),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_168),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_153),
.A2(n_47),
.B1(n_48),
.B2(n_104),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_169),
.A2(n_177),
.B1(n_213),
.B2(n_225),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_103),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_170),
.B(n_173),
.Y(n_267)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_111),
.Y(n_171)
);

INVx11_ASAP7_75t_L g231 ( 
.A(n_171),
.Y(n_231)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_130),
.Y(n_172)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_172),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_93),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_174),
.A2(n_193),
.B1(n_200),
.B2(n_221),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_118),
.B(n_92),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_175),
.B(n_186),
.Y(n_229)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_176),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_161),
.A2(n_85),
.B1(n_73),
.B2(n_72),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_178),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_115),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_180),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_181),
.Y(n_256)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_109),
.Y(n_182)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_182),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_112),
.Y(n_184)
);

INVx11_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

INVx11_ASAP7_75t_L g185 ( 
.A(n_111),
.Y(n_185)
);

BUFx4f_ASAP7_75t_SL g234 ( 
.A(n_185),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_118),
.B(n_74),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_110),
.Y(n_187)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_187),
.Y(n_260)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_188),
.Y(n_245)
);

OR2x2_ASAP7_75t_SL g189 ( 
.A(n_116),
.B(n_74),
.Y(n_189)
);

OR2x2_ASAP7_75t_SL g236 ( 
.A(n_189),
.B(n_209),
.Y(n_236)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_128),
.Y(n_191)
);

INVx13_ASAP7_75t_L g266 ( 
.A(n_191),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_135),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_192),
.B(n_196),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_114),
.A2(n_157),
.B1(n_155),
.B2(n_159),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_116),
.B(n_71),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_194),
.B(n_201),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_134),
.B(n_136),
.Y(n_195)
);

OAI21xp33_ASAP7_75t_L g249 ( 
.A1(n_195),
.A2(n_216),
.B(n_220),
.Y(n_249)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_120),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_124),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_197),
.B(n_199),
.Y(n_253)
);

A2O1A1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_123),
.A2(n_99),
.B(n_2),
.C(n_3),
.Y(n_198)
);

A2O1A1Ixp33_ASAP7_75t_L g273 ( 
.A1(n_198),
.A2(n_217),
.B(n_218),
.C(n_211),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_120),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_160),
.A2(n_139),
.B1(n_137),
.B2(n_143),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_126),
.B(n_1),
.Y(n_201)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_121),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_202),
.B(n_206),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_133),
.B(n_1),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_203),
.B(n_10),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_105),
.A2(n_135),
.B(n_121),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_204),
.A2(n_165),
.B(n_8),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_107),
.B(n_3),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_205),
.B(n_219),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_106),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_161),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_207),
.B(n_208),
.Y(n_261)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_148),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_131),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_211),
.B(n_212),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_119),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_142),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_149),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_214),
.B(n_215),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_154),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_105),
.B(n_4),
.C(n_5),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_217),
.B(n_182),
.C(n_172),
.Y(n_274)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_139),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_113),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_133),
.Y(n_222)
);

BUFx12_ASAP7_75t_L g263 ( 
.A(n_222),
.Y(n_263)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_113),
.Y(n_223)
);

NOR3xp33_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_224),
.C(n_138),
.Y(n_239)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_158),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_112),
.Y(n_225)
);

AND2x2_ASAP7_75t_SL g226 ( 
.A(n_175),
.B(n_158),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_226),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_170),
.B(n_163),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_228),
.B(n_252),
.Y(n_275)
);

O2A1O1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_204),
.A2(n_186),
.B(n_194),
.C(n_210),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_235),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_237),
.A2(n_242),
.B(n_273),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_170),
.A2(n_163),
.B1(n_138),
.B2(n_129),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_238),
.A2(n_251),
.B1(n_226),
.B2(n_267),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_239),
.Y(n_303)
);

OR2x4_ASAP7_75t_L g242 ( 
.A(n_173),
.B(n_7),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_193),
.A2(n_165),
.B1(n_129),
.B2(n_9),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_243),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_174),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_244),
.A2(n_255),
.B1(n_236),
.B2(n_233),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_249),
.Y(n_318)
);

INVx2_ASAP7_75t_R g250 ( 
.A(n_189),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_250),
.A2(n_180),
.B(n_181),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_173),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_200),
.A2(n_10),
.B1(n_13),
.B2(n_210),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_257),
.A2(n_262),
.B1(n_254),
.B2(n_256),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_203),
.B(n_205),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_265),
.Y(n_277)
);

CKINVDCx9p33_ASAP7_75t_R g264 ( 
.A(n_198),
.Y(n_264)
);

INVx8_ASAP7_75t_L g299 ( 
.A(n_264),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_190),
.B(n_201),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_183),
.B(n_187),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_176),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_274),
.B(n_247),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_276),
.A2(n_256),
.B1(n_241),
.B2(n_231),
.Y(n_332)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_253),
.Y(n_278)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_278),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_279),
.B(n_286),
.Y(n_322)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_241),
.Y(n_280)
);

INVx5_ASAP7_75t_L g344 ( 
.A(n_280),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_261),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_281),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_227),
.A2(n_178),
.B1(n_197),
.B2(n_208),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_282),
.A2(n_284),
.B1(n_290),
.B2(n_301),
.Y(n_323)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_230),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g347 ( 
.A(n_283),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_227),
.A2(n_171),
.B1(n_225),
.B2(n_184),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_252),
.B(n_202),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_260),
.Y(n_287)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_287),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_248),
.B(n_196),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_288),
.B(n_309),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_272),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_289),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_226),
.A2(n_264),
.B1(n_267),
.B2(n_237),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_291),
.B(n_316),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_248),
.B(n_206),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_292),
.B(n_308),
.Y(n_355)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_260),
.Y(n_293)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_293),
.Y(n_342)
);

OAI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_259),
.A2(n_185),
.B1(n_250),
.B2(n_236),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_294),
.A2(n_311),
.B1(n_299),
.B2(n_312),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_295),
.A2(n_317),
.B1(n_234),
.B2(n_240),
.Y(n_345)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_232),
.Y(n_296)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_296),
.Y(n_353)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_232),
.Y(n_297)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_297),
.Y(n_356)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_268),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_298),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_226),
.A2(n_267),
.B1(n_238),
.B2(n_228),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_268),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_302),
.Y(n_329)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_230),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_304),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_259),
.A2(n_257),
.B1(n_250),
.B2(n_245),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_305),
.A2(n_313),
.B(n_234),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_235),
.A2(n_255),
.B1(n_251),
.B2(n_270),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g328 ( 
.A1(n_306),
.A2(n_289),
.B1(n_299),
.B2(n_309),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_246),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_308),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_262),
.B(n_229),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_258),
.B(n_229),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_310),
.B(n_319),
.Y(n_339)
);

OAI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_273),
.A2(n_242),
.B1(n_262),
.B2(n_247),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_245),
.A2(n_256),
.B1(n_241),
.B2(n_269),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_230),
.Y(n_314)
);

INVx6_ASAP7_75t_L g330 ( 
.A(n_314),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_315),
.B(n_245),
.C(n_266),
.Y(n_334)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_269),
.Y(n_316)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_271),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_317),
.A2(n_300),
.B(n_291),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_326),
.A2(n_340),
.B(n_351),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_312),
.A2(n_274),
.B1(n_265),
.B2(n_231),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_327),
.A2(n_332),
.B1(n_346),
.B2(n_350),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_328),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_334),
.B(n_336),
.C(n_338),
.Y(n_382)
);

AO21x1_ASAP7_75t_L g378 ( 
.A1(n_335),
.A2(n_359),
.B(n_302),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_315),
.B(n_266),
.C(n_263),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_337),
.B(n_355),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_310),
.B(n_266),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_300),
.A2(n_234),
.B(n_263),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_277),
.B(n_263),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_343),
.B(n_345),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_276),
.A2(n_240),
.B1(n_234),
.B2(n_263),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_285),
.B(n_277),
.C(n_301),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_348),
.B(n_349),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_275),
.B(n_290),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_295),
.A2(n_307),
.B1(n_299),
.B2(n_285),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_278),
.A2(n_281),
.B(n_279),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_275),
.B(n_286),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_352),
.B(n_338),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_284),
.A2(n_282),
.B1(n_303),
.B2(n_319),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_357),
.A2(n_323),
.B1(n_327),
.B2(n_321),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_288),
.A2(n_316),
.B(n_287),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_331),
.B(n_318),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_360),
.B(n_368),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_359),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_361),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_326),
.A2(n_280),
.B(n_293),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_362),
.A2(n_381),
.B(n_388),
.Y(n_400)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_325),
.Y(n_365)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_365),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_351),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_366),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_321),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_331),
.B(n_296),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_369),
.B(n_374),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_354),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_372),
.B(n_376),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_320),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_340),
.A2(n_304),
.B(n_297),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_375),
.A2(n_378),
.B(n_356),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_341),
.B(n_298),
.Y(n_377)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_377),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_341),
.B(n_283),
.Y(n_379)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_379),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_339),
.B(n_314),
.Y(n_380)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_380),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_320),
.A2(n_350),
.B(n_345),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_354),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_383),
.B(n_385),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_339),
.B(n_322),
.Y(n_384)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_384),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_322),
.Y(n_385)
);

AO22x1_ASAP7_75t_L g386 ( 
.A1(n_337),
.A2(n_323),
.B1(n_320),
.B2(n_346),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_386),
.B(n_390),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_387),
.A2(n_363),
.B1(n_386),
.B2(n_364),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_348),
.A2(n_333),
.B(n_334),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_325),
.Y(n_389)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_389),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_333),
.B(n_352),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_342),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_391),
.B(n_392),
.Y(n_418)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_342),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_353),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_393),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_344),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_394),
.B(n_344),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_371),
.A2(n_386),
.B1(n_367),
.B2(n_361),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_395),
.A2(n_396),
.B1(n_406),
.B2(n_420),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_386),
.A2(n_349),
.B1(n_343),
.B2(n_335),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_382),
.B(n_373),
.C(n_336),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_398),
.B(n_408),
.C(n_416),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_373),
.B(n_356),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_399),
.B(n_419),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_403),
.A2(n_363),
.B1(n_381),
.B2(n_378),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_367),
.A2(n_358),
.B1(n_347),
.B2(n_353),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_407),
.A2(n_414),
.B(n_423),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_382),
.B(n_324),
.C(n_329),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_411),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_364),
.A2(n_330),
.B(n_366),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_382),
.B(n_330),
.C(n_388),
.Y(n_416)
);

XNOR2x1_ASAP7_75t_L g419 ( 
.A(n_376),
.B(n_388),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_385),
.A2(n_387),
.B1(n_363),
.B2(n_374),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_390),
.B(n_374),
.C(n_370),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_422),
.B(n_365),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_370),
.A2(n_378),
.B(n_381),
.Y(n_423)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_409),
.Y(n_426)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_426),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_404),
.B(n_369),
.Y(n_427)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_427),
.Y(n_459)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_409),
.Y(n_429)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_429),
.Y(n_461)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_418),
.Y(n_430)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_430),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_421),
.B(n_383),
.Y(n_431)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_431),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_413),
.B(n_377),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_432),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_433),
.A2(n_438),
.B1(n_440),
.B2(n_445),
.Y(n_467)
);

INVxp33_ASAP7_75t_L g434 ( 
.A(n_401),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_434),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_403),
.A2(n_362),
.B1(n_375),
.B2(n_372),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_395),
.A2(n_360),
.B1(n_368),
.B2(n_384),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_439),
.A2(n_441),
.B1(n_443),
.B2(n_448),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_418),
.Y(n_440)
);

INVx13_ASAP7_75t_L g441 ( 
.A(n_411),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_407),
.A2(n_362),
.B(n_379),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_442),
.B(n_444),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_411),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_398),
.B(n_380),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_401),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_446),
.B(n_449),
.Y(n_457)
);

BUFx12_ASAP7_75t_L g448 ( 
.A(n_412),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_421),
.A2(n_389),
.B1(n_391),
.B2(n_392),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_402),
.A2(n_393),
.B1(n_394),
.B2(n_405),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_450),
.A2(n_451),
.B1(n_429),
.B2(n_426),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_424),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_447),
.B(n_416),
.C(n_408),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_453),
.B(n_456),
.C(n_460),
.Y(n_486)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_454),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_447),
.B(n_399),
.C(n_419),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_422),
.C(n_400),
.Y(n_460)
);

FAx1_ASAP7_75t_SL g463 ( 
.A(n_437),
.B(n_417),
.CI(n_396),
.CON(n_463),
.SN(n_463)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_463),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_437),
.B(n_400),
.C(n_414),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_464),
.B(n_472),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_436),
.A2(n_402),
.B1(n_405),
.B2(n_410),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_465),
.A2(n_466),
.B1(n_473),
.B2(n_438),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_436),
.A2(n_410),
.B1(n_415),
.B2(n_420),
.Y(n_466)
);

FAx1_ASAP7_75t_SL g470 ( 
.A(n_432),
.B(n_417),
.CI(n_415),
.CON(n_470),
.SN(n_470)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_470),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_428),
.B(n_423),
.C(n_406),
.Y(n_472)
);

OR2x4_ASAP7_75t_L g473 ( 
.A(n_430),
.B(n_397),
.Y(n_473)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_474),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_452),
.B(n_428),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_475),
.B(n_476),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_464),
.B(n_433),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_469),
.B(n_412),
.Y(n_477)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_477),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_471),
.B(n_451),
.Y(n_479)
);

CKINVDCx14_ASAP7_75t_R g491 ( 
.A(n_479),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_454),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_480),
.B(n_483),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_470),
.B(n_445),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_452),
.B(n_442),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_484),
.B(n_457),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_462),
.B(n_440),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_487),
.B(n_488),
.Y(n_498)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_458),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_467),
.B(n_427),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_489),
.B(n_435),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_SL g490 ( 
.A1(n_459),
.A2(n_443),
.B1(n_435),
.B2(n_425),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_490),
.A2(n_455),
.B1(n_465),
.B2(n_466),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_481),
.A2(n_482),
.B1(n_478),
.B2(n_468),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_492),
.B(n_496),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_486),
.B(n_453),
.C(n_460),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_494),
.B(n_500),
.C(n_450),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_485),
.B(n_472),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_497),
.B(n_502),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_486),
.B(n_476),
.C(n_456),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_501),
.B(n_504),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_475),
.B(n_457),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_484),
.B(n_463),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_505),
.B(n_441),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_499),
.A2(n_482),
.B1(n_461),
.B2(n_489),
.Y(n_506)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_506),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_508),
.B(n_514),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_496),
.A2(n_479),
.B(n_483),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_509),
.A2(n_511),
.B(n_498),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_495),
.A2(n_487),
.B1(n_449),
.B2(n_473),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_510),
.A2(n_491),
.B1(n_503),
.B2(n_505),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_494),
.A2(n_477),
.B(n_425),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_500),
.B(n_397),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_515),
.B(n_516),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_493),
.B(n_448),
.C(n_504),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_517),
.B(n_520),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_508),
.A2(n_493),
.B(n_497),
.Y(n_521)
);

CKINVDCx16_ASAP7_75t_R g527 ( 
.A(n_521),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_513),
.B(n_448),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_523),
.B(n_510),
.Y(n_525)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_525),
.Y(n_529)
);

NOR2x1_ASAP7_75t_L g526 ( 
.A(n_522),
.B(n_506),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_526),
.B(n_516),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_527),
.B(n_519),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_528),
.B(n_529),
.Y(n_532)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_530),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_523),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_531),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_534),
.B(n_524),
.C(n_507),
.Y(n_535)
);

AO21x1_ASAP7_75t_L g536 ( 
.A1(n_535),
.A2(n_526),
.B(n_518),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_536),
.B(n_512),
.C(n_448),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_512),
.Y(n_538)
);


endmodule