module real_aes_17768_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_635;
wire n_287;
wire n_503;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_666;
wire n_320;
wire n_551;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_860;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_898;
wire n_115;
wire n_604;
wire n_110;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_237;
wire n_797;
wire n_862;
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_0), .Y(n_244) );
AND2x4_ASAP7_75t_L g114 ( .A(n_1), .B(n_115), .Y(n_114) );
XNOR2x2_ASAP7_75t_L g899 ( .A(n_2), .B(n_900), .Y(n_899) );
BUFx3_ASAP7_75t_L g185 ( .A(n_3), .Y(n_185) );
INVx1_ASAP7_75t_L g115 ( .A(n_4), .Y(n_115) );
AOI22x1_ASAP7_75t_SL g513 ( .A1(n_5), .A2(n_27), .B1(n_514), .B2(n_515), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_5), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_6), .B(n_157), .Y(n_156) );
BUFx2_ASAP7_75t_L g120 ( .A(n_7), .Y(n_120) );
OR2x2_ASAP7_75t_L g131 ( .A(n_7), .B(n_21), .Y(n_131) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_8), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_9), .B(n_179), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_10), .B(n_179), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_11), .B(n_204), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_12), .A2(n_83), .B1(n_154), .B2(n_179), .Y(n_253) );
OAI21x1_ASAP7_75t_L g149 ( .A1(n_13), .A2(n_37), .B(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_14), .B(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_15), .B(n_194), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g581 ( .A(n_16), .Y(n_581) );
AO32x2_ASAP7_75t_L g250 ( .A1(n_17), .A2(n_171), .A3(n_172), .B1(n_251), .B2(n_254), .Y(n_250) );
AO32x1_ASAP7_75t_L g288 ( .A1(n_17), .A2(n_171), .A3(n_172), .B1(n_251), .B2(n_254), .Y(n_288) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_18), .B(n_566), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_19), .B(n_171), .Y(n_615) );
CKINVDCx5p33_ASAP7_75t_R g594 ( .A(n_20), .Y(n_594) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_21), .Y(n_118) );
AOI22xp33_ASAP7_75t_L g260 ( .A1(n_22), .A2(n_43), .B1(n_182), .B2(n_194), .Y(n_260) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_23), .A2(n_92), .B1(n_154), .B2(n_162), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_24), .B(n_161), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g585 ( .A(n_25), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_26), .B(n_217), .Y(n_277) );
INVx1_ASAP7_75t_L g515 ( .A(n_27), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_28), .A2(n_63), .B1(n_162), .B2(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g636 ( .A(n_29), .B(n_179), .Y(n_636) );
INVx2_ASAP7_75t_L g126 ( .A(n_30), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_31), .B(n_158), .Y(n_667) );
INVx1_ASAP7_75t_L g110 ( .A(n_32), .Y(n_110) );
BUFx3_ASAP7_75t_L g537 ( .A(n_32), .Y(n_537) );
CKINVDCx5p33_ASAP7_75t_R g524 ( .A(n_33), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g896 ( .A1(n_34), .A2(n_56), .B1(n_897), .B2(n_898), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_34), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_35), .B(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_36), .B(n_572), .Y(n_673) );
AND2x2_ASAP7_75t_L g587 ( .A(n_38), .B(n_572), .Y(n_587) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_39), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_40), .B(n_216), .Y(n_609) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_41), .B(n_566), .Y(n_565) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_42), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_44), .B(n_599), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g215 ( .A1(n_45), .A2(n_77), .B1(n_216), .B2(n_217), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_46), .B(n_259), .Y(n_570) );
A2O1A1Ixp33_ASAP7_75t_L g579 ( .A1(n_47), .A2(n_195), .B(n_242), .C(n_580), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g178 ( .A1(n_48), .A2(n_79), .B1(n_154), .B2(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g150 ( .A(n_49), .Y(n_150) );
AND2x4_ASAP7_75t_L g168 ( .A(n_50), .B(n_169), .Y(n_168) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_51), .A2(n_52), .B1(n_162), .B2(n_182), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_53), .B(n_171), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_54), .B(n_572), .Y(n_611) );
CKINVDCx5p33_ASAP7_75t_R g586 ( .A(n_55), .Y(n_586) );
INVxp67_ASAP7_75t_SL g898 ( .A(n_56), .Y(n_898) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_57), .B(n_162), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_58), .B(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g169 ( .A(n_59), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_60), .B(n_171), .Y(n_170) );
A2O1A1Ixp33_ASAP7_75t_L g241 ( .A1(n_61), .A2(n_242), .B(n_243), .C(n_245), .Y(n_241) );
NAND3xp33_ASAP7_75t_L g166 ( .A(n_62), .B(n_154), .C(n_164), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g647 ( .A(n_64), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_65), .B(n_171), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_66), .A2(n_518), .B1(n_519), .B2(n_520), .Y(n_517) );
INVx1_ASAP7_75t_L g519 ( .A(n_66), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_67), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g247 ( .A(n_68), .B(n_248), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_69), .Y(n_263) );
NAND3xp33_ASAP7_75t_L g668 ( .A(n_70), .B(n_158), .C(n_194), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_71), .A2(n_96), .B1(n_179), .B2(n_216), .Y(n_220) );
INVx2_ASAP7_75t_L g159 ( .A(n_72), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_73), .B(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_74), .B(n_564), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_75), .B(n_179), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_76), .B(n_219), .Y(n_606) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_78), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_80), .B(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_81), .B(n_198), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_82), .A2(n_91), .B1(n_566), .B2(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_84), .B(n_179), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_85), .B(n_164), .Y(n_163) );
NAND2xp33_ASAP7_75t_SL g610 ( .A(n_86), .B(n_157), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_87), .A2(n_105), .B1(n_121), .B2(n_903), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_88), .B(n_192), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_89), .A2(n_103), .B1(n_162), .B2(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_90), .B(n_217), .Y(n_274) );
INVx1_ASAP7_75t_SL g900 ( .A(n_93), .Y(n_900) );
INVx1_ASAP7_75t_L g113 ( .A(n_94), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_95), .B(n_204), .Y(n_280) );
NAND2xp33_ASAP7_75t_L g619 ( .A(n_97), .B(n_157), .Y(n_619) );
INVx1_ASAP7_75t_L g518 ( .A(n_98), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_98), .B(n_572), .Y(n_571) );
NAND3xp33_ASAP7_75t_L g607 ( .A(n_99), .B(n_157), .C(n_219), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_100), .B(n_564), .Y(n_638) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_101), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_102), .B(n_566), .Y(n_569) );
CKINVDCx11_ASAP7_75t_R g903 ( .A(n_105), .Y(n_903) );
CKINVDCx11_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
OR2x6_ASAP7_75t_L g106 ( .A(n_107), .B(n_116), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
NOR2x1p5_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
AND3x2_ASAP7_75t_L g129 ( .A(n_109), .B(n_112), .C(n_130), .Y(n_129) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_114), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g535 ( .A(n_113), .Y(n_535) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
NOR2x1p5_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_538), .Y(n_121) );
OAI21xp33_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_127), .B(n_526), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx3_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_126), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g542 ( .A(n_126), .Y(n_542) );
AOI21x1_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_132), .B(n_523), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx4_ASAP7_75t_L g525 ( .A(n_129), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_130), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NOR2x1_ASAP7_75t_L g536 ( .A(n_131), .B(n_537), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_510), .B1(n_511), .B2(n_521), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_135), .Y(n_522) );
INVx2_ASAP7_75t_L g550 ( .A(n_135), .Y(n_550) );
OR2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_420), .Y(n_135) );
NAND4xp25_ASAP7_75t_L g136 ( .A(n_137), .B(n_325), .C(n_352), .D(n_388), .Y(n_136) );
AOI221x1_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_230), .B1(n_264), .B2(n_300), .C(n_304), .Y(n_137) );
NAND3xp33_ASAP7_75t_L g138 ( .A(n_139), .B(n_206), .C(n_228), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_173), .Y(n_141) );
INVx2_ASAP7_75t_L g265 ( .A(n_142), .Y(n_265) );
AND2x2_ASAP7_75t_L g438 ( .A(n_142), .B(n_382), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_142), .B(n_229), .Y(n_447) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g453 ( .A(n_143), .Y(n_453) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g298 ( .A(n_144), .Y(n_298) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OR2x2_ASAP7_75t_L g381 ( .A(n_145), .B(n_227), .Y(n_381) );
OAI21x1_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_151), .B(n_170), .Y(n_145) );
OAI21xp5_ASAP7_75t_L g310 ( .A1(n_146), .A2(n_151), .B(n_170), .Y(n_310) );
OAI21x1_ASAP7_75t_L g560 ( .A1(n_146), .A2(n_561), .B(n_571), .Y(n_560) );
OAI21xp5_ASAP7_75t_L g591 ( .A1(n_146), .A2(n_592), .B(n_600), .Y(n_591) );
OAI21x1_ASAP7_75t_L g690 ( .A1(n_146), .A2(n_592), .B(n_600), .Y(n_690) );
OAI21xp33_ASAP7_75t_SL g781 ( .A1(n_146), .A2(n_561), .B(n_571), .Y(n_781) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g572 ( .A(n_147), .Y(n_572) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g205 ( .A(n_148), .Y(n_205) );
INVx2_ASAP7_75t_L g225 ( .A(n_148), .Y(n_225) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_149), .Y(n_172) );
OAI21x1_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_160), .B(n_167), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_156), .B(n_158), .Y(n_152) );
INVx2_ASAP7_75t_SL g217 ( .A(n_154), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_154), .B(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_155), .Y(n_157) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_155), .Y(n_162) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_155), .Y(n_179) );
INVx1_ASAP7_75t_L g182 ( .A(n_155), .Y(n_182) );
INVx1_ASAP7_75t_L g192 ( .A(n_155), .Y(n_192) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_155), .Y(n_194) );
INVx1_ASAP7_75t_L g216 ( .A(n_155), .Y(n_216) );
INVx1_ASAP7_75t_L g242 ( .A(n_155), .Y(n_242) );
INVx3_ASAP7_75t_L g564 ( .A(n_155), .Y(n_564) );
INVx1_ASAP7_75t_L g567 ( .A(n_155), .Y(n_567) );
INVx2_ASAP7_75t_L g599 ( .A(n_157), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g177 ( .A1(n_158), .A2(n_178), .B1(n_180), .B2(n_181), .Y(n_177) );
INVx6_ASAP7_75t_L g180 ( .A(n_158), .Y(n_180) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_158), .A2(n_195), .B1(n_252), .B2(n_253), .Y(n_251) );
O2A1O1Ixp5_ASAP7_75t_L g593 ( .A1(n_158), .A2(n_191), .B(n_594), .C(n_595), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_158), .A2(n_638), .B(n_639), .Y(n_637) );
BUFx8_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g165 ( .A(n_159), .Y(n_165) );
INVx2_ASAP7_75t_L g200 ( .A(n_159), .Y(n_200) );
INVx1_ASAP7_75t_L g219 ( .A(n_159), .Y(n_219) );
OAI21xp5_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_163), .B(n_166), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
OAI22xp33_ASAP7_75t_L g584 ( .A1(n_162), .A2(n_564), .B1(n_585), .B2(n_586), .Y(n_584) );
INVx2_ASAP7_75t_L g644 ( .A(n_162), .Y(n_644) );
OAI21xp5_ASAP7_75t_L g666 ( .A1(n_162), .A2(n_667), .B(n_668), .Y(n_666) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
BUFx4f_ASAP7_75t_L g195 ( .A(n_165), .Y(n_195) );
AOI31xp67_ASAP7_75t_L g175 ( .A1(n_167), .A2(n_176), .A3(n_177), .B(n_183), .Y(n_175) );
OAI21x1_ASAP7_75t_L g188 ( .A1(n_167), .A2(n_189), .B(n_196), .Y(n_188) );
OAI21x1_ASAP7_75t_L g561 ( .A1(n_167), .A2(n_562), .B(n_568), .Y(n_561) );
OAI21x1_ASAP7_75t_L g592 ( .A1(n_167), .A2(n_593), .B(n_596), .Y(n_592) );
OAI21x1_ASAP7_75t_L g604 ( .A1(n_167), .A2(n_605), .B(n_608), .Y(n_604) );
AND2x4_ASAP7_75t_SL g624 ( .A(n_167), .B(n_172), .Y(n_624) );
OAI21x1_ASAP7_75t_L g633 ( .A1(n_167), .A2(n_634), .B(n_637), .Y(n_633) );
OAI21x1_ASAP7_75t_L g665 ( .A1(n_167), .A2(n_666), .B(n_669), .Y(n_665) );
BUFx10_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g222 ( .A(n_168), .Y(n_222) );
INVx1_ASAP7_75t_L g246 ( .A(n_168), .Y(n_246) );
AO31x2_ASAP7_75t_L g256 ( .A1(n_168), .A2(n_213), .A3(n_257), .B(n_262), .Y(n_256) );
BUFx10_ASAP7_75t_L g577 ( .A(n_168), .Y(n_577) );
INVx2_ASAP7_75t_L g176 ( .A(n_171), .Y(n_176) );
INVx4_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_172), .B(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g187 ( .A(n_172), .Y(n_187) );
BUFx3_ASAP7_75t_L g213 ( .A(n_172), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_172), .B(n_263), .Y(n_262) );
INVx2_ASAP7_75t_SL g271 ( .A(n_172), .Y(n_271) );
INVx1_ASAP7_75t_SL g603 ( .A(n_172), .Y(n_603) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_173), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_173), .B(n_409), .Y(n_408) );
INVxp67_ASAP7_75t_L g451 ( .A(n_173), .Y(n_451) );
AND2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_186), .Y(n_173) );
AND2x2_ASAP7_75t_L g229 ( .A(n_174), .B(n_212), .Y(n_229) );
INVx2_ASAP7_75t_L g307 ( .A(n_174), .Y(n_307) );
AND2x2_ASAP7_75t_L g372 ( .A(n_174), .B(n_310), .Y(n_372) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g227 ( .A(n_175), .Y(n_227) );
INVx3_ASAP7_75t_L g279 ( .A(n_179), .Y(n_279) );
OAI21xp5_ASAP7_75t_L g605 ( .A1(n_179), .A2(n_606), .B(n_607), .Y(n_605) );
INVx1_ASAP7_75t_L g672 ( .A(n_179), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g214 ( .A1(n_180), .A2(n_215), .B1(n_218), .B2(n_220), .Y(n_214) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_180), .A2(n_258), .B1(n_260), .B2(n_261), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_180), .A2(n_277), .B(n_278), .Y(n_276) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_180), .A2(n_583), .B1(n_643), .B2(n_645), .Y(n_642) );
INVx1_ASAP7_75t_L g201 ( .A(n_182), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_182), .A2(n_194), .B1(n_238), .B2(n_239), .Y(n_237) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g299 ( .A(n_186), .Y(n_299) );
AND2x2_ASAP7_75t_L g309 ( .A(n_186), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g371 ( .A(n_186), .B(n_212), .Y(n_371) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_203), .Y(n_186) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_187), .A2(n_188), .B(n_203), .Y(n_209) );
OAI21x1_ASAP7_75t_L g632 ( .A1(n_187), .A2(n_633), .B(n_640), .Y(n_632) );
OAI21x1_ASAP7_75t_L g664 ( .A1(n_187), .A2(n_665), .B(n_673), .Y(n_664) );
OA21x2_ASAP7_75t_L g676 ( .A1(n_187), .A2(n_665), .B(n_673), .Y(n_676) );
OAI21x1_ASAP7_75t_L g679 ( .A1(n_187), .A2(n_633), .B(n_640), .Y(n_679) );
O2A1O1Ixp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_193), .C(n_195), .Y(n_189) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g259 ( .A(n_194), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_195), .A2(n_563), .B(n_565), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_195), .A2(n_609), .B(n_610), .Y(n_608) );
AOI21xp5_ASAP7_75t_L g617 ( .A1(n_195), .A2(n_618), .B(n_619), .Y(n_617) );
AOI21xp5_ASAP7_75t_L g634 ( .A1(n_195), .A2(n_635), .B(n_636), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_199), .B1(n_201), .B2(n_202), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g596 ( .A1(n_198), .A2(n_597), .B(n_598), .Y(n_596) );
INVx2_ASAP7_75t_SL g198 ( .A(n_199), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_199), .A2(n_621), .B1(n_622), .B2(n_623), .Y(n_620) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
BUFx3_ASAP7_75t_L g245 ( .A(n_200), .Y(n_245) );
INVx2_ASAP7_75t_L g234 ( .A(n_204), .Y(n_234) );
NOR2xp67_ASAP7_75t_SL g575 ( .A(n_204), .B(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AO31x2_ASAP7_75t_L g641 ( .A1(n_205), .A2(n_577), .A3(n_642), .B(n_646), .Y(n_641) );
INVx1_ASAP7_75t_L g336 ( .A(n_206), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_207), .B(n_210), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_208), .B(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_208), .B(n_351), .Y(n_350) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_208), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_208), .B(n_406), .Y(n_413) );
INVx2_ASAP7_75t_SL g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g382 ( .A(n_209), .B(n_357), .Y(n_382) );
OR2x2_ASAP7_75t_L g384 ( .A(n_209), .B(n_310), .Y(n_384) );
INVx1_ASAP7_75t_L g443 ( .A(n_209), .Y(n_443) );
BUFx2_ASAP7_75t_L g457 ( .A(n_209), .Y(n_457) );
OR2x2_ASAP7_75t_L g485 ( .A(n_209), .B(n_212), .Y(n_485) );
INVx1_ASAP7_75t_L g504 ( .A(n_210), .Y(n_504) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g351 ( .A(n_211), .Y(n_351) );
OR2x2_ASAP7_75t_L g364 ( .A(n_211), .B(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g383 ( .A(n_211), .B(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_226), .Y(n_211) );
INVx2_ASAP7_75t_L g303 ( .A(n_212), .Y(n_303) );
AND2x2_ASAP7_75t_L g319 ( .A(n_212), .B(n_226), .Y(n_319) );
INVx1_ASAP7_75t_L g357 ( .A(n_212), .Y(n_357) );
INVx1_ASAP7_75t_L g400 ( .A(n_212), .Y(n_400) );
AND2x2_ASAP7_75t_L g442 ( .A(n_212), .B(n_443), .Y(n_442) );
AO31x2_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .A3(n_221), .B(n_223), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_216), .B(n_244), .Y(n_243) );
INVx1_ASAP7_75t_SL g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g240 ( .A(n_219), .Y(n_240) );
INVx2_ASAP7_75t_SL g221 ( .A(n_222), .Y(n_221) );
INVx2_ASAP7_75t_SL g254 ( .A(n_222), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
INVx2_ASAP7_75t_L g248 ( .A(n_225), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_225), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g498 ( .A(n_228), .Y(n_498) );
AND2x4_ASAP7_75t_L g436 ( .A(n_229), .B(n_296), .Y(n_436) );
INVx2_ASAP7_75t_L g465 ( .A(n_229), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_229), .B(n_457), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_230), .B(n_455), .Y(n_454) );
AND2x4_ASAP7_75t_L g230 ( .A(n_231), .B(n_249), .Y(n_230) );
AND2x2_ASAP7_75t_L g376 ( .A(n_231), .B(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g397 ( .A(n_231), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
OR2x2_ASAP7_75t_L g268 ( .A(n_232), .B(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g292 ( .A(n_232), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g323 ( .A(n_232), .Y(n_323) );
AND2x2_ASAP7_75t_L g363 ( .A(n_232), .B(n_255), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_232), .B(n_347), .Y(n_404) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g316 ( .A(n_233), .Y(n_316) );
AOI21x1_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_247), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_241), .B(n_246), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_237), .B(n_240), .Y(n_236) );
AOI21x1_ASAP7_75t_L g669 ( .A1(n_240), .A2(n_670), .B(n_671), .Y(n_669) );
INVx1_ASAP7_75t_L g622 ( .A(n_242), .Y(n_622) );
INVx2_ASAP7_75t_L g261 ( .A(n_245), .Y(n_261) );
INVx2_ASAP7_75t_L g583 ( .A(n_245), .Y(n_583) );
INVx3_ASAP7_75t_L g282 ( .A(n_249), .Y(n_282) );
AND2x2_ASAP7_75t_L g327 ( .A(n_249), .B(n_322), .Y(n_327) );
AND2x2_ASAP7_75t_L g482 ( .A(n_249), .B(n_286), .Y(n_482) );
AND2x4_ASAP7_75t_L g249 ( .A(n_250), .B(n_255), .Y(n_249) );
INVx1_ASAP7_75t_L g333 ( .A(n_250), .Y(n_333) );
AND2x2_ASAP7_75t_L g361 ( .A(n_250), .B(n_269), .Y(n_361) );
OAI21x1_ASAP7_75t_L g272 ( .A1(n_254), .A2(n_273), .B(n_276), .Y(n_272) );
AND2x4_ASAP7_75t_L g314 ( .A(n_255), .B(n_315), .Y(n_314) );
INVx3_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g287 ( .A(n_256), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g324 ( .A(n_256), .B(n_288), .Y(n_324) );
AND2x2_ASAP7_75t_L g334 ( .A(n_256), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_256), .B(n_269), .Y(n_386) );
AND2x2_ASAP7_75t_L g392 ( .A(n_256), .B(n_316), .Y(n_392) );
AOI21x1_ASAP7_75t_L g273 ( .A1(n_261), .A2(n_274), .B(n_275), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_261), .A2(n_569), .B(n_570), .Y(n_568) );
OAI21xp33_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_266), .B(n_283), .Y(n_264) );
OAI21xp33_ASAP7_75t_L g425 ( .A1(n_265), .A2(n_426), .B(n_430), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_265), .B(n_456), .Y(n_503) );
NAND2x1_ASAP7_75t_SL g266 ( .A(n_267), .B(n_281), .Y(n_266) );
INVx1_ASAP7_75t_L g509 ( .A(n_267), .Y(n_509) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
BUFx2_ASAP7_75t_L g286 ( .A(n_269), .Y(n_286) );
INVx2_ASAP7_75t_L g291 ( .A(n_269), .Y(n_291) );
INVxp67_ASAP7_75t_L g312 ( .A(n_269), .Y(n_312) );
AND2x2_ASAP7_75t_L g332 ( .A(n_269), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g343 ( .A(n_269), .B(n_344), .Y(n_343) );
INVx3_ASAP7_75t_L g347 ( .A(n_269), .Y(n_347) );
INVx1_ASAP7_75t_L g365 ( .A(n_269), .Y(n_365) );
OR2x2_ASAP7_75t_L g398 ( .A(n_269), .B(n_333), .Y(n_398) );
INVx1_ASAP7_75t_L g469 ( .A(n_269), .Y(n_469) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OAI21x1_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_272), .B(n_280), .Y(n_270) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OAI21xp33_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_289), .B(n_294), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OAI22xp33_ASAP7_75t_L g407 ( .A1(n_285), .A2(n_408), .B1(n_410), .B2(n_413), .Y(n_407) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_286), .B(n_334), .Y(n_368) );
BUFx2_ASAP7_75t_L g427 ( .A(n_286), .Y(n_427) );
INVx2_ASAP7_75t_L g377 ( .A(n_287), .Y(n_377) );
OR2x2_ASAP7_75t_L g461 ( .A(n_287), .B(n_291), .Y(n_461) );
INVx1_ASAP7_75t_L g293 ( .A(n_288), .Y(n_293) );
INVx1_ASAP7_75t_L g342 ( .A(n_288), .Y(n_342) );
NOR2x1p5_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
INVxp67_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_291), .Y(n_412) );
OR2x2_ASAP7_75t_L g496 ( .A(n_291), .B(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g499 ( .A(n_291), .B(n_334), .Y(n_499) );
INVxp67_ASAP7_75t_SL g462 ( .A(n_292), .Y(n_462) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_296), .B(n_356), .Y(n_418) );
AND2x2_ASAP7_75t_L g508 ( .A(n_296), .B(n_306), .Y(n_508) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g417 ( .A(n_297), .B(n_306), .Y(n_417) );
NAND2x1p5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
AND2x2_ASAP7_75t_L g374 ( .A(n_298), .B(n_307), .Y(n_374) );
AND2x2_ASAP7_75t_L g409 ( .A(n_298), .B(n_303), .Y(n_409) );
INVxp67_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g328 ( .A(n_301), .B(n_309), .Y(n_328) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx2_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g468 ( .A(n_303), .B(n_469), .Y(n_468) );
OAI22xp33_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_311), .B1(n_317), .B2(n_320), .Y(n_304) );
O2A1O1Ixp33_ASAP7_75t_L g505 ( .A1(n_305), .A2(n_506), .B(n_507), .C(n_509), .Y(n_505) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g356 ( .A(n_307), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g424 ( .A(n_307), .Y(n_424) );
OR2x2_ASAP7_75t_L g471 ( .A(n_308), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
AND2x2_ASAP7_75t_L g326 ( .A(n_312), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g429 ( .A(n_315), .Y(n_429) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g335 ( .A(n_316), .Y(n_335) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_316), .Y(n_344) );
INVx1_ASAP7_75t_L g416 ( .A(n_316), .Y(n_416) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g472 ( .A(n_319), .Y(n_472) );
AND2x2_ASAP7_75t_L g494 ( .A(n_319), .B(n_457), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_320), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g346 ( .A(n_324), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g402 ( .A(n_324), .B(n_403), .Y(n_402) );
INVx2_ASAP7_75t_SL g497 ( .A(n_324), .Y(n_497) );
AOI221xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_328), .B1(n_329), .B2(n_336), .C(n_337), .Y(n_325) );
INVxp67_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_334), .Y(n_331) );
INVx2_ASAP7_75t_L g419 ( .A(n_332), .Y(n_419) );
BUFx2_ASAP7_75t_L g439 ( .A(n_334), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_345), .B(n_348), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_340), .B(n_343), .Y(n_339) );
AND2x2_ASAP7_75t_L g481 ( .A(n_340), .B(n_403), .Y(n_481) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g387 ( .A(n_342), .Y(n_387) );
AND2x2_ASAP7_75t_L g477 ( .A(n_342), .B(n_347), .Y(n_477) );
INVx1_ASAP7_75t_L g360 ( .A(n_344), .Y(n_360) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AOI211xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_354), .B(n_366), .C(n_378), .Y(n_352) );
OAI22xp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_358), .B1(n_362), .B2(n_364), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
BUFx2_ASAP7_75t_L g394 ( .A(n_361), .Y(n_394) );
AND2x2_ASAP7_75t_L g487 ( .A(n_361), .B(n_429), .Y(n_487) );
OAI21xp33_ASAP7_75t_L g490 ( .A1(n_362), .A2(n_491), .B(n_493), .Y(n_490) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_369), .B1(n_373), .B2(n_375), .Y(n_366) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_369), .B(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
INVxp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x4_ASAP7_75t_L g441 ( .A(n_374), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x4_ASAP7_75t_L g428 ( .A(n_377), .B(n_429), .Y(n_428) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_377), .Y(n_444) );
AOI21xp33_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_383), .B(n_385), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
AND2x2_ASAP7_75t_L g455 ( .A(n_380), .B(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g492 ( .A(n_380), .B(n_457), .Y(n_492) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g406 ( .A(n_381), .Y(n_406) );
OR2x2_ASAP7_75t_L g484 ( .A(n_381), .B(n_485), .Y(n_484) );
OR2x2_ASAP7_75t_L g399 ( .A(n_384), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g431 ( .A(n_384), .Y(n_431) );
OR2x2_ASAP7_75t_L g464 ( .A(n_384), .B(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g435 ( .A(n_385), .Y(n_435) );
OR2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
NOR3xp33_ASAP7_75t_L g388 ( .A(n_389), .B(n_407), .C(n_414), .Y(n_388) );
OAI322xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_393), .A3(n_395), .B1(n_397), .B2(n_399), .C1(n_401), .C2(n_405), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
A2O1A1Ixp33_ASAP7_75t_L g466 ( .A1(n_391), .A2(n_431), .B(n_467), .C(n_470), .Y(n_466) );
BUFx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g411 ( .A(n_392), .B(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g448 ( .A(n_392), .Y(n_448) );
AND2x4_ASAP7_75t_L g476 ( .A(n_392), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AOI32xp33_ASAP7_75t_L g445 ( .A1(n_394), .A2(n_432), .A3(n_446), .B1(n_448), .B2(n_449), .Y(n_445) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g432 ( .A(n_398), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_400), .B(n_453), .Y(n_452) );
INVxp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
O2A1O1Ixp33_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_417), .B(n_418), .C(n_419), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_421), .B(n_478), .Y(n_420) );
AOI211xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_425), .B(n_433), .C(n_458), .Y(n_421) );
INVxp67_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
O2A1O1Ixp33_ASAP7_75t_SL g500 ( .A1(n_426), .A2(n_501), .B(n_502), .C(n_504), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
OAI31xp33_ASAP7_75t_L g480 ( .A1(n_428), .A2(n_481), .A3(n_482), .B(n_483), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx2_ASAP7_75t_L g440 ( .A(n_432), .Y(n_440) );
NAND4xp25_ASAP7_75t_SL g433 ( .A(n_434), .B(n_437), .C(n_445), .D(n_454), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
AOI32xp33_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_439), .A3(n_440), .B1(n_441), .B2(n_444), .Y(n_437) );
INVx1_ASAP7_75t_L g489 ( .A(n_441), .Y(n_489) );
INVx1_ASAP7_75t_L g501 ( .A(n_444), .Y(n_501) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND3xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_466), .C(n_473), .Y(n_458) );
OAI21xp5_ASAP7_75t_SL g459 ( .A1(n_460), .A2(n_462), .B(n_463), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_467), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_476), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NOR4xp25_ASAP7_75t_L g478 ( .A(n_479), .B(n_490), .C(n_500), .D(n_505), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_486), .Y(n_479) );
OAI21xp33_ASAP7_75t_L g486 ( .A1(n_481), .A2(n_487), .B(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B1(n_498), .B2(n_499), .Y(n_493) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_497), .Y(n_506) );
INVxp67_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
CKINVDCx5p33_ASAP7_75t_R g510 ( .A(n_511), .Y(n_510) );
OAI22xp5_ASAP7_75t_SL g511 ( .A1(n_512), .A2(n_513), .B1(n_516), .B2(n_517), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_518), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_523), .B(n_527), .Y(n_526) );
NOR2x1_ASAP7_75t_R g523 ( .A(n_524), .B(n_525), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx10_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_535), .Y(n_549) );
BUFx8_ASAP7_75t_SL g894 ( .A(n_535), .Y(n_894) );
INVx1_ASAP7_75t_L g544 ( .A(n_537), .Y(n_544) );
NOR2xp67_ASAP7_75t_L g538 ( .A(n_539), .B(n_545), .Y(n_538) );
CKINVDCx5p33_ASAP7_75t_R g539 ( .A(n_540), .Y(n_539) );
BUFx12f_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x6_ASAP7_75t_SL g541 ( .A(n_542), .B(n_543), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_895), .B1(n_901), .B2(n_902), .Y(n_545) );
INVx1_ASAP7_75t_L g901 ( .A(n_546), .Y(n_901) );
OA21x2_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_550), .B(n_551), .Y(n_546) );
INVx8_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
BUFx12f_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_894), .Y(n_551) );
NAND2x1p5_ASAP7_75t_L g552 ( .A(n_553), .B(n_789), .Y(n_552) );
NOR2x1_ASAP7_75t_L g553 ( .A(n_554), .B(n_724), .Y(n_553) );
NAND3xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_648), .C(n_697), .Y(n_554) );
A2O1A1Ixp33_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_588), .B(n_612), .C(n_629), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OR2x2_ASAP7_75t_L g863 ( .A(n_557), .B(n_782), .Y(n_863) );
OR2x2_ASAP7_75t_L g874 ( .A(n_557), .B(n_875), .Y(n_874) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_558), .B(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g765 ( .A(n_558), .B(n_655), .Y(n_765) );
AND2x2_ASAP7_75t_L g886 ( .A(n_558), .B(n_696), .Y(n_886) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_573), .Y(n_558) );
INVx2_ASAP7_75t_L g716 ( .A(n_559), .Y(n_716) );
AND2x2_ASAP7_75t_L g731 ( .A(n_559), .B(n_683), .Y(n_731) );
AND2x2_ASAP7_75t_L g740 ( .A(n_559), .B(n_614), .Y(n_740) );
AND2x2_ASAP7_75t_L g809 ( .A(n_559), .B(n_695), .Y(n_809) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g627 ( .A(n_560), .Y(n_627) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g780 ( .A(n_573), .B(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g628 ( .A(n_574), .B(n_602), .Y(n_628) );
INVx2_ASAP7_75t_L g653 ( .A(n_574), .Y(n_653) );
AOI21x1_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_578), .B(n_587), .Y(n_574) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_582), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
AND2x2_ASAP7_75t_L g817 ( .A(n_588), .B(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_601), .Y(n_589) );
INVx1_ASAP7_75t_L g837 ( .A(n_590), .Y(n_837) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g675 ( .A(n_591), .B(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g758 ( .A(n_591), .B(n_664), .Y(n_758) );
AND2x2_ASAP7_75t_L g684 ( .A(n_601), .B(n_627), .Y(n_684) );
INVxp67_ASAP7_75t_L g833 ( .A(n_601), .Y(n_833) );
OR2x2_ASAP7_75t_L g875 ( .A(n_601), .B(n_614), .Y(n_875) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g657 ( .A(n_602), .Y(n_657) );
OAI21x1_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .B(n_611), .Y(n_602) );
AND2x4_ASAP7_75t_L g612 ( .A(n_613), .B(n_625), .Y(n_612) );
INVx1_ASAP7_75t_L g730 ( .A(n_613), .Y(n_730) );
AND2x2_ASAP7_75t_L g884 ( .A(n_613), .B(n_780), .Y(n_884) );
BUFx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g656 ( .A(n_614), .Y(n_656) );
INVx4_ASAP7_75t_L g695 ( .A(n_614), .Y(n_695) );
AND2x4_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
OAI21x1_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_620), .B(n_624), .Y(n_616) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_628), .Y(n_625) );
AND2x2_ASAP7_75t_L g711 ( .A(n_626), .B(n_694), .Y(n_711) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_L g748 ( .A(n_627), .B(n_696), .Y(n_748) );
INVx2_ASAP7_75t_L g714 ( .A(n_628), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_628), .B(n_719), .Y(n_882) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_631), .B(n_795), .Y(n_794) );
BUFx2_ASAP7_75t_L g867 ( .A(n_631), .Y(n_867) );
AND2x2_ASAP7_75t_L g881 ( .A(n_631), .B(n_703), .Y(n_881) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_641), .Y(n_631) );
INVx1_ASAP7_75t_L g662 ( .A(n_632), .Y(n_662) );
AND2x2_ASAP7_75t_L g816 ( .A(n_632), .B(n_723), .Y(n_816) );
OR2x2_ASAP7_75t_L g853 ( .A(n_632), .B(n_641), .Y(n_853) );
AND2x2_ASAP7_75t_L g663 ( .A(n_641), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g677 ( .A(n_641), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g723 ( .A(n_641), .Y(n_723) );
OR2x2_ASAP7_75t_L g736 ( .A(n_641), .B(n_676), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_641), .B(n_676), .Y(n_769) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_658), .B(n_680), .Y(n_648) );
INVxp67_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AOI31xp33_ASAP7_75t_L g726 ( .A1(n_650), .A2(n_727), .A3(n_729), .B(n_732), .Y(n_726) );
OR2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_654), .Y(n_650) );
AND2x2_ASAP7_75t_L g739 ( .A(n_651), .B(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g749 ( .A(n_652), .Y(n_749) );
HB1xp67_ASAP7_75t_L g755 ( .A(n_652), .Y(n_755) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx2_ASAP7_75t_L g683 ( .A(n_653), .Y(n_683) );
AND2x2_ASAP7_75t_L g712 ( .A(n_653), .B(n_696), .Y(n_712) );
INVx2_ASAP7_75t_L g762 ( .A(n_653), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_654), .B(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g787 ( .A(n_655), .B(n_788), .Y(n_787) );
AND2x2_ASAP7_75t_L g836 ( .A(n_655), .B(n_837), .Y(n_836) );
AOI33xp33_ASAP7_75t_L g891 ( .A1(n_655), .A2(n_721), .A3(n_731), .B1(n_758), .B2(n_867), .B3(n_892), .Y(n_891) );
AND2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
INVx2_ASAP7_75t_L g696 ( .A(n_657), .Y(n_696) );
INVx1_ASAP7_75t_L g783 ( .A(n_657), .Y(n_783) );
INVxp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_660), .B(n_674), .Y(n_659) );
INVx2_ASAP7_75t_L g691 ( .A(n_660), .Y(n_691) );
AND2x2_ASAP7_75t_L g772 ( .A(n_660), .B(n_773), .Y(n_772) );
AND2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_663), .Y(n_660) );
INVx1_ASAP7_75t_L g734 ( .A(n_661), .Y(n_734) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g802 ( .A(n_662), .B(n_689), .Y(n_802) );
AND2x2_ASAP7_75t_L g752 ( .A(n_663), .B(n_746), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_663), .B(n_770), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_663), .B(n_802), .Y(n_851) );
AND2x2_ASAP7_75t_L g688 ( .A(n_664), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g707 ( .A(n_664), .B(n_702), .Y(n_707) );
INVx1_ASAP7_75t_L g722 ( .A(n_664), .Y(n_722) );
AND2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_677), .Y(n_674) );
INVx1_ASAP7_75t_L g777 ( .A(n_675), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_675), .B(n_870), .Y(n_872) );
AND2x2_ASAP7_75t_L g885 ( .A(n_675), .B(n_701), .Y(n_885) );
AND2x2_ASAP7_75t_L g703 ( .A(n_676), .B(n_689), .Y(n_703) );
INVx2_ASAP7_75t_L g685 ( .A(n_677), .Y(n_685) );
AND2x2_ASAP7_75t_L g799 ( .A(n_677), .B(n_800), .Y(n_799) );
AND2x2_ASAP7_75t_L g858 ( .A(n_677), .B(n_770), .Y(n_858) );
BUFx2_ASAP7_75t_L g840 ( .A(n_678), .Y(n_840) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
BUFx3_ASAP7_75t_L g702 ( .A(n_679), .Y(n_702) );
OAI32xp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_685), .A3(n_686), .B1(n_691), .B2(n_692), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
INVx2_ASAP7_75t_L g788 ( .A(n_683), .Y(n_788) );
AND2x2_ASAP7_75t_L g818 ( .A(n_683), .B(n_740), .Y(n_818) );
AND2x2_ASAP7_75t_L g760 ( .A(n_684), .B(n_761), .Y(n_760) );
AND3x2_ASAP7_75t_L g767 ( .A(n_684), .B(n_694), .C(n_762), .Y(n_767) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_687), .A2(n_709), .B1(n_718), .B2(n_720), .Y(n_717) );
OAI322xp33_ASAP7_75t_L g865 ( .A1(n_687), .A2(n_786), .A3(n_866), .B1(n_867), .B2(n_868), .C1(n_869), .C2(n_872), .Y(n_865) );
INVx2_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g887 ( .A(n_688), .B(n_870), .Y(n_887) );
INVxp67_ASAP7_75t_SL g706 ( .A(n_689), .Y(n_706) );
INVxp67_ASAP7_75t_SL g746 ( .A(n_689), .Y(n_746) );
BUFx3_ASAP7_75t_L g770 ( .A(n_689), .Y(n_770) );
INVx1_ASAP7_75t_L g796 ( .A(n_689), .Y(n_796) );
INVx1_ASAP7_75t_L g800 ( .A(n_689), .Y(n_800) );
INVx3_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g754 ( .A(n_693), .B(n_755), .Y(n_754) );
AND2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .Y(n_693) );
INVx1_ASAP7_75t_L g805 ( .A(n_694), .Y(n_805) );
NAND2xp5_ASAP7_75t_SL g856 ( .A(n_694), .B(n_762), .Y(n_856) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
NAND2x1_ASAP7_75t_L g715 ( .A(n_695), .B(n_716), .Y(n_715) );
BUFx2_ASAP7_75t_L g719 ( .A(n_695), .Y(n_719) );
AND2x2_ASAP7_75t_L g761 ( .A(n_695), .B(n_762), .Y(n_761) );
OR2x2_ASAP7_75t_L g782 ( .A(n_695), .B(n_783), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_696), .B(n_809), .Y(n_866) );
O2A1O1Ixp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_704), .B(n_708), .C(n_717), .Y(n_697) );
INVxp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AOI31xp33_ASAP7_75t_L g859 ( .A1(n_699), .A2(n_860), .A3(n_862), .B(n_863), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_700), .B(n_703), .Y(n_699) );
AND2x4_ASAP7_75t_L g812 ( .A(n_700), .B(n_721), .Y(n_812) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_701), .Y(n_744) );
INVx3_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NOR2xp67_ASAP7_75t_L g828 ( .A(n_702), .B(n_722), .Y(n_828) );
BUFx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AND2x4_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
NAND2x1_ASAP7_75t_L g708 ( .A(n_709), .B(n_713), .Y(n_708) );
INVx3_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AND2x4_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
INVx1_ASAP7_75t_L g868 ( .A(n_711), .Y(n_868) );
AND2x2_ASAP7_75t_L g728 ( .A(n_712), .B(n_719), .Y(n_728) );
OAI22xp33_ASAP7_75t_L g797 ( .A1(n_713), .A2(n_798), .B1(n_801), .B2(n_803), .Y(n_797) );
OR2x6_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
INVx1_ASAP7_75t_SL g855 ( .A(n_716), .Y(n_855) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g825 ( .A(n_721), .B(n_770), .Y(n_825) );
INVx2_ASAP7_75t_L g871 ( .A(n_721), .Y(n_871) );
AND2x4_ASAP7_75t_L g879 ( .A(n_721), .B(n_800), .Y(n_879) );
AND2x4_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
NAND3xp33_ASAP7_75t_L g724 ( .A(n_725), .B(n_741), .C(n_771), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_726), .B(n_737), .Y(n_725) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_728), .B(n_858), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
AND2x4_ASAP7_75t_L g792 ( .A(n_730), .B(n_747), .Y(n_792) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_733), .B(n_739), .Y(n_738) );
AND2x4_ASAP7_75t_L g733 ( .A(n_734), .B(n_735), .Y(n_733) );
AND2x2_ASAP7_75t_L g823 ( .A(n_735), .B(n_802), .Y(n_823) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_736), .Y(n_743) );
INVx1_ASAP7_75t_L g861 ( .A(n_736), .Y(n_861) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g890 ( .A(n_739), .Y(n_890) );
HB1xp67_ASAP7_75t_L g775 ( .A(n_740), .Y(n_775) );
AOI211xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_747), .B(n_750), .C(n_763), .Y(n_741) );
NOR3x1_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .C(n_745), .Y(n_742) );
NAND2x1_ASAP7_75t_L g811 ( .A(n_745), .B(n_812), .Y(n_811) );
BUFx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NOR2x1p5_ASAP7_75t_SL g747 ( .A(n_748), .B(n_749), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_753), .B1(n_756), .B2(n_759), .Y(n_750) );
INVxp67_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g844 ( .A(n_755), .Y(n_844) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
BUFx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
AND2x2_ASAP7_75t_L g839 ( .A(n_758), .B(n_840), .Y(n_839) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g893 ( .A(n_761), .Y(n_893) );
AOI21xp33_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_766), .B(n_768), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g847 ( .A(n_768), .Y(n_847) );
OR2x2_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
INVx2_ASAP7_75t_L g774 ( .A(n_770), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_770), .B(n_828), .Y(n_827) );
AOI21xp33_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_775), .B(n_776), .Y(n_771) );
INVxp67_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_774), .B(n_861), .Y(n_860) );
OAI22xp33_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_778), .B1(n_784), .B2(n_786), .Y(n_776) );
OR2x2_ASAP7_75t_L g778 ( .A(n_779), .B(n_782), .Y(n_778) );
INVx1_ASAP7_75t_L g829 ( .A(n_779), .Y(n_829) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
AND2x2_ASAP7_75t_L g804 ( .A(n_780), .B(n_805), .Y(n_804) );
BUFx2_ASAP7_75t_L g821 ( .A(n_781), .Y(n_821) );
INVx1_ASAP7_75t_L g841 ( .A(n_782), .Y(n_841) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
NOR2x1_ASAP7_75t_L g789 ( .A(n_790), .B(n_845), .Y(n_789) );
NAND3xp33_ASAP7_75t_SL g790 ( .A(n_791), .B(n_806), .C(n_819), .Y(n_790) );
AOI21xp5_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_793), .B(n_797), .Y(n_791) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
OR2x2_ASAP7_75t_L g852 ( .A(n_795), .B(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
NAND2x1p5_ASAP7_75t_L g849 ( .A(n_804), .B(n_832), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_810), .B1(n_813), .B2(n_817), .Y(n_806) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx2_ASAP7_75t_L g862 ( .A(n_812), .Y(n_862) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
OAI21xp33_ASAP7_75t_L g834 ( .A1(n_814), .A2(n_835), .B(n_838), .Y(n_834) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
HB1xp67_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_830), .B1(n_834), .B2(n_842), .Y(n_819) );
OAI21xp33_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_822), .B(n_824), .Y(n_820) );
INVxp67_ASAP7_75t_SL g822 ( .A(n_823), .Y(n_822) );
OAI21xp5_ASAP7_75t_L g824 ( .A1(n_825), .A2(n_826), .B(n_829), .Y(n_824) );
INVx1_ASAP7_75t_L g889 ( .A(n_825), .Y(n_889) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g878 ( .A(n_828), .Y(n_878) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
BUFx2_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_839), .B(n_841), .Y(n_838) );
INVx2_ASAP7_75t_L g870 ( .A(n_840), .Y(n_870) );
INVxp67_ASAP7_75t_SL g842 ( .A(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_846), .B(n_864), .Y(n_845) );
AOI211xp5_ASAP7_75t_L g846 ( .A1(n_847), .A2(n_848), .B(n_850), .C(n_859), .Y(n_846) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
A2O1A1Ixp33_ASAP7_75t_L g850 ( .A1(n_851), .A2(n_852), .B(n_854), .C(n_857), .Y(n_850) );
OR2x2_ASAP7_75t_L g854 ( .A(n_855), .B(n_856), .Y(n_854) );
NOR3xp33_ASAP7_75t_L g864 ( .A(n_865), .B(n_873), .C(n_888), .Y(n_864) );
OR2x2_ASAP7_75t_L g869 ( .A(n_870), .B(n_871), .Y(n_869) );
OAI221xp5_ASAP7_75t_L g873 ( .A1(n_874), .A2(n_876), .B1(n_880), .B2(n_882), .C(n_883), .Y(n_873) );
NOR2xp67_ASAP7_75t_L g876 ( .A(n_877), .B(n_879), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx2_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_884), .A2(n_885), .B1(n_886), .B2(n_887), .Y(n_883) );
OAI21xp33_ASAP7_75t_SL g888 ( .A1(n_889), .A2(n_890), .B(n_891), .Y(n_888) );
INVx1_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
CKINVDCx5p33_ASAP7_75t_R g902 ( .A(n_895), .Y(n_902) );
XNOR2x2_ASAP7_75t_L g895 ( .A(n_896), .B(n_899), .Y(n_895) );
endmodule