module fake_jpeg_8684_n_64 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_64);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_64;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_35),
.B1(n_28),
.B2(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_36),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_29),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_3),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_4),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_38),
.Y(n_47)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_33),
.B(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_42),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_43),
.B(n_44),
.Y(n_51)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_5),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_7),
.C(n_9),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_45),
.A2(n_16),
.B1(n_19),
.B2(n_20),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_36),
.B(n_14),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_46),
.A2(n_49),
.B1(n_21),
.B2(n_24),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_48),
.A2(n_26),
.B1(n_22),
.B2(n_23),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_15),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_53),
.Y(n_56)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_55),
.B(n_50),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_47),
.Y(n_59)
);

FAx1_ASAP7_75t_SL g60 ( 
.A(n_59),
.B(n_56),
.CI(n_51),
.CON(n_60),
.SN(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_47),
.B1(n_41),
.B2(n_49),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_62),
.A2(n_60),
.B(n_41),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_53),
.Y(n_64)
);


endmodule