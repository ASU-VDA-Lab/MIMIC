module fake_aes_9330_n_39 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
AOI22xp5_ASAP7_75t_L g11 ( .A1(n_1), .A2(n_8), .B1(n_6), .B2(n_0), .Y(n_11) );
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_4), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_1), .B(n_2), .Y(n_13) );
INVx4_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
CKINVDCx8_ASAP7_75t_R g15 ( .A(n_2), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_8), .Y(n_16) );
AND2x2_ASAP7_75t_SL g17 ( .A(n_14), .B(n_3), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_16), .B(n_3), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_14), .Y(n_19) );
AND2x6_ASAP7_75t_L g20 ( .A(n_13), .B(n_10), .Y(n_20) );
OA21x2_ASAP7_75t_L g21 ( .A1(n_18), .A2(n_11), .B(n_14), .Y(n_21) );
OAI21x1_ASAP7_75t_L g22 ( .A1(n_19), .A2(n_15), .B(n_5), .Y(n_22) );
BUFx6f_ASAP7_75t_L g23 ( .A(n_20), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
OR2x2_ASAP7_75t_L g25 ( .A(n_21), .B(n_18), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
INVx2_ASAP7_75t_L g27 ( .A(n_24), .Y(n_27) );
AOI21xp33_ASAP7_75t_SL g28 ( .A1(n_26), .A2(n_17), .B(n_21), .Y(n_28) );
NOR4xp25_ASAP7_75t_SL g29 ( .A(n_27), .B(n_22), .C(n_12), .D(n_21), .Y(n_29) );
AOI21xp5_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_27), .B(n_23), .Y(n_30) );
NAND2xp33_ASAP7_75t_SL g31 ( .A(n_28), .B(n_12), .Y(n_31) );
AND5x1_ASAP7_75t_L g32 ( .A(n_28), .B(n_21), .C(n_20), .D(n_6), .E(n_7), .Y(n_32) );
NAND2xp5_ASAP7_75t_L g33 ( .A(n_31), .B(n_20), .Y(n_33) );
OAI22xp5_ASAP7_75t_SL g34 ( .A1(n_32), .A2(n_4), .B1(n_5), .B2(n_7), .Y(n_34) );
NOR2x1_ASAP7_75t_L g35 ( .A(n_30), .B(n_23), .Y(n_35) );
NAND2xp5_ASAP7_75t_L g36 ( .A(n_34), .B(n_9), .Y(n_36) );
NAND2x1_ASAP7_75t_L g37 ( .A(n_35), .B(n_23), .Y(n_37) );
AO22x2_ASAP7_75t_L g38 ( .A1(n_36), .A2(n_33), .B1(n_9), .B2(n_23), .Y(n_38) );
OAI221xp5_ASAP7_75t_R g39 ( .A1(n_38), .A2(n_23), .B1(n_37), .B2(n_11), .C(n_12), .Y(n_39) );
endmodule