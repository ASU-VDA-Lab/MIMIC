module fake_netlist_5_1747_n_1104 (n_137, n_210, n_168, n_260, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_248, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_237, n_90, n_241, n_127, n_75, n_101, n_180, n_184, n_226, n_235, n_65, n_78, n_74, n_144, n_207, n_240, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_229, n_108, n_231, n_257, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_236, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_249, n_46, n_233, n_21, n_94, n_203, n_245, n_205, n_113, n_38, n_123, n_139, n_105, n_246, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_234, n_17, n_92, n_19, n_149, n_120, n_232, n_135, n_30, n_156, n_5, n_33, n_126, n_254, n_14, n_225, n_84, n_23, n_202, n_130, n_219, n_157, n_258, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_244, n_251, n_25, n_53, n_160, n_198, n_223, n_247, n_188, n_190, n_8, n_201, n_158, n_263, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_243, n_239, n_175, n_252, n_169, n_59, n_262, n_26, n_255, n_133, n_238, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_242, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_259, n_222, n_230, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_253, n_261, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_256, n_48, n_204, n_50, n_250, n_52, n_88, n_110, n_216, n_1104);

input n_137;
input n_210;
input n_168;
input n_260;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_237;
input n_90;
input n_241;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_235;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_240;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_229;
input n_108;
input n_231;
input n_257;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_236;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_249;
input n_46;
input n_233;
input n_21;
input n_94;
input n_203;
input n_245;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_246;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_234;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_232;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_254;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_258;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_244;
input n_251;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_247;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_243;
input n_239;
input n_175;
input n_252;
input n_169;
input n_59;
input n_262;
input n_26;
input n_255;
input n_133;
input n_238;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_242;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_259;
input n_222;
input n_230;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_253;
input n_261;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_256;
input n_48;
input n_204;
input n_50;
input n_250;
input n_52;
input n_88;
input n_110;
input n_216;

output n_1104;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_419;
wire n_380;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_316;
wire n_785;
wire n_389;
wire n_855;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_912;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_605;
wire n_776;
wire n_928;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_823;
wire n_983;
wire n_725;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_719;
wire n_372;
wire n_293;
wire n_443;
wire n_677;
wire n_864;
wire n_859;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_946;
wire n_417;
wire n_1048;
wire n_932;
wire n_612;
wire n_1001;
wire n_385;
wire n_498;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_509;
wire n_568;
wire n_936;
wire n_373;
wire n_820;
wire n_757;
wire n_947;
wire n_1090;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_1063;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_394;
wire n_579;
wire n_992;
wire n_1049;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_406;
wire n_519;
wire n_470;
wire n_919;
wire n_782;
wire n_908;
wire n_325;
wire n_449;
wire n_1073;
wire n_1100;
wire n_862;
wire n_1016;
wire n_724;
wire n_856;
wire n_546;
wire n_900;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_942;
wire n_381;
wire n_291;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_976;
wire n_1095;
wire n_1096;
wire n_343;
wire n_428;
wire n_308;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_853;
wire n_603;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_660;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_1062;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_680;
wire n_974;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_342;
wire n_482;
wire n_517;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_1075;
wire n_1069;
wire n_388;
wire n_761;
wire n_1012;
wire n_1019;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_1031;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1015;
wire n_1000;
wire n_891;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_332;
wire n_1053;
wire n_1101;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_289;
wire n_745;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_767;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_1059;
wire n_1084;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_425;
wire n_513;
wire n_679;
wire n_407;
wire n_527;
wire n_710;
wire n_707;
wire n_795;
wire n_857;
wire n_695;
wire n_832;
wire n_1072;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_1027;
wire n_971;
wire n_490;
wire n_805;
wire n_910;
wire n_326;
wire n_794;
wire n_768;
wire n_996;
wire n_921;
wire n_404;
wire n_686;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_596;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_1080;
wire n_266;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_352;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_803;
wire n_868;
wire n_1092;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_817;
wire n_1032;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

INVx1_ASAP7_75t_L g264 ( 
.A(n_252),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_17),
.Y(n_265)
);

BUFx10_ASAP7_75t_L g266 ( 
.A(n_77),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_115),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_211),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_144),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_185),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_155),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_238),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_205),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_50),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_214),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_123),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_170),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_253),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_163),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_112),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_53),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_126),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_104),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_213),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_227),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_93),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_132),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_183),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_26),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_156),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_219),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_122),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_145),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_129),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_47),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_233),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_16),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_14),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_188),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_140),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_173),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_45),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_105),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_235),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_102),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_48),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_160),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_192),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_52),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_203),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_106),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_216),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_150),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_177),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_9),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_199),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_40),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_29),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_197),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_98),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_76),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_41),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_92),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_25),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_256),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_247),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_157),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_287),
.B(n_0),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_268),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_270),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_315),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_274),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_324),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_287),
.B(n_277),
.Y(n_334)
);

NOR2xp67_ASAP7_75t_L g335 ( 
.A(n_289),
.B(n_0),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_265),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_271),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_294),
.B(n_1),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_297),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_311),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_311),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_278),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_298),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_280),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_290),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_264),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_267),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_275),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_276),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_279),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_282),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_269),
.B(n_1),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_318),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_281),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_299),
.Y(n_355)
);

INVxp33_ASAP7_75t_SL g356 ( 
.A(n_283),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_300),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_302),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_327),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_303),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_284),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_305),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_285),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_306),
.B(n_307),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_314),
.Y(n_365)
);

BUFx6f_ASAP7_75t_SL g366 ( 
.A(n_266),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_316),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_320),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_271),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_266),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_347),
.B(n_341),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_346),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_348),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_337),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_349),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_350),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_337),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_354),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_355),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_336),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_336),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_369),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_366),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_357),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_369),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_334),
.B(n_271),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_358),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_366),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_360),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_362),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_328),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_365),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_367),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_341),
.B(n_313),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_368),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_356),
.B(n_326),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_331),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_352),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_333),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_340),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_329),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_330),
.B(n_325),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_364),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_335),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_338),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_332),
.Y(n_406)
);

INVx4_ASAP7_75t_L g407 ( 
.A(n_342),
.Y(n_407)
);

NAND2x1_ASAP7_75t_L g408 ( 
.A(n_344),
.B(n_271),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_351),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_359),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_361),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_363),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_339),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_339),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_343),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_343),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_353),
.B(n_323),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_345),
.Y(n_418)
);

AND2x6_ASAP7_75t_L g419 ( 
.A(n_370),
.B(n_272),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_371),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_371),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_371),
.B(n_370),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_391),
.B(n_272),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_410),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_377),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_377),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_377),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_406),
.B(n_353),
.Y(n_428)
);

OR2x6_ASAP7_75t_L g429 ( 
.A(n_418),
.B(n_272),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_405),
.B(n_286),
.Y(n_430)
);

INVx6_ASAP7_75t_L g431 ( 
.A(n_391),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_416),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_377),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_391),
.B(n_398),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_401),
.B(n_288),
.Y(n_435)
);

INVx5_ASAP7_75t_L g436 ( 
.A(n_377),
.Y(n_436)
);

INVx6_ASAP7_75t_L g437 ( 
.A(n_391),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_385),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_394),
.B(n_291),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_419),
.B(n_396),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_385),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_401),
.B(n_292),
.Y(n_442)
);

INVx4_ASAP7_75t_SL g443 ( 
.A(n_419),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_399),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_418),
.Y(n_445)
);

INVx5_ASAP7_75t_L g446 ( 
.A(n_385),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_391),
.B(n_272),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_385),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_372),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_417),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_373),
.Y(n_451)
);

NOR3xp33_ASAP7_75t_L g452 ( 
.A(n_386),
.B(n_295),
.C(n_293),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_406),
.B(n_359),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_402),
.B(n_322),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_403),
.B(n_296),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_385),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_374),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_393),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_374),
.Y(n_459)
);

BUFx8_ASAP7_75t_SL g460 ( 
.A(n_416),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_398),
.B(n_273),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_394),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_375),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_394),
.B(n_301),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_382),
.Y(n_465)
);

BUFx10_ASAP7_75t_L g466 ( 
.A(n_409),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_376),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_382),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_378),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_403),
.B(n_308),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_393),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_379),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_393),
.Y(n_473)
);

OAI22xp33_ASAP7_75t_L g474 ( 
.A1(n_404),
.A2(n_321),
.B1(n_310),
.B2(n_312),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_400),
.B(n_309),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_384),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_387),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_398),
.B(n_273),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_390),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_395),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_401),
.B(n_319),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_407),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_393),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_386),
.A2(n_317),
.B1(n_304),
.B2(n_273),
.Y(n_484)
);

INVx5_ASAP7_75t_L g485 ( 
.A(n_398),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_455),
.B(n_412),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_428),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_457),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_434),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_424),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_454),
.B(n_398),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_434),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g493 ( 
.A(n_475),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_444),
.Y(n_494)
);

AO22x2_ASAP7_75t_L g495 ( 
.A1(n_484),
.A2(n_414),
.B1(n_415),
.B2(n_413),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_449),
.Y(n_496)
);

NAND3xp33_ASAP7_75t_SL g497 ( 
.A(n_424),
.B(n_414),
.C(n_381),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_460),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_432),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_432),
.B(n_418),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_470),
.B(n_420),
.Y(n_501)
);

AO22x2_ASAP7_75t_L g502 ( 
.A1(n_484),
.A2(n_411),
.B1(n_407),
.B2(n_412),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_451),
.Y(n_503)
);

OAI221xp5_ASAP7_75t_L g504 ( 
.A1(n_452),
.A2(n_400),
.B1(n_392),
.B2(n_397),
.C(n_389),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_422),
.Y(n_505)
);

AO22x2_ASAP7_75t_L g506 ( 
.A1(n_450),
.A2(n_407),
.B1(n_412),
.B2(n_388),
.Y(n_506)
);

AO22x2_ASAP7_75t_L g507 ( 
.A1(n_452),
.A2(n_383),
.B1(n_408),
.B2(n_419),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_421),
.B(n_416),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_463),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_467),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_469),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_459),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_472),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_482),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_465),
.Y(n_515)
);

OAI221xp5_ASAP7_75t_L g516 ( 
.A1(n_440),
.A2(n_392),
.B1(n_397),
.B2(n_389),
.C(n_408),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_476),
.Y(n_517)
);

BUFx8_ASAP7_75t_L g518 ( 
.A(n_445),
.Y(n_518)
);

AO22x2_ASAP7_75t_L g519 ( 
.A1(n_430),
.A2(n_419),
.B1(n_4),
.B2(n_2),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_468),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_466),
.Y(n_521)
);

NAND2x1p5_ASAP7_75t_L g522 ( 
.A(n_462),
.B(n_389),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_453),
.Y(n_523)
);

AO22x2_ASAP7_75t_L g524 ( 
.A1(n_439),
.A2(n_419),
.B1(n_4),
.B2(n_2),
.Y(n_524)
);

NAND2x1p5_ASAP7_75t_L g525 ( 
.A(n_485),
.B(n_477),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_479),
.Y(n_526)
);

OAI221xp5_ASAP7_75t_L g527 ( 
.A1(n_440),
.A2(n_393),
.B1(n_304),
.B2(n_273),
.C(n_416),
.Y(n_527)
);

AO22x2_ASAP7_75t_L g528 ( 
.A1(n_439),
.A2(n_419),
.B1(n_6),
.B2(n_3),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_480),
.Y(n_529)
);

NAND2x1p5_ASAP7_75t_L g530 ( 
.A(n_485),
.B(n_416),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_431),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_431),
.Y(n_532)
);

AO22x2_ASAP7_75t_L g533 ( 
.A1(n_464),
.A2(n_6),
.B1(n_3),
.B2(n_5),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_475),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_431),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_466),
.Y(n_536)
);

AO22x2_ASAP7_75t_L g537 ( 
.A1(n_464),
.A2(n_8),
.B1(n_5),
.B2(n_7),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_437),
.A2(n_304),
.B1(n_380),
.B2(n_9),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_437),
.Y(n_539)
);

NAND2x1p5_ASAP7_75t_L g540 ( 
.A(n_485),
.B(n_304),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_429),
.Y(n_541)
);

AND2x2_ASAP7_75t_SL g542 ( 
.A(n_461),
.B(n_7),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_437),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_429),
.B(n_36),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_423),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_429),
.B(n_37),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_423),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_435),
.B(n_8),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_447),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_447),
.Y(n_550)
);

OR2x6_ASAP7_75t_L g551 ( 
.A(n_442),
.B(n_10),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_461),
.Y(n_552)
);

AO22x2_ASAP7_75t_L g553 ( 
.A1(n_481),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_553)
);

AO22x2_ASAP7_75t_L g554 ( 
.A1(n_443),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_485),
.B(n_38),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_478),
.B(n_13),
.Y(n_556)
);

AO22x2_ASAP7_75t_L g557 ( 
.A1(n_443),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_478),
.B(n_39),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_471),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_486),
.B(n_487),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_523),
.B(n_474),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_501),
.B(n_474),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_514),
.B(n_493),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_508),
.B(n_443),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_534),
.B(n_483),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_500),
.B(n_473),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_489),
.B(n_458),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_499),
.B(n_544),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_494),
.B(n_496),
.Y(n_569)
);

NAND2xp33_ASAP7_75t_SL g570 ( 
.A(n_521),
.B(n_473),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_544),
.B(n_473),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_546),
.B(n_458),
.Y(n_572)
);

NAND2xp33_ASAP7_75t_SL g573 ( 
.A(n_536),
.B(n_548),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_SL g574 ( 
.A(n_538),
.B(n_425),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_546),
.B(n_426),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_491),
.B(n_490),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_503),
.B(n_426),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_509),
.B(n_426),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_510),
.B(n_433),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_511),
.B(n_427),
.Y(n_580)
);

NAND2xp33_ASAP7_75t_SL g581 ( 
.A(n_556),
.B(n_427),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_513),
.B(n_427),
.Y(n_582)
);

NAND2xp33_ASAP7_75t_SL g583 ( 
.A(n_498),
.B(n_441),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_517),
.B(n_441),
.Y(n_584)
);

NAND2xp33_ASAP7_75t_SL g585 ( 
.A(n_526),
.B(n_441),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_489),
.B(n_438),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_492),
.B(n_438),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_529),
.B(n_448),
.Y(n_588)
);

NAND2xp33_ASAP7_75t_SL g589 ( 
.A(n_545),
.B(n_448),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_505),
.B(n_456),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_547),
.B(n_456),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_542),
.B(n_436),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_530),
.B(n_436),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_522),
.B(n_436),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_541),
.B(n_436),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_488),
.B(n_446),
.Y(n_596)
);

NAND2xp33_ASAP7_75t_SL g597 ( 
.A(n_549),
.B(n_15),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_SL g598 ( 
.A(n_550),
.B(n_17),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_512),
.B(n_446),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_515),
.B(n_446),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_520),
.B(n_446),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_552),
.B(n_42),
.Y(n_602)
);

NAND2xp33_ASAP7_75t_SL g603 ( 
.A(n_558),
.B(n_18),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_SL g604 ( 
.A(n_531),
.B(n_18),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_539),
.B(n_532),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_535),
.B(n_543),
.Y(n_606)
);

NAND2xp33_ASAP7_75t_SL g607 ( 
.A(n_555),
.B(n_19),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_518),
.B(n_43),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_518),
.B(n_44),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_525),
.B(n_46),
.Y(n_610)
);

NAND2xp33_ASAP7_75t_SL g611 ( 
.A(n_506),
.B(n_19),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_SL g612 ( 
.A(n_506),
.B(n_20),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_551),
.B(n_49),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_502),
.B(n_20),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_559),
.B(n_51),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_540),
.B(n_54),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_524),
.B(n_528),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_524),
.B(n_55),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_528),
.B(n_56),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_502),
.B(n_57),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_551),
.B(n_21),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_507),
.B(n_58),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_507),
.B(n_59),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_569),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_569),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_562),
.B(n_495),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_568),
.Y(n_627)
);

NAND2xp33_ASAP7_75t_L g628 ( 
.A(n_561),
.B(n_519),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_613),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_SL g630 ( 
.A(n_613),
.B(n_497),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_575),
.A2(n_516),
.B(n_527),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_560),
.A2(n_495),
.B1(n_504),
.B2(n_519),
.Y(n_632)
);

BUFx10_ASAP7_75t_L g633 ( 
.A(n_565),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_571),
.A2(n_557),
.B(n_554),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_576),
.B(n_553),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_565),
.B(n_553),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_572),
.A2(n_557),
.B(n_554),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_579),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_579),
.B(n_533),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_567),
.B(n_533),
.Y(n_640)
);

NAND2x1_ASAP7_75t_L g641 ( 
.A(n_586),
.B(n_537),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_563),
.B(n_21),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_587),
.B(n_537),
.Y(n_643)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_590),
.B(n_583),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_621),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_591),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_588),
.Y(n_647)
);

O2A1O1Ixp5_ASAP7_75t_L g648 ( 
.A1(n_620),
.A2(n_159),
.B(n_262),
.C(n_261),
.Y(n_648)
);

OR2x2_ASAP7_75t_L g649 ( 
.A(n_573),
.B(n_22),
.Y(n_649)
);

INVxp67_ASAP7_75t_L g650 ( 
.A(n_614),
.Y(n_650)
);

INVx4_ASAP7_75t_L g651 ( 
.A(n_570),
.Y(n_651)
);

NAND3xp33_ASAP7_75t_L g652 ( 
.A(n_597),
.B(n_22),
.C(n_23),
.Y(n_652)
);

BUFx5_ASAP7_75t_L g653 ( 
.A(n_564),
.Y(n_653)
);

OAI21xp33_ASAP7_75t_L g654 ( 
.A1(n_592),
.A2(n_23),
.B(n_24),
.Y(n_654)
);

OAI21x1_ASAP7_75t_L g655 ( 
.A1(n_566),
.A2(n_61),
.B(n_60),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_605),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_618),
.B(n_24),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_619),
.B(n_25),
.Y(n_658)
);

AO31x2_ASAP7_75t_L g659 ( 
.A1(n_611),
.A2(n_26),
.A3(n_27),
.B(n_28),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_606),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_617),
.B(n_27),
.Y(n_661)
);

OAI21x1_ASAP7_75t_L g662 ( 
.A1(n_577),
.A2(n_63),
.B(n_62),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_595),
.Y(n_663)
);

OAI21xp5_ASAP7_75t_SL g664 ( 
.A1(n_608),
.A2(n_28),
.B(n_29),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_622),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_574),
.B(n_30),
.Y(n_666)
);

OAI21x1_ASAP7_75t_L g667 ( 
.A1(n_578),
.A2(n_65),
.B(n_64),
.Y(n_667)
);

NAND2xp33_ASAP7_75t_R g668 ( 
.A(n_623),
.B(n_66),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_580),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g670 ( 
.A1(n_602),
.A2(n_68),
.B(n_67),
.Y(n_670)
);

OAI21x1_ASAP7_75t_L g671 ( 
.A1(n_582),
.A2(n_584),
.B(n_596),
.Y(n_671)
);

AO22x2_ASAP7_75t_L g672 ( 
.A1(n_609),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_612),
.B(n_31),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_599),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_604),
.Y(n_675)
);

AO22x2_ASAP7_75t_L g676 ( 
.A1(n_598),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_610),
.B(n_33),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_594),
.B(n_34),
.Y(n_678)
);

NAND3xp33_ASAP7_75t_L g679 ( 
.A(n_603),
.B(n_35),
.C(n_69),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_607),
.Y(n_680)
);

OAI21x1_ASAP7_75t_L g681 ( 
.A1(n_600),
.A2(n_71),
.B(n_70),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_601),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_615),
.Y(n_683)
);

BUFx4f_ASAP7_75t_L g684 ( 
.A(n_585),
.Y(n_684)
);

OAI21x1_ASAP7_75t_L g685 ( 
.A1(n_655),
.A2(n_593),
.B(n_616),
.Y(n_685)
);

AOI21xp33_ASAP7_75t_SL g686 ( 
.A1(n_629),
.A2(n_642),
.B(n_672),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_638),
.Y(n_687)
);

OAI21x1_ASAP7_75t_L g688 ( 
.A1(n_671),
.A2(n_589),
.B(n_581),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_624),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_625),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_650),
.B(n_35),
.Y(n_691)
);

OAI21x1_ASAP7_75t_L g692 ( 
.A1(n_662),
.A2(n_72),
.B(n_73),
.Y(n_692)
);

OAI21x1_ASAP7_75t_L g693 ( 
.A1(n_667),
.A2(n_681),
.B(n_631),
.Y(n_693)
);

NAND2x1p5_ASAP7_75t_L g694 ( 
.A(n_651),
.B(n_74),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_630),
.A2(n_75),
.B1(n_78),
.B2(n_79),
.Y(n_695)
);

NOR2xp67_ASAP7_75t_L g696 ( 
.A(n_627),
.B(n_80),
.Y(n_696)
);

NAND2x1p5_ASAP7_75t_L g697 ( 
.A(n_675),
.B(n_81),
.Y(n_697)
);

AO21x2_ASAP7_75t_L g698 ( 
.A1(n_666),
.A2(n_626),
.B(n_632),
.Y(n_698)
);

OAI21x1_ASAP7_75t_L g699 ( 
.A1(n_648),
.A2(n_82),
.B(n_83),
.Y(n_699)
);

BUFx12f_ASAP7_75t_L g700 ( 
.A(n_633),
.Y(n_700)
);

OAI21x1_ASAP7_75t_L g701 ( 
.A1(n_670),
.A2(n_84),
.B(n_85),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_656),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_645),
.Y(n_703)
);

OAI21xp5_ASAP7_75t_L g704 ( 
.A1(n_628),
.A2(n_86),
.B(n_87),
.Y(n_704)
);

OAI21x1_ASAP7_75t_L g705 ( 
.A1(n_646),
.A2(n_683),
.B(n_647),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_653),
.Y(n_706)
);

AO21x1_ASAP7_75t_L g707 ( 
.A1(n_634),
.A2(n_88),
.B(n_89),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_633),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_663),
.B(n_90),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_680),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_639),
.B(n_91),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_SL g712 ( 
.A1(n_641),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_660),
.Y(n_713)
);

O2A1O1Ixp33_ASAP7_75t_L g714 ( 
.A1(n_673),
.A2(n_97),
.B(n_99),
.C(n_100),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_653),
.Y(n_715)
);

O2A1O1Ixp33_ASAP7_75t_L g716 ( 
.A1(n_643),
.A2(n_101),
.B(n_103),
.C(n_107),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_652),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_717)
);

INVx4_ASAP7_75t_L g718 ( 
.A(n_665),
.Y(n_718)
);

BUFx2_ASAP7_75t_L g719 ( 
.A(n_661),
.Y(n_719)
);

OAI21x1_ASAP7_75t_L g720 ( 
.A1(n_637),
.A2(n_111),
.B(n_113),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_676),
.A2(n_114),
.B1(n_116),
.B2(n_117),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_640),
.B(n_118),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_668),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_SL g724 ( 
.A1(n_672),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_636),
.B(n_124),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_684),
.A2(n_125),
.B(n_127),
.Y(n_726)
);

OAI21x1_ASAP7_75t_L g727 ( 
.A1(n_669),
.A2(n_128),
.B(n_130),
.Y(n_727)
);

A2O1A1Ixp33_ASAP7_75t_L g728 ( 
.A1(n_657),
.A2(n_131),
.B(n_133),
.C(n_134),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_674),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_665),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_L g731 ( 
.A1(n_635),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_676),
.A2(n_654),
.B1(n_679),
.B2(n_658),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_644),
.B(n_138),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_677),
.A2(n_139),
.B(n_141),
.Y(n_734)
);

OAI21x1_ASAP7_75t_L g735 ( 
.A1(n_682),
.A2(n_142),
.B(n_143),
.Y(n_735)
);

OR2x2_ASAP7_75t_L g736 ( 
.A(n_678),
.B(n_649),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_665),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_737)
);

AOI22x1_ASAP7_75t_L g738 ( 
.A1(n_653),
.A2(n_149),
.B1(n_151),
.B2(n_152),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_659),
.Y(n_739)
);

OAI21x1_ASAP7_75t_L g740 ( 
.A1(n_653),
.A2(n_153),
.B(n_154),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_706),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_739),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_702),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_713),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_698),
.B(n_659),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_698),
.B(n_659),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_704),
.A2(n_664),
.B(n_161),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_729),
.Y(n_748)
);

HB1xp67_ASAP7_75t_L g749 ( 
.A(n_710),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_705),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_715),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_720),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_719),
.B(n_158),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_688),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_735),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_727),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_722),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_730),
.Y(n_758)
);

OAI21x1_ASAP7_75t_L g759 ( 
.A1(n_693),
.A2(n_162),
.B(n_164),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_722),
.Y(n_760)
);

BUFx12f_ASAP7_75t_L g761 ( 
.A(n_700),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_707),
.Y(n_762)
);

OAI21x1_ASAP7_75t_L g763 ( 
.A1(n_692),
.A2(n_165),
.B(n_166),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_689),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_687),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_690),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_699),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_740),
.Y(n_768)
);

OAI21x1_ASAP7_75t_L g769 ( 
.A1(n_685),
.A2(n_167),
.B(n_168),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_SL g770 ( 
.A1(n_723),
.A2(n_169),
.B1(n_171),
.B2(n_172),
.Y(n_770)
);

OAI21x1_ASAP7_75t_L g771 ( 
.A1(n_701),
.A2(n_174),
.B(n_175),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_733),
.A2(n_176),
.B1(n_178),
.B2(n_179),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_738),
.Y(n_773)
);

OAI21x1_ASAP7_75t_L g774 ( 
.A1(n_704),
.A2(n_180),
.B(n_181),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_725),
.B(n_263),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_718),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_718),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_697),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_697),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_736),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_731),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_731),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_709),
.Y(n_783)
);

AO21x2_ASAP7_75t_L g784 ( 
.A1(n_686),
.A2(n_182),
.B(n_184),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_696),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_732),
.B(n_186),
.Y(n_786)
);

BUFx2_ASAP7_75t_L g787 ( 
.A(n_708),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_708),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_709),
.Y(n_789)
);

AO21x1_ASAP7_75t_L g790 ( 
.A1(n_716),
.A2(n_187),
.B(n_189),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_703),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_733),
.B(n_260),
.Y(n_792)
);

INVx1_ASAP7_75t_SL g793 ( 
.A(n_711),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_691),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_694),
.Y(n_795)
);

OAI21xp5_ASAP7_75t_L g796 ( 
.A1(n_732),
.A2(n_190),
.B(n_191),
.Y(n_796)
);

AO32x2_ASAP7_75t_L g797 ( 
.A1(n_712),
.A2(n_193),
.A3(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_797)
);

OAI21x1_ASAP7_75t_SL g798 ( 
.A1(n_734),
.A2(n_198),
.B(n_200),
.Y(n_798)
);

AND2x4_ASAP7_75t_L g799 ( 
.A(n_726),
.B(n_201),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_694),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_724),
.B(n_259),
.Y(n_801)
);

INVx1_ASAP7_75t_SL g802 ( 
.A(n_691),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_724),
.A2(n_202),
.B1(n_204),
.B2(n_206),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_717),
.B(n_258),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_780),
.B(n_721),
.Y(n_805)
);

BUFx4f_ASAP7_75t_L g806 ( 
.A(n_758),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_R g807 ( 
.A(n_761),
.B(n_737),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_743),
.Y(n_808)
);

XNOR2xp5_ASAP7_75t_L g809 ( 
.A(n_749),
.B(n_695),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_780),
.B(n_721),
.Y(n_810)
);

NAND2xp33_ASAP7_75t_R g811 ( 
.A(n_799),
.B(n_726),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_758),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_793),
.B(n_737),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_794),
.B(n_734),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_802),
.B(n_717),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_757),
.B(n_716),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_783),
.B(n_789),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_R g818 ( 
.A(n_761),
.B(n_207),
.Y(n_818)
);

INVxp67_ASAP7_75t_L g819 ( 
.A(n_791),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_758),
.B(n_728),
.Y(n_820)
);

INVxp67_ASAP7_75t_L g821 ( 
.A(n_791),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_758),
.Y(n_822)
);

BUFx10_ASAP7_75t_L g823 ( 
.A(n_758),
.Y(n_823)
);

NAND2xp33_ASAP7_75t_R g824 ( 
.A(n_799),
.B(n_208),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_743),
.Y(n_825)
);

NAND2xp33_ASAP7_75t_R g826 ( 
.A(n_799),
.B(n_209),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_R g827 ( 
.A(n_788),
.B(n_785),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_R g828 ( 
.A(n_788),
.B(n_210),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_787),
.Y(n_829)
);

OR2x2_ASAP7_75t_L g830 ( 
.A(n_757),
.B(n_760),
.Y(n_830)
);

INVxp67_ASAP7_75t_L g831 ( 
.A(n_787),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_R g832 ( 
.A(n_775),
.B(n_212),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_783),
.B(n_789),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_R g834 ( 
.A(n_775),
.B(n_215),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_778),
.B(n_217),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_R g836 ( 
.A(n_792),
.B(n_218),
.Y(n_836)
);

NAND2xp33_ASAP7_75t_R g837 ( 
.A(n_801),
.B(n_220),
.Y(n_837)
);

CKINVDCx20_ASAP7_75t_R g838 ( 
.A(n_753),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_742),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_776),
.B(n_221),
.Y(n_840)
);

OR2x6_ASAP7_75t_L g841 ( 
.A(n_795),
.B(n_714),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_760),
.B(n_714),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_776),
.Y(n_843)
);

NAND2xp33_ASAP7_75t_R g844 ( 
.A(n_801),
.B(n_222),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_777),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_R g846 ( 
.A(n_741),
.B(n_781),
.Y(n_846)
);

NAND2xp33_ASAP7_75t_R g847 ( 
.A(n_786),
.B(n_223),
.Y(n_847)
);

BUFx10_ASAP7_75t_L g848 ( 
.A(n_748),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_744),
.B(n_224),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_744),
.Y(n_850)
);

HB1xp67_ASAP7_75t_L g851 ( 
.A(n_766),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_765),
.B(n_766),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_R g853 ( 
.A(n_741),
.B(n_257),
.Y(n_853)
);

INVxp67_ASAP7_75t_L g854 ( 
.A(n_765),
.Y(n_854)
);

OR2x6_ASAP7_75t_L g855 ( 
.A(n_795),
.B(n_225),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_R g856 ( 
.A(n_741),
.B(n_255),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_778),
.B(n_779),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_779),
.B(n_226),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_777),
.B(n_228),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_764),
.B(n_229),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_R g861 ( 
.A(n_781),
.B(n_254),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_850),
.B(n_764),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_SL g863 ( 
.A1(n_855),
.A2(n_796),
.B(n_747),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_839),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_808),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_814),
.B(n_782),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_851),
.B(n_745),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_831),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_825),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_809),
.A2(n_803),
.B1(n_786),
.B2(n_772),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_805),
.B(n_745),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_830),
.Y(n_872)
);

BUFx2_ASAP7_75t_L g873 ( 
.A(n_827),
.Y(n_873)
);

OR2x2_ASAP7_75t_L g874 ( 
.A(n_842),
.B(n_746),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_852),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_816),
.B(n_746),
.Y(n_876)
);

INVxp67_ASAP7_75t_SL g877 ( 
.A(n_854),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_857),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_810),
.B(n_742),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_845),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_857),
.Y(n_881)
);

HB1xp67_ASAP7_75t_L g882 ( 
.A(n_846),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_817),
.B(n_833),
.Y(n_883)
);

OR2x2_ASAP7_75t_L g884 ( 
.A(n_829),
.B(n_754),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_817),
.Y(n_885)
);

AND2x4_ASAP7_75t_SL g886 ( 
.A(n_848),
.B(n_800),
.Y(n_886)
);

INVx5_ASAP7_75t_L g887 ( 
.A(n_841),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_813),
.B(n_782),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_841),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_837),
.A2(n_804),
.B1(n_790),
.B2(n_800),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_812),
.B(n_750),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_815),
.B(n_754),
.Y(n_892)
);

INVxp67_ASAP7_75t_SL g893 ( 
.A(n_811),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_843),
.B(n_751),
.Y(n_894)
);

OR2x2_ASAP7_75t_L g895 ( 
.A(n_819),
.B(n_750),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_822),
.B(n_768),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_843),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_821),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_860),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_849),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_835),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_820),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_838),
.B(n_751),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_823),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_835),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_858),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_858),
.B(n_797),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_806),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_859),
.Y(n_909)
);

INVx2_ASAP7_75t_SL g910 ( 
.A(n_840),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_855),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_824),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_861),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_832),
.B(n_797),
.Y(n_914)
);

NAND2x1p5_ASAP7_75t_SL g915 ( 
.A(n_847),
.B(n_773),
.Y(n_915)
);

OR2x2_ASAP7_75t_L g916 ( 
.A(n_826),
.B(n_762),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_853),
.Y(n_917)
);

OAI22xp5_ASAP7_75t_L g918 ( 
.A1(n_870),
.A2(n_770),
.B1(n_762),
.B2(n_844),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_871),
.B(n_797),
.Y(n_919)
);

INVxp67_ASAP7_75t_SL g920 ( 
.A(n_892),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_871),
.B(n_797),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_889),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_877),
.B(n_784),
.Y(n_923)
);

INVx4_ASAP7_75t_L g924 ( 
.A(n_887),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_865),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_890),
.A2(n_790),
.B1(n_784),
.B2(n_774),
.Y(n_926)
);

OAI221xp5_ASAP7_75t_L g927 ( 
.A1(n_863),
.A2(n_768),
.B1(n_807),
.B2(n_773),
.C(n_755),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_864),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_867),
.B(n_797),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_909),
.B(n_784),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_867),
.B(n_767),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_879),
.B(n_767),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_912),
.A2(n_836),
.B1(n_798),
.B2(n_834),
.Y(n_933)
);

INVx1_ASAP7_75t_SL g934 ( 
.A(n_873),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_879),
.B(n_752),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_865),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_869),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_874),
.B(n_752),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_872),
.Y(n_939)
);

OAI31xp33_ASAP7_75t_L g940 ( 
.A1(n_916),
.A2(n_912),
.A3(n_913),
.B(n_914),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_869),
.Y(n_941)
);

AOI221xp5_ASAP7_75t_L g942 ( 
.A1(n_915),
.A2(n_818),
.B1(n_798),
.B2(n_828),
.C(n_856),
.Y(n_942)
);

INVx4_ASAP7_75t_L g943 ( 
.A(n_887),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_874),
.B(n_756),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_875),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_880),
.Y(n_946)
);

AOI221xp5_ASAP7_75t_L g947 ( 
.A1(n_915),
.A2(n_756),
.B1(n_755),
.B2(n_774),
.C(n_234),
.Y(n_947)
);

INVxp67_ASAP7_75t_SL g948 ( 
.A(n_892),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_895),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_876),
.B(n_769),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_876),
.B(n_769),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_875),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_907),
.B(n_759),
.Y(n_953)
);

OAI33xp33_ASAP7_75t_L g954 ( 
.A1(n_888),
.A2(n_230),
.A3(n_231),
.B1(n_232),
.B2(n_236),
.B3(n_237),
.Y(n_954)
);

INVx2_ASAP7_75t_SL g955 ( 
.A(n_886),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_866),
.B(n_771),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_925),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_920),
.B(n_948),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_928),
.Y(n_959)
);

OR2x2_ASAP7_75t_L g960 ( 
.A(n_949),
.B(n_889),
.Y(n_960)
);

OR2x2_ASAP7_75t_L g961 ( 
.A(n_944),
.B(n_868),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_936),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_936),
.Y(n_963)
);

OR2x2_ASAP7_75t_L g964 ( 
.A(n_944),
.B(n_878),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_925),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_937),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_922),
.B(n_893),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_937),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_922),
.B(n_885),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_938),
.B(n_895),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_953),
.B(n_885),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_955),
.Y(n_972)
);

OR2x6_ASAP7_75t_L g973 ( 
.A(n_924),
.B(n_863),
.Y(n_973)
);

OR2x2_ASAP7_75t_L g974 ( 
.A(n_953),
.B(n_878),
.Y(n_974)
);

AND2x4_ASAP7_75t_SL g975 ( 
.A(n_924),
.B(n_882),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_938),
.B(n_881),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_934),
.B(n_885),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_945),
.B(n_862),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_931),
.B(n_881),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_941),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_939),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_927),
.B(n_916),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_929),
.B(n_907),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_945),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_952),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_952),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_935),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_982),
.A2(n_918),
.B1(n_942),
.B2(n_926),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_982),
.B(n_940),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_961),
.B(n_930),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_970),
.B(n_950),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_970),
.B(n_950),
.Y(n_992)
);

AO221x2_ASAP7_75t_L g993 ( 
.A1(n_981),
.A2(n_903),
.B1(n_911),
.B2(n_917),
.C(n_923),
.Y(n_993)
);

NOR2x1_ASAP7_75t_L g994 ( 
.A(n_972),
.B(n_943),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_960),
.B(n_946),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_967),
.B(n_951),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_959),
.B(n_978),
.Y(n_997)
);

OAI221xp5_ASAP7_75t_L g998 ( 
.A1(n_973),
.A2(n_933),
.B1(n_947),
.B2(n_902),
.C(n_955),
.Y(n_998)
);

AO221x2_ASAP7_75t_L g999 ( 
.A1(n_978),
.A2(n_904),
.B1(n_897),
.B2(n_905),
.C(n_956),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_975),
.Y(n_1000)
);

A2O1A1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_975),
.A2(n_914),
.B(n_887),
.C(n_919),
.Y(n_1001)
);

OAI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_973),
.A2(n_887),
.B1(n_943),
.B2(n_924),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_958),
.B(n_951),
.Y(n_1003)
);

BUFx12f_ASAP7_75t_L g1004 ( 
.A(n_1000),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_994),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_997),
.Y(n_1006)
);

NAND2x1_ASAP7_75t_SL g1007 ( 
.A(n_988),
.B(n_987),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_1003),
.Y(n_1008)
);

OR2x2_ASAP7_75t_L g1009 ( 
.A(n_990),
.B(n_976),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_999),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_991),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_993),
.Y(n_1012)
);

INVx1_ASAP7_75t_SL g1013 ( 
.A(n_989),
.Y(n_1013)
);

INVx1_ASAP7_75t_SL g1014 ( 
.A(n_996),
.Y(n_1014)
);

OR2x2_ASAP7_75t_L g1015 ( 
.A(n_992),
.B(n_964),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_1001),
.B(n_973),
.Y(n_1016)
);

INVx1_ASAP7_75t_SL g1017 ( 
.A(n_1004),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_1013),
.B(n_995),
.Y(n_1018)
);

INVx1_ASAP7_75t_SL g1019 ( 
.A(n_1007),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_1012),
.B(n_987),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1006),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1008),
.Y(n_1022)
);

AOI21xp33_ASAP7_75t_L g1023 ( 
.A1(n_1013),
.A2(n_1002),
.B(n_998),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_1012),
.B(n_971),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_1017),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_1018),
.B(n_1010),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1021),
.Y(n_1027)
);

OR2x2_ASAP7_75t_L g1028 ( 
.A(n_1022),
.B(n_1014),
.Y(n_1028)
);

INVx1_ASAP7_75t_SL g1029 ( 
.A(n_1019),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1020),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_1025),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1030),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1028),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_1027),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1029),
.Y(n_1035)
);

BUFx4f_ASAP7_75t_SL g1036 ( 
.A(n_1029),
.Y(n_1036)
);

OAI211xp5_ASAP7_75t_SL g1037 ( 
.A1(n_1035),
.A2(n_1026),
.B(n_1023),
.C(n_1005),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_1033),
.A2(n_1020),
.B(n_1024),
.Y(n_1038)
);

NAND3xp33_ASAP7_75t_L g1039 ( 
.A(n_1031),
.B(n_1024),
.C(n_1016),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_1036),
.Y(n_1040)
);

NOR3xp33_ASAP7_75t_L g1041 ( 
.A(n_1032),
.B(n_1016),
.C(n_954),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_1034),
.B(n_1014),
.Y(n_1042)
);

NOR4xp25_ASAP7_75t_L g1043 ( 
.A(n_1034),
.B(n_1011),
.C(n_1009),
.D(n_980),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_SL g1044 ( 
.A1(n_1034),
.A2(n_898),
.B(n_886),
.Y(n_1044)
);

AOI222xp33_ASAP7_75t_L g1045 ( 
.A1(n_1042),
.A2(n_887),
.B1(n_880),
.B2(n_921),
.C1(n_919),
.C2(n_929),
.Y(n_1045)
);

AOI211xp5_ASAP7_75t_L g1046 ( 
.A1(n_1037),
.A2(n_977),
.B(n_1015),
.C(n_897),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_1040),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_1039),
.A2(n_943),
.B1(n_966),
.B2(n_968),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_1041),
.A2(n_899),
.B1(n_896),
.B2(n_910),
.Y(n_1049)
);

NAND3xp33_ASAP7_75t_L g1050 ( 
.A(n_1038),
.B(n_899),
.C(n_894),
.Y(n_1050)
);

XOR2xp5_ASAP7_75t_L g1051 ( 
.A(n_1047),
.B(n_1044),
.Y(n_1051)
);

INVxp67_ASAP7_75t_SL g1052 ( 
.A(n_1048),
.Y(n_1052)
);

XNOR2xp5_ASAP7_75t_L g1053 ( 
.A(n_1049),
.B(n_1043),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_1050),
.B(n_962),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_1046),
.B(n_983),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_1045),
.A2(n_900),
.B(n_963),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1049),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_1052),
.B(n_1053),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_R g1059 ( 
.A(n_1057),
.B(n_239),
.Y(n_1059)
);

NAND2xp33_ASAP7_75t_SL g1060 ( 
.A(n_1055),
.B(n_1051),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1054),
.B(n_957),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_1056),
.B(n_969),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_1051),
.B(n_986),
.Y(n_1063)
);

XNOR2x2_ASAP7_75t_L g1064 ( 
.A(n_1053),
.B(n_759),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_R g1065 ( 
.A(n_1053),
.B(n_240),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_R g1066 ( 
.A(n_1053),
.B(n_241),
.Y(n_1066)
);

NAND2xp33_ASAP7_75t_SL g1067 ( 
.A(n_1053),
.B(n_908),
.Y(n_1067)
);

OAI22x1_ASAP7_75t_L g1068 ( 
.A1(n_1058),
.A2(n_1063),
.B1(n_1062),
.B2(n_1061),
.Y(n_1068)
);

OA22x2_ASAP7_75t_L g1069 ( 
.A1(n_1064),
.A2(n_984),
.B1(n_957),
.B2(n_965),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_1059),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_1060),
.Y(n_1071)
);

NAND3x1_ASAP7_75t_L g1072 ( 
.A(n_1065),
.B(n_908),
.C(n_965),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_1067),
.Y(n_1073)
);

NOR2x1p5_ASAP7_75t_L g1074 ( 
.A(n_1066),
.B(n_908),
.Y(n_1074)
);

NOR3xp33_ASAP7_75t_L g1075 ( 
.A(n_1060),
.B(n_900),
.C(n_771),
.Y(n_1075)
);

NAND3xp33_ASAP7_75t_L g1076 ( 
.A(n_1060),
.B(n_985),
.C(n_896),
.Y(n_1076)
);

XNOR2xp5_ASAP7_75t_L g1077 ( 
.A(n_1058),
.B(n_910),
.Y(n_1077)
);

XNOR2x1_ASAP7_75t_L g1078 ( 
.A(n_1058),
.B(n_242),
.Y(n_1078)
);

OAI22x1_ASAP7_75t_L g1079 ( 
.A1(n_1058),
.A2(n_985),
.B1(n_971),
.B2(n_983),
.Y(n_1079)
);

NAND4xp75_ASAP7_75t_L g1080 ( 
.A(n_1058),
.B(n_921),
.C(n_935),
.D(n_931),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1070),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_1074),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_1071),
.B(n_979),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1068),
.Y(n_1084)
);

INVxp67_ASAP7_75t_SL g1085 ( 
.A(n_1072),
.Y(n_1085)
);

INVx3_ASAP7_75t_L g1086 ( 
.A(n_1073),
.Y(n_1086)
);

NOR2x1p5_ASAP7_75t_L g1087 ( 
.A(n_1076),
.B(n_906),
.Y(n_1087)
);

INVxp67_ASAP7_75t_SL g1088 ( 
.A(n_1078),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1086),
.B(n_1077),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_1084),
.A2(n_1075),
.B1(n_1079),
.B2(n_1069),
.Y(n_1090)
);

AOI211x1_ASAP7_75t_L g1091 ( 
.A1(n_1081),
.A2(n_1080),
.B(n_932),
.C(n_883),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1083),
.B(n_974),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1085),
.A2(n_763),
.B(n_896),
.Y(n_1093)
);

AOI31xp33_ASAP7_75t_L g1094 ( 
.A1(n_1089),
.A2(n_1088),
.A3(n_1082),
.B(n_1086),
.Y(n_1094)
);

AOI31xp33_ASAP7_75t_L g1095 ( 
.A1(n_1090),
.A2(n_1087),
.A3(n_906),
.B(n_901),
.Y(n_1095)
);

AOI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_1092),
.A2(n_891),
.B1(n_932),
.B2(n_884),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_1093),
.A2(n_891),
.B1(n_884),
.B2(n_901),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_1094),
.A2(n_1091),
.B(n_244),
.C(n_245),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_1098),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_SL g1100 ( 
.A1(n_1098),
.A2(n_1095),
.B1(n_1097),
.B2(n_1096),
.Y(n_1100)
);

OR2x6_ASAP7_75t_L g1101 ( 
.A(n_1099),
.B(n_763),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1100),
.Y(n_1102)
);

OAI221xp5_ASAP7_75t_R g1103 ( 
.A1(n_1102),
.A2(n_243),
.B1(n_246),
.B2(n_248),
.C(n_249),
.Y(n_1103)
);

AOI211xp5_ASAP7_75t_L g1104 ( 
.A1(n_1103),
.A2(n_1101),
.B(n_250),
.C(n_251),
.Y(n_1104)
);


endmodule