module fake_jpeg_5370_n_265 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_182;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx5_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVxp33_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_30),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_57),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

BUFx4f_ASAP7_75t_SL g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_42),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_48),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_45),
.B(n_60),
.Y(n_76)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_51),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_55),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_58),
.A2(n_21),
.B1(n_22),
.B2(n_28),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_18),
.B(n_1),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_18),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_29),
.B(n_2),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_58),
.A2(n_21),
.B1(n_35),
.B2(n_25),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_63),
.A2(n_88),
.B1(n_101),
.B2(n_32),
.Y(n_118)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_74),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_71),
.A2(n_98),
.B1(n_27),
.B2(n_24),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_38),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_91),
.Y(n_113)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_40),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_80),
.Y(n_106)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_86),
.Y(n_105)
);

CKINVDCx6p67_ASAP7_75t_R g85 ( 
.A(n_55),
.Y(n_85)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_42),
.A2(n_26),
.B(n_3),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_87),
.A2(n_100),
.B(n_37),
.C(n_19),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_46),
.A2(n_22),
.B1(n_21),
.B2(n_35),
.Y(n_88)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_92),
.Y(n_119)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

CKINVDCx12_ASAP7_75t_R g93 ( 
.A(n_42),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_97),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_44),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_94),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_95),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_38),
.Y(n_96)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_57),
.A2(n_22),
.B1(n_25),
.B2(n_31),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_56),
.A2(n_33),
.B1(n_31),
.B2(n_36),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_61),
.A2(n_33),
.B1(n_36),
.B2(n_30),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_102),
.A2(n_110),
.B1(n_112),
.B2(n_129),
.Y(n_137)
);

AND2x2_ASAP7_75t_SL g104 ( 
.A(n_64),
.B(n_47),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_104),
.A2(n_73),
.B(n_66),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_109),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_41),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_108),
.B(n_114),
.Y(n_140)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_78),
.A2(n_20),
.B1(n_24),
.B2(n_27),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_64),
.B(n_32),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_116),
.Y(n_144)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_121),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_118),
.A2(n_117),
.B1(n_132),
.B2(n_114),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_70),
.B(n_49),
.C(n_19),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_87),
.C(n_71),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_75),
.B(n_2),
.Y(n_125)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_127),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_77),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_128),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_79),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_65),
.B(n_3),
.Y(n_130)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_98),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_133),
.B(n_141),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_136),
.C(n_157),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_76),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_63),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_88),
.B1(n_101),
.B2(n_99),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_143),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_95),
.Y(n_145)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_147),
.A2(n_161),
.B(n_131),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_95),
.Y(n_148)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_111),
.B(n_90),
.Y(n_149)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_149),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_89),
.Y(n_150)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_5),
.Y(n_151)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_106),
.B(n_5),
.Y(n_152)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_104),
.A2(n_67),
.B1(n_84),
.B2(n_62),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_104),
.A2(n_108),
.B1(n_106),
.B2(n_120),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_110),
.A2(n_84),
.B1(n_62),
.B2(n_12),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_11),
.C(n_14),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_105),
.B(n_7),
.Y(n_158)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_159),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_16),
.C(n_8),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_115),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_162),
.B(n_168),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_165),
.Y(n_191)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_169),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_144),
.Y(n_168)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_173),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_171),
.A2(n_174),
.B(n_145),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_131),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_141),
.A2(n_103),
.B(n_122),
.Y(n_174)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_181),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_179),
.Y(n_203)
);

CKINVDCx10_ASAP7_75t_R g181 ( 
.A(n_154),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_126),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_142),
.B(n_116),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_184),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_188),
.A2(n_196),
.B1(n_202),
.B2(n_175),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_148),
.C(n_133),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_193),
.Y(n_217)
);

AOI32xp33_ASAP7_75t_L g192 ( 
.A1(n_181),
.A2(n_153),
.A3(n_135),
.B1(n_147),
.B2(n_136),
.Y(n_192)
);

NOR3xp33_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_175),
.C(n_172),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_150),
.C(n_155),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_143),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_171),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_174),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_204),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_185),
.A2(n_137),
.B1(n_151),
.B2(n_152),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_142),
.Y(n_200)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_200),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_201),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_167),
.A2(n_109),
.B1(n_124),
.B2(n_138),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_138),
.Y(n_205)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_186),
.Y(n_207)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_208),
.B(n_214),
.Y(n_230)
);

INVxp33_ASAP7_75t_L g209 ( 
.A(n_197),
.Y(n_209)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_192),
.Y(n_233)
);

NOR3xp33_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_218),
.C(n_177),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_178),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_215),
.A2(n_221),
.B1(n_172),
.B2(n_206),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_198),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_187),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_165),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_219),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_173),
.Y(n_221)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_223),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_190),
.C(n_193),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_231),
.C(n_233),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_229),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_216),
.A2(n_203),
.B1(n_196),
.B2(n_180),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_227),
.A2(n_228),
.B1(n_221),
.B2(n_211),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_218),
.A2(n_179),
.B1(n_204),
.B2(n_200),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_188),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_217),
.C(n_220),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_234),
.C(n_166),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_208),
.Y(n_238)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_238),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_242),
.Y(n_246)
);

MAJx2_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_221),
.C(n_191),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_209),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_223),
.B(n_222),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_199),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_213),
.C(n_164),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_231),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_247),
.C(n_248),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_226),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_250),
.C(n_236),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_235),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_251),
.A2(n_252),
.B(n_183),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_246),
.A2(n_240),
.B(n_241),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_249),
.A2(n_234),
.B1(n_250),
.B2(n_191),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_255),
.C(n_182),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_256),
.A2(n_259),
.B1(n_119),
.B2(n_170),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_258),
.Y(n_260)
);

MAJx2_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_225),
.C(n_157),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_161),
.C(n_158),
.Y(n_259)
);

AOI322xp5_ASAP7_75t_L g262 ( 
.A1(n_261),
.A2(n_126),
.A3(n_128),
.B1(n_16),
.B2(n_107),
.C1(n_9),
.C2(n_7),
.Y(n_262)
);

NOR3xp33_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_263),
.C(n_7),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_260),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_8),
.Y(n_265)
);


endmodule