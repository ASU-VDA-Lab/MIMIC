module real_aes_7680_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_725;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_754;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_762;
wire n_210;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g112 ( .A(n_0), .Y(n_112) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_1), .A2(n_145), .B(n_149), .C(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g198 ( .A(n_2), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_3), .A2(n_140), .B(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_4), .B(n_162), .Y(n_479) );
AOI21xp33_ASAP7_75t_L g166 ( .A1(n_5), .A2(n_140), .B(n_167), .Y(n_166) );
AND2x6_ASAP7_75t_L g145 ( .A(n_6), .B(n_146), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_7), .A2(n_248), .B(n_249), .Y(n_247) );
INVx1_ASAP7_75t_L g110 ( .A(n_8), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_8), .B(n_41), .Y(n_737) );
INVx1_ASAP7_75t_L g535 ( .A(n_9), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_10), .B(n_171), .Y(n_514) );
INVx1_ASAP7_75t_L g173 ( .A(n_11), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_12), .B(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g138 ( .A(n_13), .Y(n_138) );
INVx1_ASAP7_75t_L g254 ( .A(n_14), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_15), .A2(n_157), .B(n_255), .C(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_16), .B(n_162), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_17), .B(n_154), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_18), .B(n_140), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_19), .B(n_563), .Y(n_562) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_20), .A2(n_181), .B(n_240), .C(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_21), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_22), .B(n_171), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_23), .A2(n_252), .B(n_253), .C(n_255), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_24), .B(n_171), .Y(n_486) );
CKINVDCx16_ASAP7_75t_R g459 ( .A(n_25), .Y(n_459) );
INVx1_ASAP7_75t_L g485 ( .A(n_26), .Y(n_485) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_27), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_28), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_29), .B(n_171), .Y(n_200) );
INVx1_ASAP7_75t_L g560 ( .A(n_30), .Y(n_560) );
INVx1_ASAP7_75t_L g187 ( .A(n_31), .Y(n_187) );
OAI22xp5_ASAP7_75t_SL g753 ( .A1(n_32), .A2(n_92), .B1(n_754), .B2(n_755), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_32), .Y(n_755) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_33), .A2(n_105), .B1(n_116), .B2(n_766), .Y(n_104) );
INVx2_ASAP7_75t_L g143 ( .A(n_34), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_35), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g476 ( .A1(n_36), .A2(n_158), .B(n_240), .C(n_477), .Y(n_476) );
INVxp67_ASAP7_75t_L g561 ( .A(n_37), .Y(n_561) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_38), .A2(n_145), .B(n_149), .C(n_212), .Y(n_211) );
CKINVDCx14_ASAP7_75t_R g475 ( .A(n_39), .Y(n_475) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_40), .A2(n_149), .B(n_484), .C(n_489), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_41), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g185 ( .A(n_42), .Y(n_185) );
OAI22xp5_ASAP7_75t_SL g749 ( .A1(n_43), .A2(n_50), .B1(n_750), .B2(n_751), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_43), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g731 ( .A1(n_44), .A2(n_64), .B1(n_732), .B2(n_733), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_44), .Y(n_733) );
OAI22xp5_ASAP7_75t_SL g729 ( .A1(n_45), .A2(n_730), .B1(n_731), .B2(n_734), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_45), .Y(n_734) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_46), .A2(n_170), .B(n_216), .C(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_47), .B(n_171), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_48), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_49), .Y(n_557) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_50), .Y(n_750) );
INVx1_ASAP7_75t_L g500 ( .A(n_51), .Y(n_500) );
CKINVDCx16_ASAP7_75t_R g188 ( .A(n_52), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_53), .B(n_140), .Y(n_242) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_54), .A2(n_149), .B1(n_181), .B2(n_183), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_55), .Y(n_220) );
CKINVDCx16_ASAP7_75t_R g195 ( .A(n_56), .Y(n_195) );
A2O1A1Ixp33_ASAP7_75t_L g169 ( .A1(n_57), .A2(n_158), .B(n_170), .C(n_172), .Y(n_169) );
CKINVDCx14_ASAP7_75t_R g532 ( .A(n_58), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_59), .Y(n_230) );
INVx1_ASAP7_75t_L g168 ( .A(n_60), .Y(n_168) );
INVx1_ASAP7_75t_L g146 ( .A(n_61), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_62), .Y(n_741) );
INVx1_ASAP7_75t_L g137 ( .A(n_63), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_64), .Y(n_732) );
INVx1_ASAP7_75t_SL g478 ( .A(n_65), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_66), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_67), .B(n_162), .Y(n_504) );
INVx1_ASAP7_75t_L g462 ( .A(n_68), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_69), .Y(n_763) );
A2O1A1Ixp33_ASAP7_75t_SL g153 ( .A1(n_70), .A2(n_154), .B(n_155), .C(n_158), .Y(n_153) );
INVxp67_ASAP7_75t_L g156 ( .A(n_71), .Y(n_156) );
INVx1_ASAP7_75t_L g115 ( .A(n_72), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_73), .A2(n_140), .B(n_531), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_74), .A2(n_728), .B1(n_729), .B2(n_735), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_74), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_75), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_76), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_77), .A2(n_140), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g223 ( .A(n_78), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_79), .A2(n_248), .B(n_556), .Y(n_555) );
CKINVDCx16_ASAP7_75t_R g482 ( .A(n_80), .Y(n_482) );
INVx1_ASAP7_75t_L g520 ( .A(n_81), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_82), .A2(n_145), .B(n_149), .C(n_225), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_83), .A2(n_140), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g523 ( .A(n_84), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_85), .B(n_199), .Y(n_213) );
INVx2_ASAP7_75t_L g135 ( .A(n_86), .Y(n_135) );
INVx1_ASAP7_75t_L g513 ( .A(n_87), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_88), .B(n_154), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_89), .A2(n_145), .B(n_149), .C(n_197), .Y(n_196) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_90), .B(n_112), .C(n_113), .Y(n_111) );
INVx2_ASAP7_75t_L g122 ( .A(n_90), .Y(n_122) );
OR2x2_ASAP7_75t_L g761 ( .A(n_90), .B(n_740), .Y(n_761) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_91), .A2(n_149), .B(n_461), .C(n_465), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_92), .B(n_175), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_92), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_93), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_94), .A2(n_145), .B(n_149), .C(n_237), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g244 ( .A(n_95), .Y(n_244) );
INVx1_ASAP7_75t_L g152 ( .A(n_96), .Y(n_152) );
CKINVDCx16_ASAP7_75t_R g250 ( .A(n_97), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_98), .B(n_199), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_99), .B(n_133), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_100), .B(n_133), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_101), .B(n_115), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_102), .A2(n_140), .B(n_147), .Y(n_139) );
INVx2_ASAP7_75t_L g503 ( .A(n_103), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVx5_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
CKINVDCx9p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
BUFx2_ASAP7_75t_L g766 ( .A(n_108), .Y(n_766) );
OR2x4_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
AND2x2_ASAP7_75t_L g736 ( .A(n_112), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
AO221x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_742), .B1(n_747), .B2(n_757), .C(n_762), .Y(n_116) );
OAI22xp5_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_736), .B1(n_738), .B2(n_741), .Y(n_117) );
XOR2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_727), .Y(n_118) );
OAI22xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_123), .B1(n_449), .B2(n_450), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g449 ( .A(n_122), .Y(n_449) );
NOR2x2_ASAP7_75t_L g739 ( .A(n_122), .B(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND4x1_ASAP7_75t_L g125 ( .A(n_126), .B(n_367), .C(n_414), .D(n_434), .Y(n_125) );
NOR3xp33_ASAP7_75t_SL g126 ( .A(n_127), .B(n_297), .C(n_322), .Y(n_126) );
OAI211xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_205), .B(n_257), .C(n_287), .Y(n_127) );
INVxp67_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_130), .B(n_176), .Y(n_129) );
INVx3_ASAP7_75t_SL g339 ( .A(n_130), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_130), .B(n_270), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_130), .B(n_192), .Y(n_420) );
AND2x2_ASAP7_75t_L g443 ( .A(n_130), .B(n_309), .Y(n_443) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_164), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g261 ( .A(n_132), .B(n_165), .Y(n_261) );
INVx3_ASAP7_75t_L g274 ( .A(n_132), .Y(n_274) );
AND2x2_ASAP7_75t_L g279 ( .A(n_132), .B(n_164), .Y(n_279) );
OR2x2_ASAP7_75t_L g330 ( .A(n_132), .B(n_271), .Y(n_330) );
BUFx2_ASAP7_75t_L g350 ( .A(n_132), .Y(n_350) );
AND2x2_ASAP7_75t_L g360 ( .A(n_132), .B(n_271), .Y(n_360) );
AND2x2_ASAP7_75t_L g366 ( .A(n_132), .B(n_177), .Y(n_366) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_139), .B(n_161), .Y(n_132) );
INVx4_ASAP7_75t_L g163 ( .A(n_133), .Y(n_163) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_133), .Y(n_472) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g178 ( .A(n_134), .Y(n_178) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
AND2x2_ASAP7_75t_SL g175 ( .A(n_135), .B(n_136), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
BUFx2_ASAP7_75t_L g248 ( .A(n_140), .Y(n_248) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_145), .Y(n_140) );
NAND2x1p5_ASAP7_75t_L g189 ( .A(n_141), .B(n_145), .Y(n_189) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
INVx1_ASAP7_75t_L g488 ( .A(n_142), .Y(n_488) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g150 ( .A(n_143), .Y(n_150) );
INVx1_ASAP7_75t_L g182 ( .A(n_143), .Y(n_182) );
INVx1_ASAP7_75t_L g151 ( .A(n_144), .Y(n_151) );
INVx1_ASAP7_75t_L g154 ( .A(n_144), .Y(n_154) );
INVx3_ASAP7_75t_L g157 ( .A(n_144), .Y(n_157) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_144), .Y(n_171) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_144), .Y(n_184) );
INVx4_ASAP7_75t_SL g160 ( .A(n_145), .Y(n_160) );
BUFx3_ASAP7_75t_L g489 ( .A(n_145), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_152), .B(n_153), .C(n_160), .Y(n_147) );
O2A1O1Ixp33_ASAP7_75t_L g167 ( .A1(n_148), .A2(n_160), .B(n_168), .C(n_169), .Y(n_167) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_148), .A2(n_160), .B(n_250), .C(n_251), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_L g474 ( .A1(n_148), .A2(n_160), .B(n_475), .C(n_476), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_SL g499 ( .A1(n_148), .A2(n_160), .B(n_500), .C(n_501), .Y(n_499) );
O2A1O1Ixp33_ASAP7_75t_SL g519 ( .A1(n_148), .A2(n_160), .B(n_520), .C(n_521), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_SL g531 ( .A1(n_148), .A2(n_160), .B(n_532), .C(n_533), .Y(n_531) );
O2A1O1Ixp33_ASAP7_75t_SL g556 ( .A1(n_148), .A2(n_160), .B(n_557), .C(n_558), .Y(n_556) );
INVx5_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x6_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_150), .Y(n_159) );
BUFx3_ASAP7_75t_L g217 ( .A(n_150), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_157), .B(n_173), .Y(n_172) );
INVx5_ASAP7_75t_L g199 ( .A(n_157), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_157), .B(n_535), .Y(n_534) );
INVx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_159), .Y(n_241) );
OAI22xp33_ASAP7_75t_L g179 ( .A1(n_160), .A2(n_180), .B1(n_188), .B2(n_189), .Y(n_179) );
INVx1_ASAP7_75t_L g465 ( .A(n_160), .Y(n_465) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_162), .A2(n_166), .B(n_174), .Y(n_165) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NOR2xp33_ASAP7_75t_SL g219 ( .A(n_163), .B(n_220), .Y(n_219) );
AO21x2_ASAP7_75t_L g457 ( .A1(n_163), .A2(n_458), .B(n_466), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_163), .B(n_491), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_163), .B(n_516), .Y(n_515) );
INVx1_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_165), .B(n_271), .Y(n_285) );
INVx2_ASAP7_75t_L g295 ( .A(n_165), .Y(n_295) );
AND2x2_ASAP7_75t_L g308 ( .A(n_165), .B(n_274), .Y(n_308) );
OR2x2_ASAP7_75t_L g319 ( .A(n_165), .B(n_271), .Y(n_319) );
AND2x2_ASAP7_75t_SL g365 ( .A(n_165), .B(n_366), .Y(n_365) );
BUFx2_ASAP7_75t_L g377 ( .A(n_165), .Y(n_377) );
AND2x2_ASAP7_75t_L g423 ( .A(n_165), .B(n_177), .Y(n_423) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx4_ASAP7_75t_L g240 ( .A(n_171), .Y(n_240) );
INVx1_ASAP7_75t_L g204 ( .A(n_175), .Y(n_204) );
INVx2_ASAP7_75t_L g234 ( .A(n_175), .Y(n_234) );
OA21x2_ASAP7_75t_L g246 ( .A1(n_175), .A2(n_247), .B(n_256), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_L g481 ( .A1(n_175), .A2(n_189), .B(n_482), .C(n_483), .Y(n_481) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_175), .A2(n_530), .B(n_536), .Y(n_529) );
INVx3_ASAP7_75t_SL g296 ( .A(n_176), .Y(n_296) );
OR2x2_ASAP7_75t_L g349 ( .A(n_176), .B(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g176 ( .A(n_177), .B(n_192), .Y(n_176) );
INVx3_ASAP7_75t_L g271 ( .A(n_177), .Y(n_271) );
AND2x2_ASAP7_75t_L g338 ( .A(n_177), .B(n_193), .Y(n_338) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_177), .Y(n_406) );
AOI33xp33_ASAP7_75t_L g410 ( .A1(n_177), .A2(n_339), .A3(n_346), .B1(n_355), .B2(n_411), .B3(n_412), .Y(n_410) );
AO21x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_190), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_178), .B(n_191), .Y(n_190) );
AO21x2_ASAP7_75t_L g193 ( .A1(n_178), .A2(n_194), .B(n_202), .Y(n_193) );
INVx2_ASAP7_75t_L g218 ( .A(n_178), .Y(n_218) );
INVx2_ASAP7_75t_L g201 ( .A(n_181), .Y(n_201) );
INVx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
OAI22xp5_ASAP7_75t_SL g183 ( .A1(n_184), .A2(n_185), .B1(n_186), .B2(n_187), .Y(n_183) );
INVx2_ASAP7_75t_L g186 ( .A(n_184), .Y(n_186) );
INVx4_ASAP7_75t_L g252 ( .A(n_184), .Y(n_252) );
INVx2_ASAP7_75t_L g463 ( .A(n_186), .Y(n_463) );
OAI21xp5_ASAP7_75t_L g194 ( .A1(n_189), .A2(n_195), .B(n_196), .Y(n_194) );
OAI21xp5_ASAP7_75t_L g222 ( .A1(n_189), .A2(n_223), .B(n_224), .Y(n_222) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_189), .A2(n_459), .B(n_460), .Y(n_458) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_189), .A2(n_510), .B(n_511), .Y(n_509) );
INVx1_ASAP7_75t_L g259 ( .A(n_192), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_192), .B(n_274), .Y(n_273) );
NOR3xp33_ASAP7_75t_L g333 ( .A(n_192), .B(n_334), .C(n_336), .Y(n_333) );
AND2x2_ASAP7_75t_L g359 ( .A(n_192), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_192), .B(n_366), .Y(n_369) );
AND2x2_ASAP7_75t_L g422 ( .A(n_192), .B(n_423), .Y(n_422) );
INVx3_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx3_ASAP7_75t_L g278 ( .A(n_193), .Y(n_278) );
OR2x2_ASAP7_75t_L g372 ( .A(n_193), .B(n_271), .Y(n_372) );
O2A1O1Ixp33_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_200), .C(n_201), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g484 ( .A1(n_199), .A2(n_485), .B(n_486), .C(n_487), .Y(n_484) );
OAI22xp33_ASAP7_75t_L g559 ( .A1(n_199), .A2(n_252), .B1(n_560), .B2(n_561), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_204), .B(n_230), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_204), .B(n_244), .Y(n_243) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_204), .A2(n_509), .B(n_515), .Y(n_508) );
OR2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_231), .Y(n_205) );
AOI32xp33_ASAP7_75t_L g323 ( .A1(n_206), .A2(n_324), .A3(n_326), .B1(n_328), .B2(n_331), .Y(n_323) );
NOR2xp67_ASAP7_75t_L g396 ( .A(n_206), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g426 ( .A(n_206), .Y(n_426) );
INVx4_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g358 ( .A(n_207), .B(n_342), .Y(n_358) );
AND2x2_ASAP7_75t_L g378 ( .A(n_207), .B(n_304), .Y(n_378) );
AND2x2_ASAP7_75t_L g446 ( .A(n_207), .B(n_364), .Y(n_446) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_221), .Y(n_207) );
INVx3_ASAP7_75t_L g267 ( .A(n_208), .Y(n_267) );
AND2x2_ASAP7_75t_L g281 ( .A(n_208), .B(n_265), .Y(n_281) );
OR2x2_ASAP7_75t_L g286 ( .A(n_208), .B(n_264), .Y(n_286) );
INVx1_ASAP7_75t_L g293 ( .A(n_208), .Y(n_293) );
AND2x2_ASAP7_75t_L g301 ( .A(n_208), .B(n_275), .Y(n_301) );
AND2x2_ASAP7_75t_L g303 ( .A(n_208), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_208), .B(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g356 ( .A(n_208), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_208), .B(n_441), .Y(n_440) );
OR2x6_ASAP7_75t_L g208 ( .A(n_209), .B(n_219), .Y(n_208) );
AOI21xp5_ASAP7_75t_SL g209 ( .A1(n_210), .A2(n_211), .B(n_218), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_215), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_215), .A2(n_226), .B(n_227), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g461 ( .A1(n_215), .A2(n_462), .B(n_463), .C(n_464), .Y(n_461) );
O2A1O1Ixp5_ASAP7_75t_L g512 ( .A1(n_215), .A2(n_463), .B(n_513), .C(n_514), .Y(n_512) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g255 ( .A(n_217), .Y(n_255) );
INVx1_ASAP7_75t_L g228 ( .A(n_218), .Y(n_228) );
INVx2_ASAP7_75t_L g265 ( .A(n_221), .Y(n_265) );
AND2x2_ASAP7_75t_L g311 ( .A(n_221), .B(n_232), .Y(n_311) );
AND2x2_ASAP7_75t_L g321 ( .A(n_221), .B(n_246), .Y(n_321) );
AO21x2_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_228), .B(n_229), .Y(n_221) );
INVx1_ASAP7_75t_L g554 ( .A(n_228), .Y(n_554) );
AO21x2_ASAP7_75t_L g570 ( .A1(n_228), .A2(n_571), .B(n_572), .Y(n_570) );
INVx2_ASAP7_75t_L g441 ( .A(n_231), .Y(n_441) );
OR2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_245), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_232), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g282 ( .A(n_232), .Y(n_282) );
AND2x2_ASAP7_75t_L g326 ( .A(n_232), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g342 ( .A(n_232), .B(n_305), .Y(n_342) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g290 ( .A(n_233), .Y(n_290) );
AND2x2_ASAP7_75t_L g304 ( .A(n_233), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g355 ( .A(n_233), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_233), .B(n_265), .Y(n_387) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_243), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_234), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g563 ( .A(n_234), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_242), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B(n_241), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_240), .B(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g266 ( .A(n_245), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g327 ( .A(n_245), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_245), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g364 ( .A(n_245), .Y(n_364) );
INVx1_ASAP7_75t_L g397 ( .A(n_245), .Y(n_397) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g275 ( .A(n_246), .B(n_265), .Y(n_275) );
INVx1_ASAP7_75t_L g305 ( .A(n_246), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_252), .B(n_254), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_252), .B(n_503), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_252), .B(n_523), .Y(n_522) );
AOI221xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_262), .B1(n_268), .B2(n_275), .C(n_276), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_259), .B(n_279), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_259), .B(n_342), .Y(n_419) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_261), .B(n_309), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_261), .B(n_270), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_261), .B(n_284), .Y(n_413) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_266), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g335 ( .A(n_265), .Y(n_335) );
AND2x2_ASAP7_75t_L g310 ( .A(n_266), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g388 ( .A(n_266), .Y(n_388) );
AND2x2_ASAP7_75t_L g320 ( .A(n_267), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_267), .B(n_290), .Y(n_336) );
AND2x2_ASAP7_75t_L g400 ( .A(n_267), .B(n_326), .Y(n_400) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_272), .Y(n_269) );
BUFx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g309 ( .A(n_271), .B(n_278), .Y(n_309) );
AND2x2_ASAP7_75t_L g405 ( .A(n_272), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_274), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_275), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_275), .B(n_282), .Y(n_370) );
AND2x2_ASAP7_75t_L g390 ( .A(n_275), .B(n_290), .Y(n_390) );
AND2x2_ASAP7_75t_L g411 ( .A(n_275), .B(n_355), .Y(n_411) );
OAI32xp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_280), .A3(n_282), .B1(n_283), .B2(n_286), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx1_ASAP7_75t_SL g284 ( .A(n_278), .Y(n_284) );
NAND2x1_ASAP7_75t_L g325 ( .A(n_278), .B(n_308), .Y(n_325) );
OR2x2_ASAP7_75t_L g329 ( .A(n_278), .B(n_330), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_278), .B(n_377), .Y(n_430) );
INVx1_ASAP7_75t_L g298 ( .A(n_279), .Y(n_298) );
OAI221xp5_ASAP7_75t_SL g416 ( .A1(n_280), .A2(n_371), .B1(n_417), .B2(n_420), .C(n_421), .Y(n_416) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g288 ( .A(n_281), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g331 ( .A(n_281), .B(n_304), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_281), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g409 ( .A(n_281), .B(n_342), .Y(n_409) );
INVxp67_ASAP7_75t_L g345 ( .A(n_282), .Y(n_345) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AND2x2_ASAP7_75t_L g415 ( .A(n_284), .B(n_402), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_284), .B(n_365), .Y(n_438) );
INVx1_ASAP7_75t_L g313 ( .A(n_286), .Y(n_313) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_286), .B(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g431 ( .A(n_286), .B(n_432), .Y(n_431) );
OAI21xp5_ASAP7_75t_SL g287 ( .A1(n_288), .A2(n_291), .B(n_294), .Y(n_287) );
AND2x2_ASAP7_75t_L g300 ( .A(n_289), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g384 ( .A(n_293), .B(n_304), .Y(n_384) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
AND2x2_ASAP7_75t_L g402 ( .A(n_295), .B(n_360), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_295), .B(n_359), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_296), .B(n_308), .Y(n_382) );
OAI211xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B(n_302), .C(n_312), .Y(n_297) );
AOI221xp5_ASAP7_75t_L g332 ( .A1(n_298), .A2(n_333), .B1(n_337), .B2(n_340), .C(n_343), .Y(n_332) );
AOI31xp33_ASAP7_75t_L g427 ( .A1(n_298), .A2(n_428), .A3(n_429), .B(n_431), .Y(n_427) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_306), .B1(n_308), .B2(n_310), .Y(n_302) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx1_ASAP7_75t_L g428 ( .A(n_308), .Y(n_428) );
INVx1_ASAP7_75t_L g391 ( .A(n_309), .Y(n_391) );
O2A1O1Ixp33_ASAP7_75t_L g434 ( .A1(n_311), .A2(n_435), .B(n_437), .C(n_439), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_314), .B1(n_316), .B2(n_320), .Y(n_312) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_317), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OAI221xp5_ASAP7_75t_SL g407 ( .A1(n_319), .A2(n_353), .B1(n_372), .B2(n_408), .C(n_410), .Y(n_407) );
INVx1_ASAP7_75t_L g403 ( .A(n_320), .Y(n_403) );
INVx1_ASAP7_75t_L g357 ( .A(n_321), .Y(n_357) );
NAND3xp33_ASAP7_75t_SL g322 ( .A(n_323), .B(n_332), .C(n_347), .Y(n_322) );
OAI21xp33_ASAP7_75t_L g373 ( .A1(n_324), .A2(n_374), .B(n_378), .Y(n_373) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_326), .B(n_426), .Y(n_425) );
INVxp67_ASAP7_75t_L g433 ( .A(n_327), .Y(n_433) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g371 ( .A(n_334), .B(n_354), .Y(n_371) );
INVx1_ASAP7_75t_L g346 ( .A(n_335), .Y(n_346) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx1_ASAP7_75t_L g344 ( .A(n_338), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_338), .B(n_376), .Y(n_375) );
NOR4xp25_ASAP7_75t_L g343 ( .A(n_339), .B(n_344), .C(n_345), .D(n_346), .Y(n_343) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AOI222xp33_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_352), .B1(n_358), .B2(n_359), .C1(n_361), .C2(n_365), .Y(n_347) );
NAND2xp5_ASAP7_75t_SL g348 ( .A(n_349), .B(n_351), .Y(n_348) );
INVx1_ASAP7_75t_L g445 ( .A(n_349), .Y(n_445) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_357), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_361), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OAI21xp5_ASAP7_75t_SL g421 ( .A1(n_366), .A2(n_422), .B(n_424), .Y(n_421) );
NOR4xp25_ASAP7_75t_L g367 ( .A(n_368), .B(n_379), .C(n_392), .D(n_407), .Y(n_367) );
OAI221xp5_ASAP7_75t_SL g368 ( .A1(n_369), .A2(n_370), .B1(n_371), .B2(n_372), .C(n_373), .Y(n_368) );
INVx1_ASAP7_75t_L g448 ( .A(n_369), .Y(n_448) );
INVx1_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_376), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
OAI222xp33_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_383), .B1(n_385), .B2(n_386), .C1(n_389), .C2(n_391), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AOI211xp5_ASAP7_75t_L g414 ( .A1(n_384), .A2(n_415), .B(n_416), .C(n_427), .Y(n_414) );
OR2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
INVx1_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
OAI222xp33_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_398), .B1(n_399), .B2(n_401), .C1(n_403), .C2(n_404), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVxp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_409), .A2(n_412), .B1(n_445), .B2(n_446), .Y(n_444) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OAI211xp5_ASAP7_75t_SL g439 ( .A1(n_440), .A2(n_442), .B(n_444), .C(n_447), .Y(n_439) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
XNOR2xp5_ASAP7_75t_L g748 ( .A(n_450), .B(n_749), .Y(n_748) );
AND2x2_ASAP7_75t_SL g450 ( .A(n_451), .B(n_682), .Y(n_450) );
NOR4xp25_ASAP7_75t_L g451 ( .A(n_452), .B(n_619), .C(n_653), .D(n_669), .Y(n_451) );
NAND4xp25_ASAP7_75t_SL g452 ( .A(n_453), .B(n_549), .C(n_583), .D(n_599), .Y(n_452) );
AOI222xp33_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_492), .B1(n_525), .B2(n_537), .C1(n_542), .C2(n_548), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AOI31xp33_ASAP7_75t_L g715 ( .A1(n_455), .A2(n_716), .A3(n_717), .B(n_719), .Y(n_715) );
OR2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_468), .Y(n_455) );
AND2x2_ASAP7_75t_L g690 ( .A(n_456), .B(n_470), .Y(n_690) );
BUFx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_SL g541 ( .A(n_457), .Y(n_541) );
AND2x2_ASAP7_75t_L g548 ( .A(n_457), .B(n_480), .Y(n_548) );
AND2x2_ASAP7_75t_L g604 ( .A(n_457), .B(n_471), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_468), .B(n_634), .Y(n_633) );
INVx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_469), .B(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_469), .B(n_552), .Y(n_594) );
AND2x2_ASAP7_75t_L g687 ( .A(n_469), .B(n_627), .Y(n_687) );
OAI321xp33_ASAP7_75t_L g721 ( .A1(n_469), .A2(n_541), .A3(n_694), .B1(n_722), .B2(n_724), .C(n_725), .Y(n_721) );
NAND4xp25_ASAP7_75t_L g725 ( .A(n_469), .B(n_528), .C(n_634), .D(n_726), .Y(n_725) );
AND2x4_ASAP7_75t_L g469 ( .A(n_470), .B(n_480), .Y(n_469) );
AND2x2_ASAP7_75t_L g589 ( .A(n_470), .B(n_539), .Y(n_589) );
AND2x2_ASAP7_75t_L g608 ( .A(n_470), .B(n_541), .Y(n_608) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g540 ( .A(n_471), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g564 ( .A(n_471), .B(n_480), .Y(n_564) );
AND2x2_ASAP7_75t_L g650 ( .A(n_471), .B(n_539), .Y(n_650) );
OA21x2_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B(n_479), .Y(n_471) );
OA21x2_ASAP7_75t_L g497 ( .A1(n_472), .A2(n_498), .B(n_504), .Y(n_497) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_472), .A2(n_518), .B(n_524), .Y(n_517) );
INVx3_ASAP7_75t_SL g539 ( .A(n_480), .Y(n_539) );
AND2x2_ASAP7_75t_L g582 ( .A(n_480), .B(n_569), .Y(n_582) );
OR2x2_ASAP7_75t_L g615 ( .A(n_480), .B(n_541), .Y(n_615) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_480), .Y(n_622) );
AND2x2_ASAP7_75t_L g651 ( .A(n_480), .B(n_540), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_480), .B(n_624), .Y(n_666) );
AND2x2_ASAP7_75t_L g698 ( .A(n_480), .B(n_690), .Y(n_698) );
AND2x2_ASAP7_75t_L g707 ( .A(n_480), .B(n_553), .Y(n_707) );
OR2x6_ASAP7_75t_L g480 ( .A(n_481), .B(n_490), .Y(n_480) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_488), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_505), .Y(n_493) );
INVx1_ASAP7_75t_SL g675 ( .A(n_494), .Y(n_675) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g544 ( .A(n_495), .B(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g527 ( .A(n_496), .B(n_507), .Y(n_527) );
AND2x2_ASAP7_75t_L g611 ( .A(n_496), .B(n_529), .Y(n_611) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g581 ( .A(n_497), .B(n_517), .Y(n_581) );
OR2x2_ASAP7_75t_L g592 ( .A(n_497), .B(n_529), .Y(n_592) );
AND2x2_ASAP7_75t_L g618 ( .A(n_497), .B(n_529), .Y(n_618) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_497), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_505), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_505), .B(n_675), .Y(n_674) );
INVx2_ASAP7_75t_SL g505 ( .A(n_506), .Y(n_505) );
OR2x2_ASAP7_75t_L g591 ( .A(n_506), .B(n_592), .Y(n_591) );
AOI322xp5_ASAP7_75t_L g677 ( .A1(n_506), .A2(n_581), .A3(n_587), .B1(n_618), .B2(n_668), .C1(n_678), .C2(n_680), .Y(n_677) );
OR2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_517), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_507), .B(n_528), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_507), .B(n_529), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_507), .B(n_545), .Y(n_598) );
AND2x2_ASAP7_75t_L g652 ( .A(n_507), .B(n_618), .Y(n_652) );
INVx1_ASAP7_75t_L g656 ( .A(n_507), .Y(n_656) );
AND2x2_ASAP7_75t_L g668 ( .A(n_507), .B(n_517), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_507), .B(n_544), .Y(n_700) );
INVx4_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g565 ( .A(n_508), .B(n_517), .Y(n_565) );
BUFx3_ASAP7_75t_L g579 ( .A(n_508), .Y(n_579) );
AND3x2_ASAP7_75t_L g661 ( .A(n_508), .B(n_641), .C(n_662), .Y(n_661) );
NAND3xp33_ASAP7_75t_L g526 ( .A(n_517), .B(n_527), .C(n_528), .Y(n_526) );
INVx1_ASAP7_75t_SL g545 ( .A(n_517), .Y(n_545) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_517), .Y(n_646) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g640 ( .A(n_527), .B(n_641), .Y(n_640) );
INVxp67_ASAP7_75t_L g647 ( .A(n_527), .Y(n_647) );
AND2x2_ASAP7_75t_L g685 ( .A(n_528), .B(n_663), .Y(n_685) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
BUFx3_ASAP7_75t_L g566 ( .A(n_529), .Y(n_566) );
AND2x2_ASAP7_75t_L g641 ( .A(n_529), .B(n_545), .Y(n_641) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
OR2x2_ASAP7_75t_L g585 ( .A(n_539), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g704 ( .A(n_539), .B(n_604), .Y(n_704) );
AND2x2_ASAP7_75t_L g718 ( .A(n_539), .B(n_541), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_540), .B(n_553), .Y(n_659) );
AND2x2_ASAP7_75t_L g706 ( .A(n_540), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g569 ( .A(n_541), .B(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g586 ( .A(n_541), .B(n_553), .Y(n_586) );
INVx1_ASAP7_75t_L g596 ( .A(n_541), .Y(n_596) );
AND2x2_ASAP7_75t_L g627 ( .A(n_541), .B(n_553), .Y(n_627) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
OAI221xp5_ASAP7_75t_L g669 ( .A1(n_543), .A2(n_670), .B1(n_674), .B2(n_676), .C(n_677), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_544), .B(n_546), .Y(n_543) );
AND2x2_ASAP7_75t_L g573 ( .A(n_544), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_547), .B(n_580), .Y(n_723) );
AOI322xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_565), .A3(n_566), .B1(n_567), .B2(n_573), .C1(n_575), .C2(n_582), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_564), .Y(n_551) );
NAND2x1p5_ASAP7_75t_L g603 ( .A(n_552), .B(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_552), .B(n_614), .Y(n_613) );
O2A1O1Ixp33_ASAP7_75t_L g637 ( .A1(n_552), .A2(n_564), .B(n_638), .C(n_639), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_552), .B(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_552), .B(n_608), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_552), .B(n_690), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_552), .B(n_718), .Y(n_717) );
BUFx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_553), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_553), .B(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g679 ( .A(n_553), .B(n_566), .Y(n_679) );
OA21x2_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_555), .B(n_562), .Y(n_553) );
INVx1_ASAP7_75t_L g571 ( .A(n_555), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_562), .Y(n_572) );
INVx1_ASAP7_75t_L g654 ( .A(n_564), .Y(n_654) );
OAI31xp33_ASAP7_75t_L g664 ( .A1(n_564), .A2(n_589), .A3(n_665), .B(n_667), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_564), .B(n_570), .Y(n_716) );
INVx1_ASAP7_75t_SL g577 ( .A(n_565), .Y(n_577) );
AND2x2_ASAP7_75t_L g610 ( .A(n_565), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g691 ( .A(n_565), .B(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g576 ( .A(n_566), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g601 ( .A(n_566), .Y(n_601) );
AND2x2_ASAP7_75t_L g628 ( .A(n_566), .B(n_581), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_566), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g720 ( .A(n_566), .B(n_668), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_568), .B(n_638), .Y(n_711) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g607 ( .A(n_570), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_SL g625 ( .A(n_570), .Y(n_625) );
NAND2xp33_ASAP7_75t_SL g575 ( .A(n_576), .B(n_578), .Y(n_575) );
OAI211xp5_ASAP7_75t_SL g619 ( .A1(n_577), .A2(n_620), .B(n_626), .C(n_642), .Y(n_619) );
OR2x2_ASAP7_75t_L g694 ( .A(n_577), .B(n_675), .Y(n_694) );
OR2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
CKINVDCx16_ASAP7_75t_R g631 ( .A(n_579), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_579), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g600 ( .A(n_581), .B(n_601), .Y(n_600) );
O2A1O1Ixp33_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_587), .B(n_590), .C(n_593), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_SL g634 ( .A(n_586), .Y(n_634) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_589), .B(n_627), .Y(n_632) );
INVx1_ASAP7_75t_L g638 ( .A(n_589), .Y(n_638) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g597 ( .A(n_592), .B(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g630 ( .A(n_592), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g692 ( .A(n_592), .Y(n_692) );
AOI21xp33_ASAP7_75t_SL g593 ( .A1(n_594), .A2(n_595), .B(n_597), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g605 ( .A1(n_595), .A2(n_606), .B(n_609), .Y(n_605) );
AOI211xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_602), .B(n_605), .C(n_612), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_600), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_603), .B(n_694), .Y(n_693) );
INVx2_ASAP7_75t_SL g616 ( .A(n_604), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g671 ( .A1(n_606), .A2(n_672), .B(n_673), .Y(n_671) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_611), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_SL g636 ( .A(n_611), .Y(n_636) );
AOI21xp33_ASAP7_75t_SL g612 ( .A1(n_613), .A2(n_616), .B(n_617), .Y(n_612) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g667 ( .A(n_618), .B(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_624), .B(n_650), .Y(n_676) );
AND2x2_ASAP7_75t_L g689 ( .A(n_624), .B(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g703 ( .A(n_624), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g713 ( .A(n_624), .B(n_651), .Y(n_713) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AOI211xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_628), .B(n_629), .C(n_637), .Y(n_626) );
INVx1_ASAP7_75t_L g673 ( .A(n_627), .Y(n_673) );
OAI22xp33_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_632), .B1(n_633), .B2(n_635), .Y(n_629) );
OR2x2_ASAP7_75t_L g635 ( .A(n_631), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g714 ( .A(n_631), .B(n_692), .Y(n_714) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g708 ( .A(n_641), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_648), .B1(n_651), .B2(n_652), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
INVx1_ASAP7_75t_L g726 ( .A(n_646), .Y(n_726) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g672 ( .A(n_650), .Y(n_672) );
OAI211xp5_ASAP7_75t_SL g653 ( .A1(n_654), .A2(n_655), .B(n_657), .C(n_664), .Y(n_653) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
INVx2_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
INVxp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVxp67_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_672), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NOR5xp2_ASAP7_75t_L g682 ( .A(n_683), .B(n_701), .C(n_709), .D(n_715), .E(n_721), .Y(n_682) );
OAI211xp5_ASAP7_75t_SL g683 ( .A1(n_684), .A2(n_686), .B(n_688), .C(n_695), .Y(n_683) );
INVxp67_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_691), .B(n_693), .Y(n_688) );
OAI21xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_698), .B(n_699), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_698), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AOI21xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_705), .B(n_708), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_SL g724 ( .A(n_704), .Y(n_724) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_712), .B(n_714), .Y(n_709) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g740 ( .A(n_736), .Y(n_740) );
INVx3_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVxp67_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
BUFx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g758 ( .A(n_746), .Y(n_758) );
OAI22xp5_ASAP7_75t_SL g747 ( .A1(n_748), .A2(n_752), .B1(n_753), .B2(n_756), .Y(n_747) );
INVx1_ASAP7_75t_L g756 ( .A(n_748), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_753), .Y(n_752) );
NOR2xp33_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g765 ( .A(n_761), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
endmodule