module fake_jpeg_3483_n_106 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_106);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_9),
.Y(n_11)
);

INVx13_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx4f_ASAP7_75t_SL g14 ( 
.A(n_0),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_22),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_19),
.B(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_11),
.B(n_3),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_SL g55 ( 
.A(n_34),
.Y(n_55)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_11),
.B(n_25),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_4),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_38),
.B(n_17),
.Y(n_45)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_21),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_26),
.B(n_23),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_46),
.B(n_30),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_27),
.A2(n_15),
.B1(n_17),
.B2(n_23),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_5),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_29),
.A2(n_16),
.B1(n_20),
.B2(n_18),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_34),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_16),
.B1(n_20),
.B2(n_18),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_21),
.B1(n_6),
.B2(n_8),
.Y(n_52)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_64),
.Y(n_74)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_73),
.B1(n_67),
.B2(n_51),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_59),
.B(n_53),
.C(n_43),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_69),
.B(n_70),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_34),
.B(n_37),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_67),
.A2(n_48),
.B(n_51),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_68),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_49),
.B(n_47),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_42),
.B(n_30),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_72),
.Y(n_76)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_47),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_68),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_71),
.B1(n_60),
.B2(n_48),
.Y(n_87)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_88),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_77),
.A2(n_73),
.B(n_71),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_86),
.A2(n_76),
.B(n_74),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_10),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_48),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_85),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_95),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_94),
.Y(n_97)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_90),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_99),
.A2(n_100),
.B(n_91),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_97),
.A2(n_85),
.B1(n_91),
.B2(n_81),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_98),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_102),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_78),
.C(n_82),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_79),
.Y(n_106)
);


endmodule