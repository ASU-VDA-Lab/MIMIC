module fake_jpeg_2581_n_431 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_431);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_431;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_SL g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_42),
.B(n_51),
.Y(n_109)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_43),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_44),
.B(n_47),
.Y(n_99)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_0),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_50),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_32),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

NAND2x1_ASAP7_75t_SL g97 ( 
.A(n_52),
.B(n_68),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_53),
.B(n_57),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_14),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_54),
.B(n_59),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_21),
.Y(n_58)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_35),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_62),
.Y(n_98)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_33),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_65),
.B(n_70),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_31),
.B(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_73),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_31),
.B(n_0),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_18),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_18),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_27),
.B(n_1),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_75),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_18),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_19),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_79),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_19),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_19),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_25),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_67),
.A2(n_17),
.B1(n_27),
.B2(n_28),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_90),
.A2(n_92),
.B1(n_110),
.B2(n_79),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_47),
.A2(n_27),
.B1(n_28),
.B2(n_38),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_93),
.B(n_114),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_58),
.A2(n_29),
.B1(n_28),
.B2(n_38),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_96),
.A2(n_124),
.B1(n_125),
.B2(n_21),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_74),
.A2(n_17),
.B1(n_37),
.B2(n_36),
.Y(n_110)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_46),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_115),
.B(n_116),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_45),
.B(n_25),
.C(n_20),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_49),
.Y(n_117)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_119),
.B(n_61),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_70),
.A2(n_24),
.B1(n_22),
.B2(n_37),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_120),
.A2(n_22),
.B1(n_24),
.B2(n_23),
.Y(n_156)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_58),
.Y(n_122)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_68),
.B(n_38),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_123),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_65),
.A2(n_29),
.B1(n_17),
.B2(n_36),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_68),
.A2(n_29),
.B1(n_37),
.B2(n_36),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_43),
.B(n_44),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_126),
.A2(n_141),
.B(n_41),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_100),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_127),
.B(n_146),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_80),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_128),
.B(n_133),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_129),
.A2(n_150),
.B1(n_163),
.B2(n_98),
.Y(n_174)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_130),
.Y(n_189)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_132),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_91),
.B(n_78),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_134),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_83),
.B(n_75),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_136),
.B(n_140),
.Y(n_202)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_83),
.B(n_73),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_43),
.B(n_51),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_145),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_99),
.B(n_64),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_57),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_147),
.B(n_149),
.Y(n_199)
);

AOI21xp33_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_43),
.B(n_34),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_148),
.A2(n_161),
.B(n_164),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_82),
.B(n_59),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_92),
.A2(n_62),
.B1(n_55),
.B2(n_56),
.Y(n_150)
);

BUFx2_ASAP7_75t_SL g152 ( 
.A(n_122),
.Y(n_152)
);

BUFx2_ASAP7_75t_SL g190 ( 
.A(n_152),
.Y(n_190)
);

INVxp33_ASAP7_75t_L g153 ( 
.A(n_109),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_82),
.B(n_53),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_154),
.B(n_155),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_112),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_156),
.A2(n_162),
.B1(n_86),
.B2(n_24),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_101),
.B(n_60),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_160),
.B(n_165),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_116),
.B(n_61),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_123),
.A2(n_48),
.B1(n_71),
.B2(n_69),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_94),
.A2(n_63),
.B1(n_72),
.B2(n_66),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_106),
.B(n_61),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_106),
.B(n_50),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_166),
.B(n_167),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_97),
.B(n_66),
.Y(n_167)
);

AOI21xp33_ASAP7_75t_L g168 ( 
.A1(n_97),
.A2(n_34),
.B(n_52),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_86),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_169),
.A2(n_173),
.B1(n_208),
.B2(n_137),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_172),
.A2(n_191),
.B(n_196),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_156),
.A2(n_98),
.B1(n_22),
.B2(n_23),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_174),
.A2(n_180),
.B1(n_187),
.B2(n_162),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_102),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_176),
.Y(n_226)
);

O2A1O1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_128),
.A2(n_89),
.B(n_103),
.C(n_113),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_179),
.A2(n_193),
.B(n_126),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_129),
.A2(n_102),
.B1(n_117),
.B2(n_88),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_185),
.Y(n_223)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_138),
.Y(n_186)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_186),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_127),
.A2(n_104),
.B1(n_94),
.B2(n_111),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_104),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_192),
.Y(n_224)
);

O2A1O1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_133),
.A2(n_89),
.B(n_103),
.C(n_113),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_141),
.B(n_95),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_135),
.B(n_164),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_135),
.C(n_161),
.Y(n_217)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_142),
.Y(n_201)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_201),
.Y(n_238)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_143),
.Y(n_203)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_203),
.Y(n_240)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_132),
.Y(n_205)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_205),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_150),
.A2(n_111),
.B1(n_108),
.B2(n_84),
.Y(n_208)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_209),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_211),
.Y(n_250)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_171),
.Y(n_212)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_212),
.Y(n_277)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_171),
.Y(n_213)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_213),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_140),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_235),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_191),
.A2(n_136),
.B(n_157),
.Y(n_216)
);

OAI21xp33_ASAP7_75t_L g255 ( 
.A1(n_216),
.A2(n_242),
.B(n_181),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_217),
.B(n_184),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_188),
.B(n_147),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_218),
.B(n_220),
.Y(n_252)
);

BUFx12_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_219),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_202),
.B(n_146),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_221),
.Y(n_272)
);

A2O1A1O1Ixp25_ASAP7_75t_L g222 ( 
.A1(n_198),
.A2(n_149),
.B(n_154),
.C(n_151),
.D(n_137),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_222),
.B(n_245),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_225),
.A2(n_227),
.B1(n_234),
.B2(n_237),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_197),
.A2(n_144),
.B1(n_108),
.B2(n_130),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_185),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_229),
.B(n_231),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_180),
.A2(n_163),
.B1(n_159),
.B2(n_131),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_230),
.A2(n_236),
.B1(n_239),
.B2(n_241),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_207),
.B(n_139),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_177),
.B(n_145),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_232),
.B(n_233),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_179),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_202),
.A2(n_130),
.B1(n_131),
.B2(n_84),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_193),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_199),
.A2(n_121),
.B1(n_81),
.B2(n_34),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_182),
.A2(n_23),
.B1(n_81),
.B2(n_121),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_182),
.A2(n_113),
.B1(n_21),
.B2(n_39),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_169),
.A2(n_113),
.B1(n_21),
.B2(n_39),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_177),
.B(n_15),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_200),
.A2(n_21),
.B1(n_39),
.B2(n_16),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_243),
.A2(n_208),
.B1(n_178),
.B2(n_183),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_170),
.B(n_1),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_184),
.Y(n_269)
);

A2O1A1O1Ixp25_ASAP7_75t_L g245 ( 
.A1(n_200),
.A2(n_21),
.B(n_15),
.C(n_14),
.D(n_16),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_170),
.Y(n_246)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_246),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_196),
.C(n_192),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_249),
.B(n_253),
.C(n_271),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_216),
.B(n_206),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_255),
.B(n_268),
.Y(n_292)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_258),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_233),
.A2(n_196),
.B1(n_192),
.B2(n_186),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_259),
.A2(n_211),
.B(n_224),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_260),
.A2(n_227),
.B1(n_234),
.B2(n_228),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_235),
.A2(n_187),
.B1(n_183),
.B2(n_203),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_261),
.A2(n_264),
.B1(n_213),
.B2(n_212),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_214),
.B(n_178),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_262),
.B(n_276),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_209),
.A2(n_201),
.B1(n_195),
.B2(n_189),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_223),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_278),
.Y(n_294)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_238),
.Y(n_270)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_210),
.B(n_194),
.C(n_175),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_243),
.C(n_229),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_226),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_274),
.B(n_1),
.Y(n_310)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_240),
.Y(n_275)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_210),
.B(n_175),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_205),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_240),
.Y(n_279)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

AO22x1_ASAP7_75t_SL g280 ( 
.A1(n_224),
.A2(n_204),
.B1(n_189),
.B2(n_190),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_280),
.B(n_281),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_231),
.B(n_204),
.Y(n_281)
);

OAI21xp33_ASAP7_75t_L g322 ( 
.A1(n_282),
.A2(n_288),
.B(n_309),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_257),
.A2(n_241),
.B1(n_230),
.B2(n_222),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_283),
.A2(n_248),
.B1(n_260),
.B2(n_281),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_263),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_284),
.B(n_293),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_246),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_286),
.B(n_269),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_276),
.Y(n_288)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_288),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_289),
.A2(n_291),
.B1(n_299),
.B2(n_305),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_257),
.A2(n_247),
.B1(n_248),
.B2(n_250),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_247),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_295),
.B(n_301),
.C(n_303),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_228),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_297),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_245),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_298),
.Y(n_323)
);

INVx3_ASAP7_75t_SL g300 ( 
.A(n_277),
.Y(n_300)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_300),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_249),
.B(n_236),
.C(n_215),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_253),
.B(n_239),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_273),
.B(n_215),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_308),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_251),
.A2(n_221),
.B1(n_219),
.B2(n_3),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_251),
.A2(n_219),
.B1(n_2),
.B2(n_3),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_306),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_277),
.Y(n_308)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_310),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_285),
.B(n_262),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_312),
.B(n_313),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_290),
.B(n_265),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_285),
.B(n_259),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_315),
.B(n_322),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_291),
.A2(n_309),
.B1(n_289),
.B2(n_298),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_317),
.A2(n_321),
.B1(n_334),
.B2(n_283),
.Y(n_338)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_287),
.Y(n_320)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_320),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_324),
.B(n_325),
.C(n_326),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_286),
.B(n_254),
.C(n_256),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_290),
.B(n_252),
.Y(n_326)
);

AOI21xp33_ASAP7_75t_L g327 ( 
.A1(n_292),
.A2(n_254),
.B(n_278),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_327),
.B(n_302),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_282),
.A2(n_266),
.B(n_261),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_328),
.A2(n_297),
.B(n_304),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_303),
.B(n_267),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_331),
.B(n_335),
.C(n_295),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_294),
.B(n_267),
.Y(n_333)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_333),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_298),
.A2(n_264),
.B1(n_272),
.B2(n_4),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_301),
.B(n_272),
.Y(n_335)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_336),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_319),
.A2(n_297),
.B(n_304),
.Y(n_337)
);

OAI21x1_ASAP7_75t_SL g371 ( 
.A1(n_337),
.A2(n_332),
.B(n_296),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_338),
.A2(n_354),
.B1(n_347),
.B2(n_339),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_318),
.B(n_307),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_340),
.B(n_343),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_287),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_344),
.A2(n_349),
.B(n_351),
.Y(n_360)
);

INVxp33_ASAP7_75t_SL g345 ( 
.A(n_317),
.Y(n_345)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_345),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_346),
.B(n_325),
.Y(n_367)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_333),
.Y(n_347)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_347),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_328),
.A2(n_294),
.B(n_302),
.Y(n_349)
);

BUFx24_ASAP7_75t_SL g350 ( 
.A(n_326),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_350),
.B(n_357),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_323),
.A2(n_308),
.B(n_300),
.Y(n_351)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_314),
.Y(n_353)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_353),
.Y(n_376)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_311),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_355),
.B(n_324),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_335),
.B(n_296),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_311),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_358),
.B(n_3),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_346),
.B(n_316),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_361),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_338),
.A2(n_321),
.B1(n_329),
.B2(n_334),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_362),
.A2(n_370),
.B1(n_375),
.B2(n_341),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_342),
.B(n_316),
.C(n_331),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_363),
.B(n_365),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_364),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_342),
.B(n_315),
.C(n_312),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_367),
.B(n_352),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_356),
.B(n_313),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_368),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_348),
.B(n_356),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_369),
.B(n_365),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_371),
.A2(n_374),
.B(n_10),
.Y(n_386)
);

A2O1A1O1Ixp25_ASAP7_75t_L g374 ( 
.A1(n_339),
.A2(n_332),
.B(n_6),
.C(n_7),
.D(n_8),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_359),
.A2(n_349),
.B1(n_355),
.B2(n_337),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_377),
.B(n_381),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_361),
.B(n_348),
.C(n_351),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_378),
.B(n_383),
.Y(n_399)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_380),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_362),
.A2(n_353),
.B1(n_341),
.B2(n_344),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_382),
.B(n_385),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_373),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_363),
.B(n_6),
.C(n_9),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_386),
.B(n_387),
.Y(n_402)
);

FAx1_ASAP7_75t_SL g387 ( 
.A(n_360),
.B(n_364),
.CI(n_368),
.CON(n_387),
.SN(n_387)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_390),
.B(n_366),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_377),
.A2(n_360),
.B(n_374),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_391),
.B(n_393),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_384),
.B(n_367),
.C(n_369),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_396),
.B(n_397),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_378),
.B(n_376),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_379),
.B(n_372),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_398),
.B(n_383),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_388),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_400),
.B(n_385),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_389),
.B(n_11),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_401),
.B(n_11),
.Y(n_413)
);

CKINVDCx14_ASAP7_75t_R g403 ( 
.A(n_381),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_403),
.B(n_402),
.Y(n_404)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_404),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_397),
.Y(n_406)
);

OAI21x1_ASAP7_75t_L g417 ( 
.A1(n_406),
.A2(n_409),
.B(n_411),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_396),
.B(n_399),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_408),
.B(n_410),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_392),
.B(n_387),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_393),
.B(n_394),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_412),
.A2(n_387),
.B(n_401),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_413),
.B(n_391),
.Y(n_415)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_415),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_405),
.B(n_402),
.C(n_395),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_416),
.B(n_404),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_407),
.B(n_395),
.Y(n_418)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_418),
.Y(n_425)
);

AOI21xp33_ASAP7_75t_L g422 ( 
.A1(n_419),
.A2(n_420),
.B(n_414),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g426 ( 
.A(n_421),
.B(n_422),
.Y(n_426)
);

NAND2x1_ASAP7_75t_L g423 ( 
.A(n_417),
.B(n_11),
.Y(n_423)
);

A2O1A1O1Ixp25_ASAP7_75t_L g427 ( 
.A1(n_423),
.A2(n_11),
.B(n_12),
.C(n_13),
.D(n_415),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_427),
.B(n_423),
.C(n_424),
.Y(n_428)
);

OAI321xp33_ASAP7_75t_L g429 ( 
.A1(n_428),
.A2(n_426),
.A3(n_425),
.B1(n_418),
.B2(n_13),
.C(n_12),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_429),
.B(n_13),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_430),
.B(n_13),
.Y(n_431)
);


endmodule