module fake_ariane_1609_n_1274 (n_295, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_294, n_197, n_176, n_34, n_172, n_183, n_299, n_12, n_133, n_66, n_205, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_214, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_327, n_77, n_15, n_23, n_87, n_279, n_207, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_267, n_291, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_11, n_129, n_126, n_282, n_328, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_238, n_136, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_221, n_321, n_86, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_324, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_26, n_246, n_0, n_159, n_105, n_30, n_131, n_263, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_258, n_118, n_121, n_22, n_241, n_29, n_191, n_80, n_211, n_97, n_322, n_251, n_116, n_39, n_155, n_127, n_1274);

input n_295;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_214;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_327;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_267;
input n_291;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_238;
input n_136;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_221;
input n_321;
input n_86;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_324;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_26;
input n_246;
input n_0;
input n_159;
input n_105;
input n_30;
input n_131;
input n_263;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_258;
input n_118;
input n_121;
input n_22;
input n_241;
input n_29;
input n_191;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_39;
input n_155;
input n_127;

output n_1274;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_423;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_338;
wire n_995;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1018;
wire n_953;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_868;
wire n_884;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_611;
wire n_365;
wire n_1013;
wire n_334;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1213;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_461;
wire n_1121;
wire n_490;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1108;
wire n_355;
wire n_444;
wire n_851;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_513;
wire n_1178;
wire n_1026;
wire n_436;
wire n_669;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_967;
wire n_1083;
wire n_746;
wire n_1079;
wire n_615;
wire n_1139;
wire n_517;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_836;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_776;
wire n_424;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_553;
wire n_814;
wire n_578;
wire n_405;
wire n_1134;
wire n_647;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1061;
wire n_681;
wire n_874;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_957;
wire n_388;
wire n_1242;
wire n_1218;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1189;
wire n_1089;
wire n_735;
wire n_1005;
wire n_527;
wire n_845;
wire n_888;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1266;
wire n_769;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_999;
wire n_456;
wire n_852;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1243;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_1257;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_687;
wire n_797;
wire n_480;
wire n_642;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_730;
wire n_386;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_752;
wire n_985;
wire n_421;
wire n_906;
wire n_1180;
wire n_806;
wire n_649;
wire n_374;
wire n_643;
wire n_682;
wire n_819;
wire n_586;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_420;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_617;
wire n_543;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_613;
wire n_1022;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_493;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_1183;
wire n_981;
wire n_1110;
wire n_1204;
wire n_994;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1057;
wire n_1011;
wire n_978;
wire n_828;
wire n_558;
wire n_653;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_332;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_679;
wire n_663;
wire n_443;
wire n_528;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1064;
wire n_633;
wire n_900;
wire n_1093;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_835;
wire n_446;
wire n_1076;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_550;
wire n_997;
wire n_635;
wire n_694;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_671;
wire n_1148;
wire n_654;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_658;
wire n_630;
wire n_362;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_371;
wire n_1114;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_895;
wire n_583;
wire n_1000;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1232;
wire n_996;
wire n_1211;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1001;
wire n_1115;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_340;
wire n_548;
wire n_523;
wire n_457;
wire n_782;
wire n_364;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_573;
wire n_796;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_255),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_107),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_191),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_266),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_143),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_103),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_319),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_185),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_194),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_102),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_181),
.B(n_7),
.Y(n_340)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_123),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_20),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_286),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_91),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_19),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_170),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_118),
.Y(n_347)
);

NOR2xp67_ASAP7_75t_L g348 ( 
.A(n_6),
.B(n_214),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_239),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_106),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_77),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_57),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_126),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_195),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_263),
.Y(n_355)
);

BUFx10_ASAP7_75t_L g356 ( 
.A(n_99),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_177),
.Y(n_357)
);

INVxp33_ASAP7_75t_SL g358 ( 
.A(n_21),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_251),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_173),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_96),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_211),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_55),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_293),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_109),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_321),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_131),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_47),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_213),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_193),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_278),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_172),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_304),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_163),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_250),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_171),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_60),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_129),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_287),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_329),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_152),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_188),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_256),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_318),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_259),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_20),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_124),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g388 ( 
.A(n_325),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_108),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_60),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_226),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_288),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_208),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_174),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_55),
.Y(n_395)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_82),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_48),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_96),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_313),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_159),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_7),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_11),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_149),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_52),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_176),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_276),
.Y(n_406)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_178),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_182),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_168),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_190),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_142),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_230),
.Y(n_412)
);

CKINVDCx14_ASAP7_75t_R g413 ( 
.A(n_224),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_183),
.Y(n_414)
);

CKINVDCx14_ASAP7_75t_R g415 ( 
.A(n_220),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_17),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_157),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_236),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_179),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_243),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_267),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_104),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_121),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_145),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_283),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_32),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_262),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_302),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_161),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_97),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_86),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_257),
.Y(n_432)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_303),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_94),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_99),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_139),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_299),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_202),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_252),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_175),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_127),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_34),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_180),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_317),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_128),
.Y(n_445)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_147),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_212),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_192),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_35),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_289),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_78),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_80),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_119),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_133),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_144),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_100),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_295),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_116),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_285),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_154),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_274),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g462 ( 
.A(n_115),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_322),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_101),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_153),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_94),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_11),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_218),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_260),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_16),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_209),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_291),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_125),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_40),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_203),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_75),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_165),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_189),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_9),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_272),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_25),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_88),
.Y(n_482)
);

CKINVDCx16_ASAP7_75t_R g483 ( 
.A(n_169),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_52),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_37),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_13),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_350),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_334),
.Y(n_488)
);

OA21x2_ASAP7_75t_L g489 ( 
.A1(n_331),
.A2(n_0),
.B(n_1),
.Y(n_489)
);

BUFx12f_ASAP7_75t_L g490 ( 
.A(n_356),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_395),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_344),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_426),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_417),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_417),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_352),
.B(n_0),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_334),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_426),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_449),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_485),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_396),
.B(n_2),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_407),
.B(n_3),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_426),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_425),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_426),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_351),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_361),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_333),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_436),
.B(n_4),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_335),
.B(n_4),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_337),
.B(n_5),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_356),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_371),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_338),
.B(n_5),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_363),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_423),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_368),
.B(n_6),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_386),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_402),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_423),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_430),
.B(n_8),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_485),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_423),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_431),
.Y(n_524)
);

OA21x2_ASAP7_75t_L g525 ( 
.A1(n_349),
.A2(n_12),
.B(n_13),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_439),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_353),
.Y(n_527)
);

CKINVDCx16_ASAP7_75t_R g528 ( 
.A(n_347),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_434),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_418),
.B(n_14),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_442),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_451),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_341),
.B(n_14),
.Y(n_533)
);

BUFx8_ASAP7_75t_L g534 ( 
.A(n_380),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_354),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_466),
.B(n_15),
.Y(n_536)
);

BUFx8_ASAP7_75t_L g537 ( 
.A(n_411),
.Y(n_537)
);

OA21x2_ASAP7_75t_L g538 ( 
.A1(n_357),
.A2(n_15),
.B(n_16),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_467),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_470),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_476),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_474),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_424),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_437),
.Y(n_544)
);

CKINVDCx8_ASAP7_75t_R g545 ( 
.A(n_446),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_360),
.B(n_18),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_479),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_481),
.B(n_482),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_437),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_364),
.B(n_22),
.Y(n_550)
);

CKINVDCx16_ASAP7_75t_R g551 ( 
.A(n_457),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_456),
.B(n_22),
.Y(n_552)
);

BUFx12f_ASAP7_75t_L g553 ( 
.A(n_342),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_365),
.Y(n_554)
);

BUFx2_ASAP7_75t_L g555 ( 
.A(n_377),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_437),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_390),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_488),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_488),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_506),
.Y(n_560)
);

BUFx6f_ASAP7_75t_SL g561 ( 
.A(n_487),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_518),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_557),
.B(n_403),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_513),
.B(n_483),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_513),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_557),
.B(n_403),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_533),
.B(n_348),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_524),
.Y(n_568)
);

BUFx10_ASAP7_75t_L g569 ( 
.A(n_502),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_529),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_532),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_539),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_552),
.B(n_336),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_543),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_497),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_526),
.B(n_341),
.Y(n_576)
);

BUFx4f_ASAP7_75t_L g577 ( 
.A(n_516),
.Y(n_577)
);

OR2x6_ASAP7_75t_L g578 ( 
.A(n_522),
.B(n_420),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_526),
.B(n_413),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_541),
.Y(n_580)
);

NAND2xp33_ASAP7_75t_L g581 ( 
.A(n_510),
.B(n_437),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_547),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_516),
.Y(n_583)
);

NAND3xp33_ASAP7_75t_L g584 ( 
.A(n_530),
.B(n_492),
.C(n_494),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_516),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_520),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_505),
.Y(n_587)
);

INVx1_ASAP7_75t_SL g588 ( 
.A(n_528),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_520),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_487),
.B(n_413),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_520),
.Y(n_591)
);

AO21x2_ASAP7_75t_L g592 ( 
.A1(n_510),
.A2(n_362),
.B(n_332),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_491),
.B(n_415),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_555),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_543),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_553),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_498),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_508),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_523),
.Y(n_599)
);

OR2x2_ASAP7_75t_L g600 ( 
.A(n_492),
.B(n_345),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_552),
.B(n_359),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_523),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_523),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_560),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_594),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_587),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_592),
.B(n_554),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_592),
.B(n_508),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_562),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_574),
.Y(n_610)
);

A2O1A1Ixp33_ASAP7_75t_L g611 ( 
.A1(n_563),
.A2(n_546),
.B(n_509),
.C(n_502),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_L g612 ( 
.A(n_574),
.B(n_511),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_594),
.B(n_551),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_577),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_574),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_569),
.B(n_530),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_569),
.B(n_509),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_558),
.Y(n_618)
);

AND2x6_ASAP7_75t_SL g619 ( 
.A(n_578),
.B(n_546),
.Y(n_619)
);

INVx8_ASAP7_75t_L g620 ( 
.A(n_561),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_595),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_568),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_592),
.B(n_527),
.Y(n_623)
);

AO221x1_ASAP7_75t_L g624 ( 
.A1(n_578),
.A2(n_522),
.B1(n_495),
.B2(n_512),
.C(n_519),
.Y(n_624)
);

NAND2xp33_ASAP7_75t_L g625 ( 
.A(n_595),
.B(n_511),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_569),
.B(n_545),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_570),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_564),
.B(n_504),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_600),
.B(n_512),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_571),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_566),
.B(n_527),
.Y(n_631)
);

NAND2xp33_ASAP7_75t_L g632 ( 
.A(n_584),
.B(n_514),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_559),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_578),
.A2(n_500),
.B1(n_542),
.B2(n_521),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_593),
.B(n_535),
.Y(n_635)
);

NAND2xp33_ASAP7_75t_L g636 ( 
.A(n_572),
.B(n_514),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_578),
.A2(n_496),
.B1(n_501),
.B2(n_358),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_580),
.Y(n_638)
);

BUFx8_ASAP7_75t_L g639 ( 
.A(n_561),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_576),
.B(n_504),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_590),
.B(n_534),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_598),
.B(n_517),
.Y(n_642)
);

BUFx12f_ASAP7_75t_SL g643 ( 
.A(n_596),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_582),
.Y(n_644)
);

BUFx6f_ASAP7_75t_SL g645 ( 
.A(n_565),
.Y(n_645)
);

INVxp67_ASAP7_75t_L g646 ( 
.A(n_600),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_588),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_565),
.B(n_537),
.Y(n_648)
);

AND2x6_ASAP7_75t_SL g649 ( 
.A(n_579),
.B(n_517),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_573),
.B(n_536),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_573),
.A2(n_601),
.B1(n_567),
.B2(n_561),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_575),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_601),
.B(n_537),
.Y(n_653)
);

NOR2xp67_ASAP7_75t_L g654 ( 
.A(n_597),
.B(n_490),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_597),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_581),
.B(n_493),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_575),
.B(n_498),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_604),
.Y(n_658)
);

NAND3xp33_ASAP7_75t_L g659 ( 
.A(n_632),
.B(n_550),
.C(n_340),
.Y(n_659)
);

O2A1O1Ixp33_ASAP7_75t_L g660 ( 
.A1(n_611),
.A2(n_340),
.B(n_519),
.C(n_515),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_616),
.B(n_343),
.Y(n_661)
);

NOR3xp33_ASAP7_75t_L g662 ( 
.A(n_634),
.B(n_398),
.C(n_397),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_631),
.B(n_415),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_631),
.B(n_346),
.Y(n_664)
);

O2A1O1Ixp33_ASAP7_75t_L g665 ( 
.A1(n_612),
.A2(n_515),
.B(n_548),
.C(n_362),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_628),
.B(n_374),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_647),
.Y(n_667)
);

A2O1A1Ixp33_ASAP7_75t_L g668 ( 
.A1(n_635),
.A2(n_332),
.B(n_433),
.C(n_388),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_625),
.A2(n_433),
.B(n_388),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_640),
.B(n_412),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_646),
.B(n_427),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_629),
.B(n_419),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_650),
.B(n_462),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_605),
.B(n_491),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_615),
.A2(n_525),
.B(n_489),
.Y(n_675)
);

AO22x1_ASAP7_75t_L g676 ( 
.A1(n_639),
.A2(n_548),
.B1(n_404),
.B2(n_416),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_610),
.B(n_432),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_609),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_613),
.B(n_454),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_641),
.B(n_401),
.Y(n_680)
);

INVxp67_ASAP7_75t_SL g681 ( 
.A(n_610),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_621),
.B(n_615),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_622),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_L g684 ( 
.A1(n_637),
.A2(n_452),
.B1(n_484),
.B2(n_435),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_653),
.B(n_486),
.Y(n_685)
);

AO21x2_ASAP7_75t_L g686 ( 
.A1(n_608),
.A2(n_623),
.B(n_607),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_SL g687 ( 
.A(n_643),
.B(n_507),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_627),
.B(n_499),
.Y(n_688)
);

O2A1O1Ixp33_ASAP7_75t_L g689 ( 
.A1(n_636),
.A2(n_531),
.B(n_540),
.C(n_503),
.Y(n_689)
);

O2A1O1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_630),
.A2(n_369),
.B(n_373),
.C(n_370),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_651),
.B(n_499),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_626),
.B(n_375),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_654),
.B(n_617),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_638),
.B(n_330),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_L g695 ( 
.A1(n_642),
.A2(n_538),
.B1(n_525),
.B2(n_383),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_606),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_644),
.B(n_339),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_655),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_620),
.B(n_583),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_607),
.B(n_355),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_656),
.Y(n_701)
);

NAND2x1p5_ASAP7_75t_L g702 ( 
.A(n_648),
.B(n_585),
.Y(n_702)
);

A2O1A1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_608),
.A2(n_379),
.B(n_385),
.C(n_384),
.Y(n_703)
);

O2A1O1Ixp33_ASAP7_75t_L g704 ( 
.A1(n_623),
.A2(n_393),
.B(n_394),
.C(n_389),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_649),
.B(n_399),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_619),
.B(n_406),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_656),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_639),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_657),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_618),
.Y(n_710)
);

AOI21x1_ASAP7_75t_L g711 ( 
.A1(n_633),
.A2(n_589),
.B(n_586),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_620),
.B(n_429),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_614),
.B(n_367),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_645),
.B(n_447),
.Y(n_714)
);

INVx11_ASAP7_75t_L g715 ( 
.A(n_645),
.Y(n_715)
);

O2A1O1Ixp33_ASAP7_75t_L g716 ( 
.A1(n_652),
.A2(n_468),
.B(n_469),
.C(n_455),
.Y(n_716)
);

NAND3xp33_ASAP7_75t_L g717 ( 
.A(n_614),
.B(n_473),
.C(n_472),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_624),
.B(n_372),
.Y(n_718)
);

AOI221xp5_ASAP7_75t_L g719 ( 
.A1(n_634),
.A2(n_478),
.B1(n_480),
.B2(n_477),
.C(n_475),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_631),
.B(n_376),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_646),
.B(n_381),
.Y(n_721)
);

A2O1A1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_611),
.A2(n_378),
.B(n_405),
.C(n_366),
.Y(n_722)
);

AOI22x1_ASAP7_75t_L g723 ( 
.A1(n_615),
.A2(n_444),
.B1(n_445),
.B2(n_409),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_612),
.A2(n_599),
.B(n_591),
.Y(n_724)
);

BUFx4f_ASAP7_75t_L g725 ( 
.A(n_620),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_631),
.B(n_382),
.Y(n_726)
);

O2A1O1Ixp33_ASAP7_75t_L g727 ( 
.A1(n_611),
.A2(n_450),
.B(n_603),
.C(n_602),
.Y(n_727)
);

BUFx2_ASAP7_75t_L g728 ( 
.A(n_643),
.Y(n_728)
);

OAI21x1_ASAP7_75t_L g729 ( 
.A1(n_635),
.A2(n_602),
.B(n_471),
.Y(n_729)
);

INVx2_ASAP7_75t_SL g730 ( 
.A(n_647),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_646),
.B(n_387),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_604),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_631),
.B(n_391),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_631),
.B(n_392),
.Y(n_734)
);

OAI21x1_ASAP7_75t_L g735 ( 
.A1(n_635),
.A2(n_471),
.B(n_440),
.Y(n_735)
);

OA22x2_ASAP7_75t_L g736 ( 
.A1(n_634),
.A2(n_408),
.B1(n_410),
.B2(n_400),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_631),
.B(n_414),
.Y(n_737)
);

OAI21xp5_ASAP7_75t_L g738 ( 
.A1(n_632),
.A2(n_422),
.B(n_421),
.Y(n_738)
);

INVxp33_ASAP7_75t_SL g739 ( 
.A(n_605),
.Y(n_739)
);

AND2x6_ASAP7_75t_L g740 ( 
.A(n_651),
.B(n_440),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_634),
.A2(n_471),
.B1(n_440),
.B2(n_556),
.Y(n_741)
);

O2A1O1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_611),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_742)
);

AOI211x1_ASAP7_75t_L g743 ( 
.A1(n_659),
.A2(n_27),
.B(n_24),
.C(n_26),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_658),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_678),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_SL g746 ( 
.A(n_667),
.B(n_428),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_739),
.B(n_438),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_682),
.A2(n_443),
.B(n_441),
.Y(n_748)
);

AOI21xp33_ASAP7_75t_L g749 ( 
.A1(n_671),
.A2(n_453),
.B(n_448),
.Y(n_749)
);

O2A1O1Ixp33_ASAP7_75t_SL g750 ( 
.A1(n_722),
.A2(n_28),
.B(n_26),
.C(n_27),
.Y(n_750)
);

OAI21xp5_ASAP7_75t_L g751 ( 
.A1(n_675),
.A2(n_459),
.B(n_458),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_728),
.B(n_730),
.Y(n_752)
);

NOR4xp25_ASAP7_75t_L g753 ( 
.A(n_660),
.B(n_30),
.C(n_28),
.D(n_29),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_715),
.Y(n_754)
);

OAI21x1_ASAP7_75t_L g755 ( 
.A1(n_729),
.A2(n_471),
.B(n_440),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_681),
.A2(n_726),
.B(n_720),
.Y(n_756)
);

INVxp67_ASAP7_75t_L g757 ( 
.A(n_687),
.Y(n_757)
);

OAI21xp5_ASAP7_75t_L g758 ( 
.A1(n_727),
.A2(n_461),
.B(n_460),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_725),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_664),
.B(n_463),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_674),
.B(n_31),
.Y(n_761)
);

INVx5_ASAP7_75t_L g762 ( 
.A(n_740),
.Y(n_762)
);

AOI21xp33_ASAP7_75t_L g763 ( 
.A1(n_721),
.A2(n_465),
.B(n_464),
.Y(n_763)
);

OAI21x1_ASAP7_75t_L g764 ( 
.A1(n_735),
.A2(n_711),
.B(n_724),
.Y(n_764)
);

AND3x4_ASAP7_75t_L g765 ( 
.A(n_662),
.B(n_33),
.C(n_34),
.Y(n_765)
);

NOR2xp67_ASAP7_75t_L g766 ( 
.A(n_708),
.B(n_105),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_683),
.Y(n_767)
);

AO31x2_ASAP7_75t_L g768 ( 
.A1(n_695),
.A2(n_549),
.A3(n_556),
.B(n_544),
.Y(n_768)
);

AO31x2_ASAP7_75t_L g769 ( 
.A1(n_700),
.A2(n_549),
.A3(n_556),
.B(n_544),
.Y(n_769)
);

INVx1_ASAP7_75t_SL g770 ( 
.A(n_693),
.Y(n_770)
);

NAND2x1p5_ASAP7_75t_L g771 ( 
.A(n_725),
.B(n_549),
.Y(n_771)
);

AO22x2_ASAP7_75t_L g772 ( 
.A1(n_684),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_676),
.Y(n_773)
);

INVx8_ASAP7_75t_L g774 ( 
.A(n_699),
.Y(n_774)
);

A2O1A1Ixp33_ASAP7_75t_L g775 ( 
.A1(n_719),
.A2(n_41),
.B(n_39),
.C(n_40),
.Y(n_775)
);

AO31x2_ASAP7_75t_L g776 ( 
.A1(n_691),
.A2(n_111),
.A3(n_112),
.B(n_110),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_677),
.B(n_39),
.Y(n_777)
);

AND2x2_ASAP7_75t_SL g778 ( 
.A(n_741),
.B(n_41),
.Y(n_778)
);

OAI21xp5_ASAP7_75t_L g779 ( 
.A1(n_659),
.A2(n_114),
.B(n_113),
.Y(n_779)
);

OAI22xp5_ASAP7_75t_L g780 ( 
.A1(n_733),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_780)
);

AO31x2_ASAP7_75t_L g781 ( 
.A1(n_709),
.A2(n_120),
.A3(n_122),
.B(n_117),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_685),
.A2(n_45),
.B1(n_42),
.B2(n_43),
.Y(n_782)
);

AND2x4_ASAP7_75t_L g783 ( 
.A(n_679),
.B(n_45),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_696),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_L g785 ( 
.A1(n_734),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_666),
.B(n_46),
.Y(n_786)
);

OAI22xp5_ASAP7_75t_L g787 ( 
.A1(n_737),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_732),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_670),
.B(n_50),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_698),
.B(n_51),
.Y(n_790)
);

AO31x2_ASAP7_75t_L g791 ( 
.A1(n_668),
.A2(n_663),
.A3(n_707),
.B(n_701),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_731),
.B(n_53),
.Y(n_792)
);

INVx4_ASAP7_75t_L g793 ( 
.A(n_698),
.Y(n_793)
);

OAI21xp5_ASAP7_75t_L g794 ( 
.A1(n_665),
.A2(n_132),
.B(n_130),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_673),
.B(n_54),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_696),
.Y(n_796)
);

OAI21xp5_ASAP7_75t_L g797 ( 
.A1(n_704),
.A2(n_135),
.B(n_134),
.Y(n_797)
);

OAI21x1_ASAP7_75t_L g798 ( 
.A1(n_723),
.A2(n_137),
.B(n_136),
.Y(n_798)
);

INVx4_ASAP7_75t_L g799 ( 
.A(n_702),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_661),
.B(n_56),
.Y(n_800)
);

NOR4xp25_ASAP7_75t_L g801 ( 
.A(n_742),
.B(n_59),
.C(n_57),
.D(n_58),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_714),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_672),
.B(n_713),
.Y(n_803)
);

AO31x2_ASAP7_75t_L g804 ( 
.A1(n_692),
.A2(n_140),
.A3(n_141),
.B(n_138),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_689),
.Y(n_805)
);

A2O1A1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_690),
.A2(n_61),
.B(n_58),
.C(n_59),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_SL g807 ( 
.A1(n_706),
.A2(n_61),
.B(n_62),
.Y(n_807)
);

A2O1A1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_705),
.A2(n_712),
.B(n_697),
.C(n_694),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_710),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_688),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_686),
.B(n_62),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_736),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_812)
);

A2O1A1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_716),
.A2(n_66),
.B(n_64),
.C(n_65),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_717),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_680),
.B(n_66),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_740),
.B(n_67),
.Y(n_816)
);

O2A1O1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_668),
.A2(n_70),
.B(n_68),
.C(n_69),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_L g818 ( 
.A1(n_675),
.A2(n_148),
.B(n_146),
.Y(n_818)
);

O2A1O1Ixp5_ASAP7_75t_L g819 ( 
.A1(n_738),
.A2(n_72),
.B(n_70),
.C(n_71),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_664),
.B(n_71),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_675),
.A2(n_151),
.B(n_150),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_658),
.Y(n_822)
);

A2O1A1Ixp33_ASAP7_75t_L g823 ( 
.A1(n_669),
.A2(n_75),
.B(n_73),
.C(n_74),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_658),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_658),
.Y(n_825)
);

AO31x2_ASAP7_75t_L g826 ( 
.A1(n_703),
.A2(n_156),
.A3(n_158),
.B(n_155),
.Y(n_826)
);

AOI211x1_ASAP7_75t_L g827 ( 
.A1(n_659),
.A2(n_76),
.B(n_77),
.C(n_78),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_728),
.Y(n_828)
);

A2O1A1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_669),
.A2(n_76),
.B(n_79),
.C(n_80),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_728),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_664),
.B(n_79),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_739),
.B(n_81),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_739),
.B(n_81),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_739),
.B(n_82),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_L g835 ( 
.A1(n_675),
.A2(n_162),
.B(n_160),
.Y(n_835)
);

OA21x2_ASAP7_75t_L g836 ( 
.A1(n_735),
.A2(n_166),
.B(n_164),
.Y(n_836)
);

NOR2xp67_ASAP7_75t_L g837 ( 
.A(n_667),
.B(n_167),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_728),
.Y(n_838)
);

BUFx2_ASAP7_75t_L g839 ( 
.A(n_728),
.Y(n_839)
);

NAND3xp33_ASAP7_75t_L g840 ( 
.A(n_671),
.B(n_83),
.C(n_84),
.Y(n_840)
);

AOI221xp5_ASAP7_75t_L g841 ( 
.A1(n_719),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.C(n_87),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_664),
.B(n_85),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_664),
.B(n_87),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_728),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_662),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_845)
);

AO32x2_ASAP7_75t_L g846 ( 
.A1(n_695),
.A2(n_89),
.A3(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_658),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_715),
.Y(n_848)
);

INVx5_ASAP7_75t_L g849 ( 
.A(n_740),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_671),
.B(n_92),
.Y(n_850)
);

OAI22x1_ASAP7_75t_L g851 ( 
.A1(n_671),
.A2(n_93),
.B1(n_95),
.B2(n_97),
.Y(n_851)
);

OAI21x1_ASAP7_75t_SL g852 ( 
.A1(n_669),
.A2(n_93),
.B(n_95),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_669),
.A2(n_98),
.B(n_184),
.C(n_186),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_664),
.B(n_98),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_664),
.B(n_187),
.Y(n_855)
);

NOR2x1_ASAP7_75t_SL g856 ( 
.A(n_701),
.B(n_196),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_664),
.B(n_197),
.Y(n_857)
);

OA21x2_ASAP7_75t_L g858 ( 
.A1(n_735),
.A2(n_198),
.B(n_199),
.Y(n_858)
);

AOI31xp67_ASAP7_75t_L g859 ( 
.A1(n_718),
.A2(n_200),
.A3(n_201),
.B(n_204),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_664),
.B(n_205),
.Y(n_860)
);

A2O1A1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_669),
.A2(n_206),
.B(n_207),
.C(n_210),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_675),
.A2(n_215),
.B(n_216),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_669),
.A2(n_217),
.B(n_219),
.C(n_221),
.Y(n_863)
);

CKINVDCx20_ASAP7_75t_R g864 ( 
.A(n_728),
.Y(n_864)
);

OA21x2_ASAP7_75t_L g865 ( 
.A1(n_735),
.A2(n_222),
.B(n_223),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_664),
.B(n_225),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_802),
.B(n_227),
.Y(n_867)
);

OR2x6_ASAP7_75t_L g868 ( 
.A(n_774),
.B(n_830),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_744),
.Y(n_869)
);

A2O1A1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_808),
.A2(n_228),
.B(n_229),
.C(n_231),
.Y(n_870)
);

OA21x2_ASAP7_75t_L g871 ( 
.A1(n_818),
.A2(n_232),
.B(n_233),
.Y(n_871)
);

BUFx2_ASAP7_75t_R g872 ( 
.A(n_754),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_759),
.Y(n_873)
);

OR2x6_ASAP7_75t_L g874 ( 
.A(n_774),
.B(n_234),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_759),
.B(n_757),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_745),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_784),
.Y(n_877)
);

AND3x2_ASAP7_75t_L g878 ( 
.A(n_746),
.B(n_235),
.C(n_237),
.Y(n_878)
);

CKINVDCx16_ASAP7_75t_R g879 ( 
.A(n_864),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_828),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_767),
.B(n_238),
.Y(n_881)
);

HB1xp67_ASAP7_75t_L g882 ( 
.A(n_839),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_756),
.A2(n_751),
.B(n_821),
.Y(n_883)
);

AOI22x1_ASAP7_75t_L g884 ( 
.A1(n_779),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_884)
);

BUFx2_ASAP7_75t_R g885 ( 
.A(n_848),
.Y(n_885)
);

CKINVDCx11_ASAP7_75t_R g886 ( 
.A(n_830),
.Y(n_886)
);

OA21x2_ASAP7_75t_L g887 ( 
.A1(n_835),
.A2(n_244),
.B(n_245),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_SL g888 ( 
.A(n_778),
.B(n_246),
.Y(n_888)
);

BUFx12f_ASAP7_75t_L g889 ( 
.A(n_773),
.Y(n_889)
);

OA21x2_ASAP7_75t_L g890 ( 
.A1(n_862),
.A2(n_247),
.B(n_248),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_803),
.B(n_249),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_855),
.A2(n_253),
.B(n_254),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_788),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_822),
.Y(n_894)
);

INVx4_ASAP7_75t_L g895 ( 
.A(n_838),
.Y(n_895)
);

OA21x2_ASAP7_75t_L g896 ( 
.A1(n_797),
.A2(n_258),
.B(n_261),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_784),
.B(n_264),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_824),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_752),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_825),
.B(n_265),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_847),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_820),
.A2(n_268),
.B(n_269),
.Y(n_902)
);

NAND2x1p5_ASAP7_75t_L g903 ( 
.A(n_793),
.B(n_270),
.Y(n_903)
);

OR2x6_ASAP7_75t_L g904 ( 
.A(n_844),
.B(n_271),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_796),
.B(n_273),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_791),
.Y(n_906)
);

AO21x2_ASAP7_75t_L g907 ( 
.A1(n_794),
.A2(n_275),
.B(n_277),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_809),
.B(n_279),
.Y(n_908)
);

BUFx2_ASAP7_75t_L g909 ( 
.A(n_783),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_850),
.B(n_280),
.Y(n_910)
);

NOR2x1_ASAP7_75t_SL g911 ( 
.A(n_857),
.B(n_281),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_860),
.A2(n_282),
.B(n_284),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_799),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_866),
.A2(n_290),
.B(n_292),
.Y(n_914)
);

NOR2x1_ASAP7_75t_R g915 ( 
.A(n_832),
.B(n_833),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_805),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_792),
.A2(n_294),
.B(n_296),
.C(n_297),
.Y(n_917)
);

OAI21x1_ASAP7_75t_L g918 ( 
.A1(n_798),
.A2(n_298),
.B(n_300),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_852),
.Y(n_919)
);

OR2x2_ASAP7_75t_L g920 ( 
.A(n_770),
.B(n_301),
.Y(n_920)
);

AOI21x1_ASAP7_75t_L g921 ( 
.A1(n_786),
.A2(n_305),
.B(n_306),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_810),
.Y(n_922)
);

NOR2xp67_ASAP7_75t_L g923 ( 
.A(n_789),
.B(n_307),
.Y(n_923)
);

OA21x2_ASAP7_75t_L g924 ( 
.A1(n_758),
.A2(n_308),
.B(n_309),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_761),
.B(n_310),
.Y(n_925)
);

BUFx12f_ASAP7_75t_L g926 ( 
.A(n_815),
.Y(n_926)
);

AO31x2_ASAP7_75t_L g927 ( 
.A1(n_856),
.A2(n_311),
.A3(n_312),
.B(n_314),
.Y(n_927)
);

OAI21x1_ASAP7_75t_SL g928 ( 
.A1(n_795),
.A2(n_315),
.B(n_316),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_762),
.B(n_849),
.Y(n_929)
);

INVx2_ASAP7_75t_SL g930 ( 
.A(n_790),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_750),
.Y(n_931)
);

AO31x2_ASAP7_75t_L g932 ( 
.A1(n_853),
.A2(n_320),
.A3(n_323),
.B(n_324),
.Y(n_932)
);

AO31x2_ASAP7_75t_L g933 ( 
.A1(n_861),
.A2(n_326),
.A3(n_327),
.B(n_328),
.Y(n_933)
);

INVxp67_ASAP7_75t_L g934 ( 
.A(n_834),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_771),
.Y(n_935)
);

CKINVDCx20_ASAP7_75t_R g936 ( 
.A(n_747),
.Y(n_936)
);

OAI21x1_ASAP7_75t_L g937 ( 
.A1(n_836),
.A2(n_865),
.B(n_858),
.Y(n_937)
);

OAI21x1_ASAP7_75t_L g938 ( 
.A1(n_836),
.A2(n_865),
.B(n_858),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_817),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_L g940 ( 
.A1(n_831),
.A2(n_854),
.B(n_843),
.Y(n_940)
);

BUFx2_ASAP7_75t_R g941 ( 
.A(n_816),
.Y(n_941)
);

NOR2xp67_ASAP7_75t_L g942 ( 
.A(n_842),
.B(n_814),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_819),
.A2(n_760),
.B(n_748),
.Y(n_943)
);

AO31x2_ASAP7_75t_L g944 ( 
.A1(n_863),
.A2(n_851),
.A3(n_829),
.B(n_823),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_749),
.B(n_800),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_762),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_765),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_849),
.B(n_766),
.Y(n_948)
);

AO21x2_ASAP7_75t_L g949 ( 
.A1(n_763),
.A2(n_777),
.B(n_837),
.Y(n_949)
);

NOR2xp67_ASAP7_75t_L g950 ( 
.A(n_840),
.B(n_782),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_772),
.B(n_812),
.Y(n_951)
);

OAI21x1_ASAP7_75t_L g952 ( 
.A1(n_780),
.A2(n_787),
.B(n_785),
.Y(n_952)
);

NAND3xp33_ASAP7_75t_L g953 ( 
.A(n_841),
.B(n_845),
.C(n_775),
.Y(n_953)
);

OAI21x1_ASAP7_75t_L g954 ( 
.A1(n_859),
.A2(n_768),
.B(n_769),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_807),
.B(n_772),
.Y(n_955)
);

OR3x4_ASAP7_75t_SL g956 ( 
.A(n_743),
.B(n_827),
.C(n_846),
.Y(n_956)
);

AOI21x1_ASAP7_75t_L g957 ( 
.A1(n_768),
.A2(n_769),
.B(n_776),
.Y(n_957)
);

INVx1_ASAP7_75t_SL g958 ( 
.A(n_753),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_801),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_813),
.A2(n_806),
.B(n_846),
.Y(n_960)
);

OAI21x1_ASAP7_75t_SL g961 ( 
.A1(n_826),
.A2(n_781),
.B(n_804),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_838),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_744),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_802),
.B(n_739),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_759),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_744),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_828),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_744),
.Y(n_968)
);

NOR2x1_ASAP7_75t_R g969 ( 
.A(n_754),
.B(n_728),
.Y(n_969)
);

NAND3xp33_ASAP7_75t_L g970 ( 
.A(n_782),
.B(n_808),
.C(n_834),
.Y(n_970)
);

OA21x2_ASAP7_75t_L g971 ( 
.A1(n_764),
.A2(n_755),
.B(n_729),
.Y(n_971)
);

NOR2x1_ASAP7_75t_SL g972 ( 
.A(n_811),
.B(n_857),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_759),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_802),
.B(n_646),
.Y(n_974)
);

AO21x2_ASAP7_75t_L g975 ( 
.A1(n_811),
.A2(n_751),
.B(n_794),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_894),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_906),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_898),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_869),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_916),
.B(n_922),
.Y(n_980)
);

AO21x2_ASAP7_75t_L g981 ( 
.A1(n_961),
.A2(n_957),
.B(n_883),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_876),
.Y(n_982)
);

BUFx2_ASAP7_75t_L g983 ( 
.A(n_880),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_974),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_875),
.B(n_868),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_895),
.Y(n_986)
);

BUFx2_ASAP7_75t_L g987 ( 
.A(n_899),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_964),
.B(n_934),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_916),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_886),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_893),
.B(n_901),
.Y(n_991)
);

BUFx2_ASAP7_75t_L g992 ( 
.A(n_895),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_893),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_877),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_901),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_929),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_875),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_963),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_909),
.B(n_947),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_966),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_966),
.Y(n_1001)
);

AO21x2_ASAP7_75t_L g1002 ( 
.A1(n_937),
.A2(n_938),
.B(n_954),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_968),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_968),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_929),
.Y(n_1005)
);

INVx8_ASAP7_75t_L g1006 ( 
.A(n_874),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_877),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_877),
.Y(n_1008)
);

BUFx2_ASAP7_75t_L g1009 ( 
.A(n_882),
.Y(n_1009)
);

BUFx2_ASAP7_75t_L g1010 ( 
.A(n_967),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_962),
.Y(n_1011)
);

BUFx10_ASAP7_75t_L g1012 ( 
.A(n_904),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_959),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_908),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_920),
.Y(n_1015)
);

HB1xp67_ASAP7_75t_L g1016 ( 
.A(n_919),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_874),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_919),
.Y(n_1018)
);

BUFx4f_ASAP7_75t_SL g1019 ( 
.A(n_889),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_951),
.A2(n_953),
.B1(n_888),
.B2(n_970),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_939),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_939),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_930),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_873),
.B(n_965),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_897),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_905),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_955),
.B(n_879),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_905),
.Y(n_1028)
);

BUFx8_ASAP7_75t_L g1029 ( 
.A(n_926),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_946),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_873),
.Y(n_1031)
);

BUFx3_ASAP7_75t_L g1032 ( 
.A(n_965),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_867),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_945),
.B(n_915),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_958),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_904),
.B(n_941),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_973),
.B(n_942),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_946),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_881),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_936),
.B(n_913),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_931),
.Y(n_1041)
);

AO21x2_ASAP7_75t_L g1042 ( 
.A1(n_975),
.A2(n_972),
.B(n_940),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_900),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_948),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_913),
.B(n_935),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_931),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_891),
.Y(n_1047)
);

AND2x4_ASAP7_75t_SL g1048 ( 
.A(n_935),
.B(n_872),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_950),
.B(n_925),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_903),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_885),
.B(n_949),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_952),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_944),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_944),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_878),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_944),
.Y(n_1056)
);

INVx2_ASAP7_75t_SL g1057 ( 
.A(n_969),
.Y(n_1057)
);

OA21x2_ASAP7_75t_L g1058 ( 
.A1(n_943),
.A2(n_960),
.B(n_918),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_923),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_910),
.B(n_911),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_911),
.Y(n_1061)
);

HB1xp67_ASAP7_75t_L g1062 ( 
.A(n_971),
.Y(n_1062)
);

OR2x6_ASAP7_75t_L g1063 ( 
.A(n_902),
.B(n_892),
.Y(n_1063)
);

INVxp67_ASAP7_75t_L g1064 ( 
.A(n_928),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_907),
.B(n_870),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_917),
.B(n_927),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_921),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_977),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_993),
.B(n_932),
.Y(n_1069)
);

AOI22xp33_ASAP7_75t_L g1070 ( 
.A1(n_1020),
.A2(n_896),
.B1(n_924),
.B2(n_884),
.Y(n_1070)
);

NOR2x1_ASAP7_75t_L g1071 ( 
.A(n_1049),
.B(n_914),
.Y(n_1071)
);

OAI221xp5_ASAP7_75t_L g1072 ( 
.A1(n_1049),
.A2(n_884),
.B1(n_890),
.B2(n_871),
.C(n_887),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_984),
.B(n_932),
.Y(n_1073)
);

NOR2x1_ASAP7_75t_L g1074 ( 
.A(n_1011),
.B(n_912),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_976),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_988),
.B(n_933),
.Y(n_1076)
);

BUFx3_ASAP7_75t_L g1077 ( 
.A(n_985),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_1041),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_1041),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_983),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_993),
.B(n_933),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_978),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_991),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_989),
.Y(n_1084)
);

HB1xp67_ASAP7_75t_L g1085 ( 
.A(n_989),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_1053),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_992),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_979),
.B(n_956),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_1009),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_982),
.B(n_971),
.Y(n_1090)
);

OR2x2_ASAP7_75t_L g1091 ( 
.A(n_1010),
.B(n_1035),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_995),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_998),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1000),
.Y(n_1094)
);

INVx5_ASAP7_75t_L g1095 ( 
.A(n_1006),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1034),
.B(n_1020),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1001),
.Y(n_1097)
);

INVx5_ASAP7_75t_L g1098 ( 
.A(n_1006),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_1006),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_1027),
.B(n_999),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_L g1101 ( 
.A1(n_1047),
.A2(n_1036),
.B1(n_1034),
.B2(n_1015),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_1040),
.B(n_1048),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1003),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_1048),
.B(n_997),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_1004),
.B(n_1021),
.Y(n_1105)
);

NOR2x1_ASAP7_75t_L g1106 ( 
.A(n_1031),
.B(n_1032),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_1022),
.B(n_1054),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1056),
.B(n_1013),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_980),
.B(n_1046),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_980),
.B(n_1016),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_1032),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1033),
.B(n_1024),
.Y(n_1112)
);

INVx4_ASAP7_75t_L g1113 ( 
.A(n_1030),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_987),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1037),
.B(n_1007),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1008),
.B(n_1012),
.Y(n_1116)
);

INVxp67_ASAP7_75t_L g1117 ( 
.A(n_1023),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1018),
.B(n_1042),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1042),
.B(n_1052),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_1017),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_990),
.B(n_994),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_990),
.B(n_1051),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_1110),
.B(n_1076),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_1095),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_1078),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_1091),
.B(n_986),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1100),
.B(n_1014),
.Y(n_1127)
);

OR2x2_ASAP7_75t_L g1128 ( 
.A(n_1089),
.B(n_1025),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1068),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1082),
.Y(n_1130)
);

HB1xp67_ASAP7_75t_L g1131 ( 
.A(n_1078),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1110),
.B(n_1062),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1088),
.B(n_1062),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1092),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_1088),
.B(n_981),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_1107),
.B(n_1061),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1109),
.B(n_981),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1109),
.B(n_1043),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1093),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_1087),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1083),
.B(n_1039),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1105),
.B(n_1028),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1094),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_1112),
.B(n_1026),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1080),
.B(n_996),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1097),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1090),
.B(n_1002),
.Y(n_1147)
);

INVx1_ASAP7_75t_SL g1148 ( 
.A(n_1114),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1103),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1090),
.B(n_1002),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1096),
.B(n_1005),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1084),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1118),
.B(n_1069),
.Y(n_1153)
);

OR2x2_ASAP7_75t_L g1154 ( 
.A(n_1084),
.B(n_1045),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1085),
.B(n_1060),
.Y(n_1155)
);

NAND2x1_ASAP7_75t_L g1156 ( 
.A(n_1074),
.B(n_1038),
.Y(n_1156)
);

INVxp67_ASAP7_75t_SL g1157 ( 
.A(n_1079),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1085),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_1087),
.Y(n_1159)
);

INVxp67_ASAP7_75t_SL g1160 ( 
.A(n_1079),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1075),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1118),
.B(n_1058),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1115),
.B(n_1038),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1122),
.B(n_1044),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1111),
.B(n_1050),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1069),
.B(n_1081),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1101),
.A2(n_1055),
.B1(n_1059),
.B2(n_1063),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1117),
.B(n_1064),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1152),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_1136),
.B(n_1108),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1158),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1168),
.B(n_1120),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1125),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1123),
.B(n_1102),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1123),
.B(n_1121),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1125),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1148),
.B(n_1019),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1131),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1131),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1140),
.B(n_1073),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1133),
.B(n_1135),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1134),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1139),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_1159),
.B(n_1113),
.Y(n_1184)
);

HB1xp67_ASAP7_75t_L g1185 ( 
.A(n_1157),
.Y(n_1185)
);

NOR2x1p5_ASAP7_75t_L g1186 ( 
.A(n_1151),
.B(n_1155),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1160),
.B(n_1081),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1136),
.B(n_1095),
.Y(n_1188)
);

O2A1O1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_1167),
.A2(n_1072),
.B(n_1063),
.C(n_1065),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1161),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1136),
.B(n_1098),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1143),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_1159),
.B(n_1098),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1129),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1146),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1137),
.B(n_1119),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1135),
.B(n_1104),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_1153),
.B(n_1098),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1149),
.Y(n_1199)
);

OR2x2_ASAP7_75t_L g1200 ( 
.A(n_1153),
.B(n_1086),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1132),
.B(n_1099),
.Y(n_1201)
);

INVx2_ASAP7_75t_SL g1202 ( 
.A(n_1126),
.Y(n_1202)
);

OAI21xp33_ASAP7_75t_L g1203 ( 
.A1(n_1173),
.A2(n_1178),
.B(n_1176),
.Y(n_1203)
);

INVx2_ASAP7_75t_SL g1204 ( 
.A(n_1185),
.Y(n_1204)
);

OR2x2_ASAP7_75t_L g1205 ( 
.A(n_1200),
.B(n_1132),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1179),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1181),
.B(n_1137),
.Y(n_1207)
);

INVxp67_ASAP7_75t_SL g1208 ( 
.A(n_1185),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1186),
.B(n_1138),
.Y(n_1209)
);

INVxp67_ASAP7_75t_L g1210 ( 
.A(n_1172),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1182),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1183),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1197),
.B(n_1147),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1180),
.B(n_1147),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1175),
.B(n_1150),
.Y(n_1215)
);

INVxp67_ASAP7_75t_SL g1216 ( 
.A(n_1187),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1174),
.B(n_1166),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1192),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1194),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1170),
.B(n_1150),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1172),
.B(n_1154),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_SL g1222 ( 
.A1(n_1189),
.A2(n_1191),
.B(n_1188),
.Y(n_1222)
);

OAI21xp33_ASAP7_75t_SL g1223 ( 
.A1(n_1193),
.A2(n_1145),
.B(n_1165),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1195),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1199),
.Y(n_1225)
);

OR2x6_ASAP7_75t_L g1226 ( 
.A(n_1189),
.B(n_1124),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1190),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1206),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1215),
.B(n_1201),
.Y(n_1229)
);

AOI32xp33_ASAP7_75t_L g1230 ( 
.A1(n_1223),
.A2(n_1167),
.A3(n_1101),
.B1(n_1066),
.B2(n_1170),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1222),
.A2(n_1070),
.B(n_1169),
.Y(n_1231)
);

OR2x6_ASAP7_75t_L g1232 ( 
.A(n_1222),
.B(n_1188),
.Y(n_1232)
);

AOI222xp33_ASAP7_75t_L g1233 ( 
.A1(n_1216),
.A2(n_1196),
.B1(n_1070),
.B2(n_1142),
.C1(n_1162),
.C2(n_1144),
.Y(n_1233)
);

OAI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1226),
.A2(n_1209),
.B1(n_1063),
.B2(n_1196),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1219),
.Y(n_1235)
);

AOI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1226),
.A2(n_1162),
.B1(n_1071),
.B2(n_1164),
.Y(n_1236)
);

OAI32xp33_ASAP7_75t_SL g1237 ( 
.A1(n_1210),
.A2(n_1177),
.A3(n_1202),
.B1(n_1171),
.B2(n_1019),
.Y(n_1237)
);

NAND2xp33_ASAP7_75t_L g1238 ( 
.A(n_1221),
.B(n_1187),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1220),
.B(n_1198),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1204),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1215),
.B(n_1198),
.Y(n_1241)
);

INVx1_ASAP7_75t_SL g1242 ( 
.A(n_1217),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1211),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1212),
.Y(n_1244)
);

AOI221xp5_ASAP7_75t_L g1245 ( 
.A1(n_1230),
.A2(n_1203),
.B1(n_1225),
.B2(n_1224),
.C(n_1218),
.Y(n_1245)
);

AOI32xp33_ASAP7_75t_L g1246 ( 
.A1(n_1238),
.A2(n_1214),
.A3(n_1220),
.B1(n_1207),
.B2(n_1213),
.Y(n_1246)
);

OAI21xp33_ASAP7_75t_L g1247 ( 
.A1(n_1231),
.A2(n_1208),
.B(n_1204),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_1242),
.B(n_1205),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1233),
.A2(n_1226),
.B(n_1227),
.Y(n_1249)
);

NOR3xp33_ASAP7_75t_L g1250 ( 
.A(n_1234),
.B(n_1156),
.C(n_1184),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1228),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1245),
.B(n_1243),
.Y(n_1252)
);

OAI211xp5_ASAP7_75t_L g1253 ( 
.A1(n_1247),
.A2(n_1237),
.B(n_1240),
.C(n_1236),
.Y(n_1253)
);

NOR2xp67_ASAP7_75t_L g1254 ( 
.A(n_1249),
.B(n_1239),
.Y(n_1254)
);

AOI21xp33_ASAP7_75t_L g1255 ( 
.A1(n_1251),
.A2(n_1232),
.B(n_1228),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1248),
.Y(n_1256)
);

NOR2x1_ASAP7_75t_L g1257 ( 
.A(n_1253),
.B(n_1232),
.Y(n_1257)
);

AOI21xp33_ASAP7_75t_L g1258 ( 
.A1(n_1252),
.A2(n_1244),
.B(n_1141),
.Y(n_1258)
);

NAND3xp33_ASAP7_75t_L g1259 ( 
.A(n_1256),
.B(n_1250),
.C(n_1246),
.Y(n_1259)
);

NOR2x1_ASAP7_75t_L g1260 ( 
.A(n_1254),
.B(n_1239),
.Y(n_1260)
);

A2O1A1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_1255),
.A2(n_1213),
.B(n_1214),
.C(n_1207),
.Y(n_1261)
);

INVxp67_ASAP7_75t_L g1262 ( 
.A(n_1257),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1258),
.B(n_1259),
.Y(n_1263)
);

NAND3x1_ASAP7_75t_L g1264 ( 
.A(n_1260),
.B(n_1241),
.C(n_1229),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1263),
.B(n_1261),
.Y(n_1265)
);

NAND3x2_ASAP7_75t_L g1266 ( 
.A(n_1264),
.B(n_1128),
.C(n_1130),
.Y(n_1266)
);

NAND2x1_ASAP7_75t_L g1267 ( 
.A(n_1265),
.B(n_1262),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1267),
.B(n_1127),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_SL g1269 ( 
.A1(n_1268),
.A2(n_1057),
.B1(n_1266),
.B2(n_1029),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1269),
.A2(n_1029),
.B(n_1106),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1270),
.B(n_1163),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1271),
.A2(n_1064),
.B(n_1184),
.Y(n_1272)
);

OR2x6_ASAP7_75t_L g1273 ( 
.A(n_1272),
.B(n_1077),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1273),
.A2(n_1116),
.B1(n_1067),
.B2(n_1235),
.Y(n_1274)
);


endmodule