module fake_aes_7817_n_36 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_36);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_36;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_13;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
HB1xp67_ASAP7_75t_L g11 ( .A(n_2), .Y(n_11) );
BUFx3_ASAP7_75t_L g12 ( .A(n_6), .Y(n_12) );
NOR2xp33_ASAP7_75t_L g13 ( .A(n_0), .B(n_2), .Y(n_13) );
AOI21x1_ASAP7_75t_L g14 ( .A1(n_3), .A2(n_10), .B(n_8), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_6), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_3), .Y(n_16) );
INVx2_ASAP7_75t_SL g17 ( .A(n_10), .Y(n_17) );
OAI22xp5_ASAP7_75t_L g18 ( .A1(n_11), .A2(n_0), .B1(n_1), .B2(n_4), .Y(n_18) );
AOI21xp5_ASAP7_75t_L g19 ( .A1(n_17), .A2(n_0), .B(n_1), .Y(n_19) );
OAI21x1_ASAP7_75t_L g20 ( .A1(n_15), .A2(n_1), .B(n_4), .Y(n_20) );
A2O1A1Ixp33_ASAP7_75t_L g21 ( .A1(n_12), .A2(n_5), .B(n_7), .C(n_8), .Y(n_21) );
OAI22x1_ASAP7_75t_L g22 ( .A1(n_14), .A2(n_5), .B1(n_7), .B2(n_9), .Y(n_22) );
AOI22xp33_ASAP7_75t_L g23 ( .A1(n_19), .A2(n_11), .B1(n_16), .B2(n_12), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_20), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_19), .B(n_17), .Y(n_25) );
OR2x2_ASAP7_75t_L g26 ( .A(n_23), .B(n_18), .Y(n_26) );
AND2x2_ASAP7_75t_L g27 ( .A(n_24), .B(n_12), .Y(n_27) );
AND2x2_ASAP7_75t_L g28 ( .A(n_24), .B(n_12), .Y(n_28) );
INVx2_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
INVx1_ASAP7_75t_SL g30 ( .A(n_27), .Y(n_30) );
AO21x1_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_28), .B(n_25), .Y(n_31) );
AOI21xp5_ASAP7_75t_L g32 ( .A1(n_29), .A2(n_26), .B(n_22), .Y(n_32) );
NAND2xp5_ASAP7_75t_L g33 ( .A(n_31), .B(n_30), .Y(n_33) );
O2A1O1Ixp33_ASAP7_75t_L g34 ( .A1(n_32), .A2(n_21), .B(n_17), .C(n_16), .Y(n_34) );
CKINVDCx16_ASAP7_75t_R g35 ( .A(n_33), .Y(n_35) );
OAI22xp5_ASAP7_75t_L g36 ( .A1(n_35), .A2(n_33), .B1(n_34), .B2(n_13), .Y(n_36) );
endmodule