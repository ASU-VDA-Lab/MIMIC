module fake_jpeg_1408_n_407 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_407);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_407;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_SL g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_10),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_16),
.B(n_13),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_45),
.B(n_56),
.Y(n_108)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_46),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_47),
.B(n_53),
.Y(n_102)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_49),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_51),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_52),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_54),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_55),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_22),
.B(n_13),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g116 ( 
.A(n_57),
.Y(n_116)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_63),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_13),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_77),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_22),
.B(n_12),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_71),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_67),
.Y(n_149)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_70),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_38),
.B(n_12),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_76),
.Y(n_145)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_81),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g128 ( 
.A(n_79),
.B(n_80),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_83),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_39),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_84),
.B(n_85),
.Y(n_132)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_86),
.B(n_87),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_38),
.B(n_0),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_39),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_89),
.Y(n_118)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_39),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_90),
.B(n_92),
.Y(n_136)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_93),
.Y(n_115)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_19),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_94),
.B(n_32),
.Y(n_140)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_95),
.B(n_35),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_18),
.B(n_0),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_96),
.B(n_42),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_64),
.A2(n_28),
.B1(n_36),
.B2(n_29),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_97),
.A2(n_120),
.B1(n_122),
.B2(n_152),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_94),
.A2(n_42),
.B1(n_26),
.B2(n_24),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_99),
.Y(n_171)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_49),
.B(n_42),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_101),
.B(n_104),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_103),
.B(n_6),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_58),
.B(n_24),
.C(n_26),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_73),
.A2(n_29),
.B1(n_36),
.B2(n_40),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_SL g121 ( 
.A(n_49),
.Y(n_121)
);

INVx11_ASAP7_75t_L g195 ( 
.A(n_121),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_50),
.A2(n_26),
.B1(n_40),
.B2(n_32),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_61),
.A2(n_41),
.B1(n_18),
.B2(n_33),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_125),
.Y(n_190)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_85),
.A2(n_36),
.B1(n_41),
.B2(n_19),
.Y(n_126)
);

AND2x4_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_150),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_48),
.A2(n_41),
.B1(n_35),
.B2(n_34),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_131),
.A2(n_151),
.B1(n_93),
.B2(n_7),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_137),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_70),
.B(n_34),
.C(n_33),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_138),
.B(n_144),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_80),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_91),
.B(n_30),
.C(n_21),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_81),
.B(n_30),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_133),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_51),
.B(n_19),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_147),
.Y(n_177)
);

OA22x2_ASAP7_75t_L g150 ( 
.A1(n_54),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_62),
.A2(n_21),
.B1(n_3),
.B2(n_4),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_55),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_155),
.B(n_161),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_156),
.Y(n_206)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_98),
.Y(n_158)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_160),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_113),
.Y(n_162)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_162),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_114),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_163),
.B(n_170),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_66),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_164),
.B(n_174),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_113),
.Y(n_165)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_106),
.B(n_68),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_166),
.B(n_173),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_118),
.Y(n_170)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_112),
.B(n_102),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_63),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_108),
.B(n_67),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_178),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_86),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_192),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_117),
.B(n_60),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_179),
.Y(n_226)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_180),
.B(n_181),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_57),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_122),
.A2(n_92),
.B1(n_69),
.B2(n_79),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_183),
.A2(n_188),
.B1(n_191),
.B2(n_132),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_98),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_184),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_135),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_185),
.Y(n_205)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_98),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_186),
.B(n_187),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_L g188 ( 
.A1(n_126),
.A2(n_75),
.B1(n_74),
.B2(n_95),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_189),
.A2(n_150),
.B1(n_119),
.B2(n_109),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_126),
.A2(n_115),
.B1(n_150),
.B2(n_128),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_101),
.B(n_147),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_100),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_193),
.Y(n_201)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_143),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_194),
.Y(n_223)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_105),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_196),
.A2(n_133),
.B1(n_100),
.B2(n_119),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_124),
.B(n_44),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_198),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_101),
.B(n_147),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_145),
.B(n_6),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_7),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_174),
.A2(n_126),
.B1(n_132),
.B2(n_115),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_200),
.B(n_219),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_159),
.A2(n_127),
.B1(n_111),
.B2(n_148),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_210),
.A2(n_216),
.B1(n_184),
.B2(n_188),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_198),
.A2(n_128),
.B(n_150),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_213),
.A2(n_157),
.B(n_155),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_175),
.A2(n_132),
.B1(n_148),
.B2(n_111),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_104),
.C(n_123),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_182),
.C(n_164),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_225),
.B(n_229),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_227),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_177),
.A2(n_149),
.B1(n_142),
.B2(n_139),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_228),
.A2(n_231),
.B1(n_195),
.B2(n_171),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_169),
.A2(n_149),
.B1(n_142),
.B2(n_139),
.Y(n_231)
);

AOI32xp33_ASAP7_75t_L g232 ( 
.A1(n_192),
.A2(n_107),
.A3(n_129),
.B1(n_153),
.B2(n_110),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_182),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_233),
.A2(n_249),
.B1(n_252),
.B2(n_200),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_234),
.B(n_240),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_209),
.Y(n_235)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_235),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_236),
.B(n_247),
.C(n_203),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_237),
.Y(n_279)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_238),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_167),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_241),
.A2(n_158),
.B(n_223),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_204),
.B(n_169),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_242),
.B(n_243),
.Y(n_263)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_245),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_163),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_204),
.C(n_224),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_231),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_250),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_216),
.A2(n_157),
.B1(n_190),
.B2(n_189),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_210),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_213),
.A2(n_157),
.B1(n_159),
.B2(n_190),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_207),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_253),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_208),
.B(n_170),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_254),
.A2(n_256),
.B(n_202),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_255),
.A2(n_257),
.B1(n_223),
.B2(n_205),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_224),
.A2(n_157),
.B(n_171),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_218),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_211),
.B(n_176),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_258),
.B(n_211),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_260),
.B(n_262),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_214),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_214),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_266),
.C(n_268),
.Y(n_289)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_265),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_217),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_248),
.A2(n_227),
.B1(n_217),
.B2(n_202),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_267),
.A2(n_249),
.B1(n_233),
.B2(n_246),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_236),
.B(n_203),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_269),
.A2(n_278),
.B(n_282),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_272),
.B(n_273),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_236),
.B(n_221),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_207),
.C(n_186),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_281),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_237),
.B(n_221),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_277),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_252),
.A2(n_219),
.B1(n_183),
.B2(n_232),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_280),
.A2(n_255),
.B1(n_225),
.B2(n_243),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_253),
.B(n_256),
.C(n_241),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_278),
.A2(n_251),
.B1(n_246),
.B2(n_244),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_283),
.A2(n_284),
.B1(n_299),
.B2(n_302),
.Y(n_309)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_275),
.Y(n_288)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_288),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_270),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_290),
.B(n_295),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_263),
.B(n_254),
.Y(n_292)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_292),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_261),
.B(n_245),
.Y(n_293)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_293),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_261),
.B(n_234),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_296),
.Y(n_317)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_271),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_298),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_267),
.A2(n_250),
.B1(n_240),
.B2(n_239),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_300),
.A2(n_301),
.B1(n_230),
.B2(n_201),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_280),
.A2(n_279),
.B1(n_269),
.B2(n_282),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_281),
.A2(n_235),
.B1(n_205),
.B2(n_238),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_260),
.B(n_235),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_303),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_259),
.B(n_235),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_304),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_284),
.A2(n_266),
.B1(n_277),
.B2(n_262),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_305),
.A2(n_313),
.B1(n_297),
.B2(n_303),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_268),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_306),
.B(n_311),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_272),
.C(n_289),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_307),
.B(n_318),
.C(n_291),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_289),
.B(n_264),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_274),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_312),
.B(n_291),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_284),
.A2(n_273),
.B1(n_276),
.B2(n_257),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_298),
.A2(n_276),
.B1(n_209),
.B2(n_230),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_315),
.A2(n_319),
.B1(n_322),
.B2(n_287),
.Y(n_332)
);

A2O1A1O1Ixp25_ASAP7_75t_L g316 ( 
.A1(n_295),
.A2(n_226),
.B(n_215),
.C(n_218),
.D(n_129),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_316),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_294),
.B(n_226),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_301),
.A2(n_215),
.B1(n_201),
.B2(n_185),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_285),
.A2(n_206),
.B(n_196),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_324),
.A2(n_296),
.B(n_288),
.Y(n_344)
);

NAND3xp33_ASAP7_75t_L g325 ( 
.A(n_292),
.B(n_206),
.C(n_109),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_325),
.B(n_206),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_293),
.Y(n_328)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_328),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_309),
.A2(n_283),
.B1(n_300),
.B2(n_302),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_330),
.A2(n_332),
.B1(n_341),
.B2(n_344),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_314),
.Y(n_331)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_331),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_333),
.B(n_334),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_286),
.C(n_291),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_339),
.C(n_305),
.Y(n_346)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_326),
.Y(n_336)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_336),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_323),
.A2(n_299),
.B1(n_287),
.B2(n_304),
.Y(n_337)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_337),
.Y(n_355)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_323),
.Y(n_338)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_338),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_306),
.B(n_311),
.C(n_318),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_319),
.A2(n_285),
.B1(n_297),
.B2(n_286),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_340),
.B(n_345),
.Y(n_349)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_308),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_342),
.B(n_320),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_343),
.B(n_316),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_320),
.B(n_297),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_346),
.B(n_352),
.Y(n_371)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_351),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_329),
.B(n_313),
.C(n_324),
.Y(n_352)
);

O2A1O1Ixp33_ASAP7_75t_L g356 ( 
.A1(n_331),
.A2(n_317),
.B(n_322),
.C(n_310),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_356),
.A2(n_344),
.B(n_337),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_345),
.B(n_172),
.Y(n_358)
);

NOR2xp67_ASAP7_75t_L g364 ( 
.A(n_358),
.B(n_359),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_350),
.B(n_329),
.C(n_335),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_361),
.B(n_368),
.C(n_370),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_349),
.A2(n_328),
.B(n_330),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_362),
.B(n_369),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_363),
.A2(n_347),
.B1(n_354),
.B2(n_355),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_349),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_365),
.B(n_366),
.Y(n_373)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_356),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_348),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_367),
.B(n_347),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_350),
.B(n_339),
.C(n_333),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_327),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_346),
.B(n_340),
.C(n_334),
.Y(n_370)
);

A2O1A1Ixp33_ASAP7_75t_SL g383 ( 
.A1(n_372),
.A2(n_369),
.B(n_365),
.C(n_370),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_361),
.B(n_352),
.C(n_355),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_375),
.B(n_376),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_360),
.B(n_353),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_377),
.B(n_378),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_363),
.A2(n_357),
.B1(n_353),
.B2(n_165),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_362),
.B(n_162),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_380),
.B(n_381),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_364),
.B(n_162),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_383),
.B(n_384),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_374),
.B(n_371),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_373),
.A2(n_368),
.B1(n_193),
.B2(n_135),
.Y(n_386)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_386),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_374),
.B(n_180),
.C(n_168),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_388),
.B(n_156),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_375),
.A2(n_130),
.B(n_110),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_389),
.A2(n_379),
.B(n_372),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_385),
.B(n_379),
.Y(n_392)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_392),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_393),
.B(n_394),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_383),
.A2(n_179),
.B(n_116),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_395),
.A2(n_382),
.B(n_107),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_391),
.B(n_387),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_396),
.A2(n_8),
.B(n_9),
.Y(n_402)
);

O2A1O1Ixp33_ASAP7_75t_SL g400 ( 
.A1(n_399),
.A2(n_390),
.B(n_156),
.C(n_195),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_400),
.A2(n_401),
.B(n_11),
.Y(n_404)
);

AOI321xp33_ASAP7_75t_L g401 ( 
.A1(n_398),
.A2(n_156),
.A3(n_194),
.B1(n_160),
.B2(n_105),
.C(n_116),
.Y(n_401)
);

OAI21x1_ASAP7_75t_L g403 ( 
.A1(n_402),
.A2(n_397),
.B(n_10),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_403),
.A2(n_404),
.B(n_9),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_405),
.A2(n_9),
.B(n_10),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_406),
.A2(n_11),
.B(n_403),
.Y(n_407)
);


endmodule