module real_jpeg_14122_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g80 ( 
.A(n_2),
.Y(n_80)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_3),
.A2(n_26),
.B(n_32),
.C(n_72),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_3),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_73),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_3),
.B(n_107),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_3),
.B(n_27),
.Y(n_141)
);

AOI21xp33_ASAP7_75t_SL g156 ( 
.A1(n_3),
.A2(n_27),
.B(n_141),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_3),
.B(n_60),
.C(n_78),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_3),
.A2(n_45),
.B1(n_49),
.B2(n_73),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_3),
.A2(n_59),
.B1(n_63),
.B2(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_3),
.B(n_55),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_39),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_4),
.A2(n_39),
.B1(n_45),
.B2(n_49),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_4),
.A2(n_39),
.B1(n_60),
.B2(n_67),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_7),
.A2(n_60),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_7),
.A2(n_45),
.B1(n_49),
.B2(n_66),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_8),
.A2(n_60),
.B1(n_67),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_8),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_10),
.A2(n_45),
.B1(n_49),
.B2(n_54),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_10),
.A2(n_54),
.B1(n_60),
.B2(n_67),
.Y(n_145)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_13),
.A2(n_45),
.B1(n_49),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_13),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_13),
.A2(n_60),
.B1(n_67),
.B2(n_84),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_37),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_14),
.A2(n_37),
.B1(n_45),
.B2(n_49),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_14),
.A2(n_37),
.B1(n_60),
.B2(n_67),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_15),
.A2(n_42),
.B1(n_45),
.B2(n_49),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_15),
.A2(n_42),
.B1(n_60),
.B2(n_67),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_124),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_122),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_108),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_20),
.B(n_108),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_74),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_56),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_36),
.B2(n_38),
.Y(n_23)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_25),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_26),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_26),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_27),
.A2(n_28),
.B1(n_47),
.B2(n_48),
.Y(n_50)
);

OAI21xp33_ASAP7_75t_L g72 ( 
.A1(n_27),
.A2(n_30),
.B(n_73),
.Y(n_72)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND3xp33_ASAP7_75t_SL g142 ( 
.A(n_28),
.B(n_47),
.C(n_49),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_36),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_43),
.B(n_51),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_41),
.A2(n_43),
.B1(n_44),
.B2(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_43),
.A2(n_44),
.B1(n_102),
.B2(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_43),
.A2(n_44),
.B1(n_121),
.B2(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_50),
.Y(n_43)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_44)
);

INVx5_ASAP7_75t_SL g49 ( 
.A(n_45),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_45),
.A2(n_49),
.B1(n_78),
.B2(n_79),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_45),
.A2(n_48),
.B(n_140),
.C(n_142),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_45),
.B(n_165),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_70),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_57),
.A2(n_70),
.B1(n_71),
.B2(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_64),
.B1(n_65),
.B2(n_68),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_58),
.A2(n_90),
.B(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_58),
.A2(n_64),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_59),
.A2(n_88),
.B(n_89),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_59),
.B(n_91),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_59),
.A2(n_63),
.B1(n_171),
.B2(n_179),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_59),
.A2(n_173),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_60),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_60),
.A2(n_67),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

BUFx4f_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_63),
.B(n_73),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_64),
.A2(n_65),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_64),
.B(n_145),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_67),
.B(n_177),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_73),
.B(n_77),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_92),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_87),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_81),
.B(n_82),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_SL g78 ( 
.A(n_79),
.Y(n_78)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_85),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_83),
.B(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_85),
.A2(n_99),
.B1(n_135),
.B2(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_85),
.A2(n_99),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_85),
.A2(n_99),
.B1(n_158),
.B2(n_168),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_100),
.C(n_103),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_94),
.B1(n_100),
.B2(n_101),
.Y(n_110)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_96),
.B(n_98),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_95),
.A2(n_134),
.B(n_136),
.Y(n_133)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_99),
.Y(n_136)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_103),
.B(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.C(n_114),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_112),
.B1(n_114),
.B2(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.C(n_120),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_132)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_120),
.B(n_132),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_203),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_146),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_127),
.B(n_130),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.C(n_137),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_133),
.A2(n_137),
.B1(n_138),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_139),
.A2(n_143),
.B1(n_144),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_159),
.B(n_202),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_148),
.B(n_151),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.C(n_157),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_154),
.A2(n_155),
.B1(n_157),
.B2(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_196),
.B(n_201),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_185),
.B(n_195),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_174),
.B(n_184),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_169),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_169),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_166),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_180),
.B(n_183),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_181),
.B(n_182),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_187),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_191),
.C(n_194),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_193),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_200),
.Y(n_201)
);


endmodule