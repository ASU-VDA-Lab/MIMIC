module fake_jpeg_23016_n_265 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_38),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_41),
.B(n_44),
.Y(n_72)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_42),
.A2(n_31),
.B1(n_30),
.B2(n_18),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_1),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_45),
.B(n_16),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_26),
.B(n_1),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_16),
.Y(n_53)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_32),
.Y(n_57)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_50),
.Y(n_89)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_48),
.A2(n_22),
.B1(n_30),
.B2(n_18),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_51),
.A2(n_27),
.B1(n_31),
.B2(n_25),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_52),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_53),
.B(n_57),
.Y(n_103)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_58),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_67),
.Y(n_96)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_63),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_29),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_61),
.B(n_65),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_41),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_SL g64 ( 
.A(n_48),
.B(n_2),
.Y(n_64)
);

OR2x2_ASAP7_75t_SL g115 ( 
.A(n_64),
.B(n_34),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_29),
.Y(n_65)
);

CKINVDCx12_ASAP7_75t_R g66 ( 
.A(n_37),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_66),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_47),
.B(n_23),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_71),
.Y(n_105)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_32),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_73),
.B(n_83),
.Y(n_112)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_78),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_42),
.B(n_35),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_77),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_42),
.B(n_35),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_36),
.A2(n_30),
.B1(n_22),
.B2(n_18),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_81),
.B1(n_31),
.B2(n_28),
.Y(n_94)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_84),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_26),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_87),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_46),
.B(n_24),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_92),
.Y(n_122)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_93),
.B(n_105),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_94),
.A2(n_104),
.B1(n_76),
.B2(n_69),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_34),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_85),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_64),
.B(n_17),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_25),
.C(n_76),
.Y(n_138)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_102),
.Y(n_123)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_109),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

HAxp5_ASAP7_75t_SL g132 ( 
.A(n_115),
.B(n_20),
.CON(n_132),
.SN(n_132)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_24),
.Y(n_116)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_102),
.Y(n_126)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_81),
.B1(n_79),
.B2(n_51),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_119),
.A2(n_90),
.B1(n_92),
.B2(n_96),
.Y(n_159)
);

AOI32xp33_ASAP7_75t_L g120 ( 
.A1(n_115),
.A2(n_70),
.A3(n_86),
.B1(n_82),
.B2(n_78),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_120),
.B(n_104),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_121),
.B(n_130),
.Y(n_152)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_128),
.Y(n_155)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_138),
.Y(n_161)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_34),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_136),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_112),
.B(n_20),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_132),
.A2(n_134),
.B(n_146),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_2),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_135),
.B(n_149),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_113),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_116),
.B(n_23),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_137),
.B(n_139),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_91),
.B(n_82),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_142),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_85),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_144),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_148),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_55),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_145),
.A2(n_93),
.B1(n_112),
.B2(n_101),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_97),
.B(n_2),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_97),
.B(n_3),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_147),
.A2(n_107),
.B(n_110),
.Y(n_163)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_15),
.Y(n_149)
);

AOI221xp5_ASAP7_75t_L g185 ( 
.A1(n_153),
.A2(n_156),
.B1(n_163),
.B2(n_165),
.C(n_147),
.Y(n_185)
);

AOI21xp33_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_96),
.B(n_101),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_171),
.B1(n_134),
.B2(n_142),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_159),
.A2(n_169),
.B1(n_131),
.B2(n_133),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_123),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_160),
.Y(n_183)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_162),
.B(n_167),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_122),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_164),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_129),
.B(n_110),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_110),
.C(n_114),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_111),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_124),
.B(n_108),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_119),
.A2(n_100),
.B1(n_114),
.B2(n_111),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_170),
.B(n_174),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_145),
.A2(n_119),
.B1(n_138),
.B2(n_132),
.Y(n_171)
);

OR2x2_ASAP7_75t_SL g172 ( 
.A(n_146),
.B(n_98),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_172),
.A2(n_131),
.B(n_118),
.Y(n_192)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_177),
.B(n_173),
.Y(n_197)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_176),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_180),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_163),
.B(n_124),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_181),
.Y(n_209)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_175),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_177),
.B(n_146),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_R g182 ( 
.A(n_165),
.B(n_147),
.Y(n_182)
);

AOI221xp5_ASAP7_75t_L g210 ( 
.A1(n_182),
.A2(n_185),
.B1(n_186),
.B2(n_190),
.C(n_192),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_168),
.B(n_119),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_188),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_168),
.B(n_13),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_155),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_191),
.Y(n_211)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_166),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_128),
.Y(n_195)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_195),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_197),
.Y(n_204)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_198),
.A2(n_159),
.B1(n_170),
.B2(n_162),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_200),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_187),
.A2(n_160),
.B(n_151),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_201),
.A2(n_181),
.B(n_188),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_191),
.A2(n_186),
.B1(n_193),
.B2(n_190),
.Y(n_203)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_207),
.C(n_212),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_161),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_196),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_215),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_161),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_183),
.A2(n_153),
.B1(n_151),
.B2(n_154),
.Y(n_214)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_214),
.Y(n_218)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_194),
.Y(n_215)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_172),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_224),
.C(n_225),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_222),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_183),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_227),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_158),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_178),
.C(n_180),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_152),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_184),
.C(n_154),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_229),
.C(n_209),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_184),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_235),
.C(n_236),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_214),
.C(n_199),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_203),
.C(n_211),
.Y(n_236)
);

AOI321xp33_ASAP7_75t_L g237 ( 
.A1(n_221),
.A2(n_213),
.A3(n_200),
.B1(n_150),
.B2(n_206),
.C(n_189),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_238),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_213),
.C(n_118),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_220),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_232),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_174),
.C(n_148),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_240),
.Y(n_242)
);

MAJx2_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_229),
.C(n_218),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_13),
.C(n_12),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_244),
.A2(n_248),
.B(n_4),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_239),
.A2(n_216),
.B1(n_226),
.B2(n_223),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_3),
.Y(n_251)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_233),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_10),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_222),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_143),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_249),
.A2(n_251),
.B(n_252),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_140),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_253),
.Y(n_257)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_254),
.B(n_10),
.CI(n_12),
.CON(n_258),
.SN(n_258)
);

NOR2xp67_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_248),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_5),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_241),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_260),
.C(n_261),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_257),
.A2(n_242),
.B(n_243),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_260),
.B(n_256),
.C(n_6),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_263),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_262),
.Y(n_265)
);


endmodule