module fake_netlist_5_1249_n_1255 (n_137, n_210, n_168, n_260, n_164, n_191, n_286, n_91, n_208, n_82, n_122, n_194, n_282, n_142, n_176, n_10, n_214, n_140, n_24, n_248, n_124, n_86, n_136, n_146, n_268, n_182, n_143, n_83, n_132, n_61, n_237, n_90, n_241, n_127, n_75, n_101, n_180, n_184, n_226, n_235, n_65, n_78, n_74, n_144, n_281, n_207, n_240, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_229, n_108, n_231, n_257, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_236, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_249, n_271, n_284, n_46, n_233, n_21, n_94, n_203, n_245, n_274, n_205, n_113, n_38, n_123, n_139, n_105, n_280, n_246, n_80, n_4, n_179, n_125, n_35, n_269, n_167, n_128, n_73, n_234, n_277, n_17, n_92, n_19, n_267, n_149, n_120, n_285, n_232, n_135, n_30, n_156, n_5, n_33, n_126, n_254, n_14, n_225, n_84, n_23, n_202, n_130, n_266, n_272, n_219, n_157, n_258, n_265, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_244, n_251, n_25, n_53, n_160, n_198, n_223, n_288, n_247, n_188, n_190, n_8, n_201, n_158, n_263, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_264, n_283, n_109, n_112, n_212, n_85, n_159, n_163, n_276, n_95, n_119, n_183, n_185, n_243, n_239, n_275, n_175, n_252, n_169, n_59, n_262, n_26, n_255, n_133, n_238, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_290, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_242, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_259, n_273, n_287, n_270, n_222, n_230, n_81, n_118, n_28, n_89, n_279, n_70, n_115, n_68, n_93, n_253, n_261, n_72, n_174, n_186, n_199, n_289, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_256, n_48, n_204, n_50, n_250, n_52, n_278, n_88, n_110, n_216, n_1255);

input n_137;
input n_210;
input n_168;
input n_260;
input n_164;
input n_191;
input n_286;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_282;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_268;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_237;
input n_90;
input n_241;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_235;
input n_65;
input n_78;
input n_74;
input n_144;
input n_281;
input n_207;
input n_240;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_229;
input n_108;
input n_231;
input n_257;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_236;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_249;
input n_271;
input n_284;
input n_46;
input n_233;
input n_21;
input n_94;
input n_203;
input n_245;
input n_274;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_280;
input n_246;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_269;
input n_167;
input n_128;
input n_73;
input n_234;
input n_277;
input n_17;
input n_92;
input n_19;
input n_267;
input n_149;
input n_120;
input n_285;
input n_232;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_254;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_266;
input n_272;
input n_219;
input n_157;
input n_258;
input n_265;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_244;
input n_251;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_288;
input n_247;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_264;
input n_283;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_276;
input n_95;
input n_119;
input n_183;
input n_185;
input n_243;
input n_239;
input n_275;
input n_175;
input n_252;
input n_169;
input n_59;
input n_262;
input n_26;
input n_255;
input n_133;
input n_238;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_290;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_242;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_259;
input n_273;
input n_287;
input n_270;
input n_222;
input n_230;
input n_81;
input n_118;
input n_28;
input n_89;
input n_279;
input n_70;
input n_115;
input n_68;
input n_93;
input n_253;
input n_261;
input n_72;
input n_174;
input n_186;
input n_199;
input n_289;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_256;
input n_48;
input n_204;
input n_50;
input n_250;
input n_52;
input n_278;
input n_88;
input n_110;
input n_216;

output n_1255;

wire n_924;
wire n_977;
wire n_611;
wire n_1126;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1198;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_688;
wire n_800;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_447;
wire n_292;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_373;
wire n_307;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_659;
wire n_1182;
wire n_579;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_291;
wire n_731;
wire n_371;
wire n_709;
wire n_317;
wire n_1236;
wire n_569;
wire n_920;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_308;
wire n_297;
wire n_1078;
wire n_775;
wire n_600;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_350;
wire n_646;
wire n_436;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_496;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1069;
wire n_1075;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_989;
wire n_1039;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1002;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_561;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_596;
wire n_558;
wire n_702;
wire n_822;
wire n_728;
wire n_1162;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_409;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_759;
wire n_806;
wire n_324;
wire n_1189;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_367;
wire n_452;
wire n_525;
wire n_649;
wire n_547;
wire n_1191;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1233;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_1121;
wire n_433;
wire n_314;
wire n_368;
wire n_604;
wire n_949;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_999;
wire n_758;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1054;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_396;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_473;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_337;
wire n_1177;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1006;
wire n_329;
wire n_582;
wire n_309;
wire n_512;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_987;
wire n_767;
wire n_993;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_513;
wire n_1094;
wire n_560;
wire n_340;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_996;
wire n_921;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1037;
wire n_1080;
wire n_426;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_960;
wire n_1123;
wire n_1047;
wire n_634;
wire n_1252;
wire n_348;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_950;
wire n_380;
wire n_419;
wire n_444;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_376;
wire n_967;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_690;
wire n_583;
wire n_302;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_385;
wire n_507;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_341;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1214;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1096;
wire n_833;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_669;
wire n_472;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_311;
wire n_830;
wire n_801;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1019;
wire n_1105;
wire n_304;
wire n_577;
wire n_338;
wire n_693;
wire n_990;
wire n_836;
wire n_975;
wire n_567;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1164;
wire n_489;
wire n_1174;
wire n_617;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1059;
wire n_1133;
wire n_557;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_393;
wire n_487;
wire n_665;
wire n_421;
wire n_910;
wire n_768;
wire n_1136;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_427;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_536;
wire n_872;
wire n_594;
wire n_1155;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_605;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_501;
wire n_823;
wire n_725;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_788;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_737;
wire n_986;
wire n_509;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_862;
wire n_760;
wire n_381;
wire n_390;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_570;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_400;
wire n_930;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_432;
wire n_839;
wire n_1210;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1012;
wire n_903;
wire n_740;
wire n_384;
wire n_1061;
wire n_333;
wire n_462;
wire n_1193;
wire n_1113;
wire n_1226;
wire n_722;
wire n_844;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_312;
wire n_1076;
wire n_1091;
wire n_494;
wire n_641;
wire n_730;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_712;
wire n_1042;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_491;
wire n_1074;
wire n_566;
wire n_565;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_334;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_533;
wire n_1251;

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_116),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_266),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_105),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_274),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_106),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_35),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_123),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_27),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_124),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_80),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_110),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_128),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_264),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_28),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_247),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_187),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_53),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_20),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_83),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_219),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_1),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g312 ( 
.A(n_120),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_125),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_269),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_138),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_209),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_223),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_202),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_160),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_200),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_270),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_25),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_212),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_210),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_181),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_268),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_230),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_87),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_50),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_287),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_151),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_234),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_115),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_281),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_66),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_108),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_77),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_55),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_76),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_99),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_17),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_191),
.Y(n_342)
);

BUFx5_ASAP7_75t_L g343 ( 
.A(n_240),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_218),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_233),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_65),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_130),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_157),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_61),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_198),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_82),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_72),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_2),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_11),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_71),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_88),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_0),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_45),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_109),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_242),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_0),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_131),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_174),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_44),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_119),
.Y(n_365)
);

INVx2_ASAP7_75t_SL g366 ( 
.A(n_189),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_13),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_265),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_232),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_194),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_251),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_197),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_173),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_52),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_248),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_192),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_178),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_195),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_253),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_63),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_214),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_142),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_97),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_38),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_23),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_26),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_94),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_102),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_118),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_127),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_284),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_9),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_107),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_271),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_205),
.Y(n_395)
);

INVx2_ASAP7_75t_SL g396 ( 
.A(n_179),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_256),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_12),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_213),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_112),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_126),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_183),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_227),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_152),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_1),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_7),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_85),
.Y(n_407)
);

BUFx8_ASAP7_75t_SL g408 ( 
.A(n_225),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_150),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_148),
.Y(n_410)
);

BUFx10_ASAP7_75t_L g411 ( 
.A(n_149),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_211),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_263),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_290),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_29),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_67),
.Y(n_416)
);

CKINVDCx14_ASAP7_75t_R g417 ( 
.A(n_259),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_286),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_278),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_79),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_136),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_175),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_272),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_6),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_221),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_2),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_5),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_216),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_236),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_147),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_57),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_182),
.Y(n_432)
);

BUFx10_ASAP7_75t_L g433 ( 
.A(n_69),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_143),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_237),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_100),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_96),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_103),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_24),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_60),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_31),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_172),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_86),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_261),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_154),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_167),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_4),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_204),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_224),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_246),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_84),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_207),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_22),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_57),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_235),
.Y(n_455)
);

BUFx10_ASAP7_75t_L g456 ( 
.A(n_48),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_169),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_32),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_92),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_44),
.Y(n_460)
);

BUFx10_ASAP7_75t_L g461 ( 
.A(n_11),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_36),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_35),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_171),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_45),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_21),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_282),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_111),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_220),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_129),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_250),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_104),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_168),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_260),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_408),
.Y(n_475)
);

NOR2x1_ASAP7_75t_L g476 ( 
.A(n_299),
.B(n_3),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_351),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_322),
.B(n_3),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_322),
.B(n_4),
.Y(n_479)
);

BUFx8_ASAP7_75t_SL g480 ( 
.A(n_466),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_292),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_299),
.B(n_5),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_341),
.Y(n_483)
);

BUFx12f_ASAP7_75t_L g484 ( 
.A(n_456),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_351),
.Y(n_485)
);

AND2x6_ASAP7_75t_L g486 ( 
.A(n_351),
.B(n_58),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_341),
.B(n_441),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_300),
.B(n_6),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_411),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_341),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_320),
.B(n_7),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_301),
.B(n_8),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_398),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_341),
.B(n_8),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_351),
.Y(n_495)
);

CKINVDCx6p67_ASAP7_75t_R g496 ( 
.A(n_424),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_309),
.B(n_9),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_441),
.Y(n_498)
);

AND2x6_ASAP7_75t_L g499 ( 
.A(n_471),
.B(n_59),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_301),
.B(n_10),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_320),
.B(n_10),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_337),
.B(n_12),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_441),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_337),
.B(n_13),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_363),
.B(n_380),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_471),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_441),
.B(n_14),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_363),
.B(n_14),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_471),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_453),
.Y(n_510)
);

INVx6_ASAP7_75t_L g511 ( 
.A(n_411),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_471),
.Y(n_512)
);

INVx5_ASAP7_75t_L g513 ( 
.A(n_453),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_453),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_433),
.Y(n_515)
);

AND2x6_ASAP7_75t_L g516 ( 
.A(n_380),
.B(n_62),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_403),
.B(n_15),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_453),
.B(n_15),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_403),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_414),
.B(n_16),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_414),
.B(n_16),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_398),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_296),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_425),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_343),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_298),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_317),
.B(n_17),
.Y(n_527)
);

BUFx12f_ASAP7_75t_L g528 ( 
.A(n_456),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_425),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_343),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_432),
.Y(n_531)
);

NOR2x1_ASAP7_75t_L g532 ( 
.A(n_326),
.B(n_18),
.Y(n_532)
);

INVx5_ASAP7_75t_L g533 ( 
.A(n_433),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_343),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_432),
.B(n_18),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_307),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_434),
.B(n_19),
.Y(n_537)
);

CKINVDCx6p67_ASAP7_75t_R g538 ( 
.A(n_461),
.Y(n_538)
);

INVx5_ASAP7_75t_L g539 ( 
.A(n_461),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_343),
.Y(n_540)
);

INVx5_ASAP7_75t_L g541 ( 
.A(n_312),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_343),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_293),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_343),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_308),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_358),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_458),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_417),
.B(n_19),
.Y(n_548)
);

INVx5_ASAP7_75t_L g549 ( 
.A(n_324),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_468),
.B(n_20),
.Y(n_550)
);

INVx5_ASAP7_75t_L g551 ( 
.A(n_349),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_434),
.Y(n_552)
);

CKINVDCx11_ASAP7_75t_R g553 ( 
.A(n_291),
.Y(n_553)
);

INVx5_ASAP7_75t_L g554 ( 
.A(n_362),
.Y(n_554)
);

BUFx8_ASAP7_75t_SL g555 ( 
.A(n_314),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_364),
.Y(n_556)
);

INVx6_ASAP7_75t_L g557 ( 
.A(n_311),
.Y(n_557)
);

INVx5_ASAP7_75t_L g558 ( 
.A(n_366),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_396),
.B(n_21),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_387),
.B(n_323),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_406),
.B(n_22),
.Y(n_561)
);

INVx5_ASAP7_75t_L g562 ( 
.A(n_458),
.Y(n_562)
);

CKINVDCx11_ASAP7_75t_R g563 ( 
.A(n_330),
.Y(n_563)
);

INVx5_ASAP7_75t_L g564 ( 
.A(n_329),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_294),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_335),
.B(n_23),
.Y(n_566)
);

INVx5_ASAP7_75t_L g567 ( 
.A(n_338),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_353),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_374),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_295),
.Y(n_570)
);

INVx4_ASAP7_75t_L g571 ( 
.A(n_297),
.Y(n_571)
);

BUFx8_ASAP7_75t_SL g572 ( 
.A(n_356),
.Y(n_572)
);

BUFx12f_ASAP7_75t_L g573 ( 
.A(n_354),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_431),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_523),
.B(n_328),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_548),
.A2(n_391),
.B1(n_377),
.B2(n_357),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_560),
.A2(n_361),
.B1(n_384),
.B2(n_367),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_498),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_526),
.B(n_420),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_568),
.B(n_303),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_545),
.B(n_306),
.Y(n_581)
);

OR2x6_ASAP7_75t_L g582 ( 
.A(n_573),
.B(n_439),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_527),
.A2(n_304),
.B1(n_386),
.B2(n_385),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_483),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_533),
.B(n_310),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_481),
.B(n_302),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_560),
.A2(n_405),
.B1(n_415),
.B2(n_392),
.Y(n_587)
);

INVx8_ASAP7_75t_L g588 ( 
.A(n_555),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_493),
.B(n_426),
.Y(n_589)
);

OAI22xp33_ASAP7_75t_SL g590 ( 
.A1(n_550),
.A2(n_454),
.B1(n_462),
.B2(n_427),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_490),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_527),
.A2(n_465),
.B1(n_463),
.B2(n_316),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_539),
.B(n_315),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_533),
.B(n_319),
.Y(n_594)
);

OAI22xp33_ASAP7_75t_L g595 ( 
.A1(n_550),
.A2(n_460),
.B1(n_447),
.B2(n_313),
.Y(n_595)
);

AO22x2_ASAP7_75t_L g596 ( 
.A1(n_482),
.A2(n_318),
.B1(n_333),
.B2(n_305),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_478),
.A2(n_325),
.B1(n_327),
.B2(n_321),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_539),
.B(n_331),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_498),
.Y(n_599)
);

OAI22xp33_ASAP7_75t_SL g600 ( 
.A1(n_566),
.A2(n_348),
.B1(n_350),
.B2(n_345),
.Y(n_600)
);

AO22x2_ASAP7_75t_L g601 ( 
.A1(n_482),
.A2(n_359),
.B1(n_365),
.B2(n_355),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_510),
.Y(n_602)
);

OAI22xp33_ASAP7_75t_L g603 ( 
.A1(n_566),
.A2(n_373),
.B1(n_376),
.B2(n_371),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_541),
.B(n_378),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_572),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_511),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_489),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_541),
.B(n_382),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_479),
.A2(n_334),
.B1(n_336),
.B2(n_332),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_488),
.A2(n_340),
.B1(n_342),
.B2(n_339),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_497),
.A2(n_496),
.B1(n_559),
.B2(n_501),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_510),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_539),
.B(n_344),
.Y(n_613)
);

AOI22x1_ASAP7_75t_L g614 ( 
.A1(n_535),
.A2(n_394),
.B1(n_399),
.B2(n_388),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_561),
.A2(n_347),
.B1(n_352),
.B2(n_346),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_503),
.Y(n_616)
);

NOR2x1p5_ASAP7_75t_L g617 ( 
.A(n_515),
.B(n_360),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_533),
.B(n_368),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_559),
.A2(n_370),
.B1(n_372),
.B2(n_369),
.Y(n_619)
);

OR2x6_ASAP7_75t_L g620 ( 
.A(n_484),
.B(n_401),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_511),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_514),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_514),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_570),
.B(n_404),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_522),
.B(n_24),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_532),
.A2(n_379),
.B1(n_381),
.B2(n_375),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_477),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_543),
.B(n_383),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_532),
.A2(n_390),
.B1(n_393),
.B2(n_389),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_477),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_477),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_543),
.B(n_395),
.Y(n_632)
);

OAI22xp33_ASAP7_75t_L g633 ( 
.A1(n_491),
.A2(n_422),
.B1(n_436),
.B2(n_416),
.Y(n_633)
);

OR2x6_ASAP7_75t_L g634 ( 
.A(n_528),
.B(n_437),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_485),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_519),
.Y(n_636)
);

OAI22xp33_ASAP7_75t_L g637 ( 
.A1(n_491),
.A2(n_446),
.B1(n_448),
.B2(n_444),
.Y(n_637)
);

OAI22xp33_ASAP7_75t_SL g638 ( 
.A1(n_501),
.A2(n_469),
.B1(n_472),
.B2(n_457),
.Y(n_638)
);

OAI22xp33_ASAP7_75t_SL g639 ( 
.A1(n_502),
.A2(n_473),
.B1(n_400),
.B2(n_402),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_565),
.B(n_397),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_557),
.A2(n_475),
.B1(n_538),
.B2(n_500),
.Y(n_641)
);

OAI22xp33_ASAP7_75t_SL g642 ( 
.A1(n_502),
.A2(n_409),
.B1(n_410),
.B2(n_407),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_557),
.A2(n_413),
.B1(n_418),
.B2(n_412),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_565),
.B(n_419),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_541),
.B(n_421),
.Y(n_645)
);

OAI22xp33_ASAP7_75t_SL g646 ( 
.A1(n_504),
.A2(n_474),
.B1(n_470),
.B2(n_467),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_SL g647 ( 
.A1(n_535),
.A2(n_464),
.B1(n_459),
.B2(n_455),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_485),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_571),
.B(n_423),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_571),
.B(n_428),
.Y(n_650)
);

AO22x2_ASAP7_75t_L g651 ( 
.A1(n_492),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_651)
);

CKINVDCx6p67_ASAP7_75t_R g652 ( 
.A(n_553),
.Y(n_652)
);

OA22x2_ASAP7_75t_L g653 ( 
.A1(n_536),
.A2(n_452),
.B1(n_451),
.B2(n_450),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_485),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_495),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_564),
.B(n_429),
.Y(n_656)
);

OAI22xp33_ASAP7_75t_L g657 ( 
.A1(n_504),
.A2(n_449),
.B1(n_445),
.B2(n_443),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_564),
.B(n_430),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_575),
.B(n_564),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_627),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_631),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_624),
.B(n_492),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_631),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_630),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_648),
.Y(n_665)
);

INVx4_ASAP7_75t_SL g666 ( 
.A(n_624),
.Y(n_666)
);

INVxp33_ASAP7_75t_L g667 ( 
.A(n_579),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_648),
.Y(n_668)
);

XNOR2x2_ASAP7_75t_L g669 ( 
.A(n_651),
.B(n_476),
.Y(n_669)
);

XOR2x2_ASAP7_75t_L g670 ( 
.A(n_583),
.B(n_476),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_655),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_655),
.Y(n_672)
);

BUFx5_ASAP7_75t_L g673 ( 
.A(n_591),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_636),
.B(n_525),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_635),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_584),
.B(n_530),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_654),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_622),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_623),
.Y(n_679)
);

NAND2xp33_ASAP7_75t_R g680 ( 
.A(n_607),
.B(n_500),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_599),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_599),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_578),
.Y(n_683)
);

INVx1_ASAP7_75t_SL g684 ( 
.A(n_589),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_578),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_616),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_586),
.B(n_549),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_602),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_602),
.Y(n_689)
);

INVxp67_ASAP7_75t_SL g690 ( 
.A(n_612),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_SL g691 ( 
.A(n_595),
.B(n_486),
.Y(n_691)
);

XOR2xp5_ASAP7_75t_L g692 ( 
.A(n_605),
.B(n_576),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_612),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_625),
.Y(n_694)
);

NOR2xp67_ASAP7_75t_L g695 ( 
.A(n_643),
.B(n_567),
.Y(n_695)
);

OAI21xp5_ASAP7_75t_L g696 ( 
.A1(n_653),
.A2(n_517),
.B(n_508),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_580),
.B(n_567),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_604),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_581),
.B(n_567),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_588),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_608),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_577),
.B(n_547),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_614),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_614),
.Y(n_704)
);

CKINVDCx20_ASAP7_75t_R g705 ( 
.A(n_652),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_596),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_596),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_601),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_601),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_656),
.Y(n_710)
);

INVx4_ASAP7_75t_L g711 ( 
.A(n_658),
.Y(n_711)
);

AND2x6_ASAP7_75t_L g712 ( 
.A(n_626),
.B(n_494),
.Y(n_712)
);

INVxp67_ASAP7_75t_SL g713 ( 
.A(n_633),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_585),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_594),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_618),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_638),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_600),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_645),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_629),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_617),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_606),
.B(n_547),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_651),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_628),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_632),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_649),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_650),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_621),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_592),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_619),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_587),
.B(n_562),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_597),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_609),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_590),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_637),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_603),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_657),
.B(n_549),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_615),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_640),
.B(n_549),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_644),
.B(n_551),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_647),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_610),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_639),
.B(n_534),
.Y(n_743)
);

AND2x2_ASAP7_75t_SL g744 ( 
.A(n_641),
.B(n_508),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_611),
.Y(n_745)
);

OR2x2_ASAP7_75t_SL g746 ( 
.A(n_646),
.B(n_517),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_588),
.Y(n_747)
);

CKINVDCx16_ASAP7_75t_R g748 ( 
.A(n_582),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_719),
.B(n_642),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_667),
.B(n_546),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_700),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_714),
.B(n_519),
.Y(n_752)
);

AND2x4_ASAP7_75t_L g753 ( 
.A(n_666),
.B(n_569),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_667),
.B(n_556),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_711),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_728),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_683),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_690),
.B(n_519),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_710),
.Y(n_759)
);

HB1xp67_ASAP7_75t_L g760 ( 
.A(n_722),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_660),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_662),
.B(n_696),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_666),
.B(n_574),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_685),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_662),
.B(n_505),
.Y(n_765)
);

NAND2x1p5_ASAP7_75t_L g766 ( 
.A(n_711),
.B(n_540),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_704),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_730),
.B(n_524),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_688),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_687),
.B(n_524),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_689),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_666),
.B(n_582),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_715),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_693),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_696),
.B(n_505),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_716),
.Y(n_776)
);

OAI21xp5_ASAP7_75t_L g777 ( 
.A1(n_703),
.A2(n_521),
.B(n_520),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_659),
.B(n_494),
.Y(n_778)
);

AND2x2_ASAP7_75t_SL g779 ( 
.A(n_691),
.B(n_744),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_676),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_745),
.B(n_507),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_681),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_682),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_727),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_713),
.B(n_507),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_676),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_674),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_713),
.B(n_518),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_702),
.B(n_620),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_674),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_687),
.B(n_529),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_720),
.B(n_435),
.Y(n_792)
);

AND2x4_ASAP7_75t_L g793 ( 
.A(n_707),
.B(n_516),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_698),
.B(n_529),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_743),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_724),
.B(n_518),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_725),
.B(n_520),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_686),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_661),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_743),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_726),
.B(n_521),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_721),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_701),
.B(n_529),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_664),
.Y(n_804)
);

INVx4_ASAP7_75t_L g805 ( 
.A(n_673),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_675),
.Y(n_806)
);

BUFx3_ASAP7_75t_L g807 ( 
.A(n_747),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_678),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_679),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_736),
.B(n_684),
.Y(n_810)
);

INVx4_ASAP7_75t_L g811 ( 
.A(n_673),
.Y(n_811)
);

INVx3_ASAP7_75t_L g812 ( 
.A(n_677),
.Y(n_812)
);

INVxp67_ASAP7_75t_L g813 ( 
.A(n_684),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_735),
.B(n_537),
.Y(n_814)
);

OR2x2_ASAP7_75t_SL g815 ( 
.A(n_741),
.B(n_537),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_663),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_665),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_668),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_742),
.B(n_553),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_671),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_672),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_680),
.Y(n_822)
);

OAI21xp5_ASAP7_75t_L g823 ( 
.A1(n_729),
.A2(n_516),
.B(n_487),
.Y(n_823)
);

BUFx2_ASAP7_75t_L g824 ( 
.A(n_712),
.Y(n_824)
);

INVx3_ASAP7_75t_L g825 ( 
.A(n_673),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_694),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_717),
.B(n_718),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_742),
.B(n_563),
.Y(n_828)
);

AND2x4_ASAP7_75t_L g829 ( 
.A(n_706),
.B(n_516),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_708),
.Y(n_830)
);

INVx1_ASAP7_75t_SL g831 ( 
.A(n_731),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_709),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_697),
.B(n_699),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_673),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_739),
.B(n_531),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_673),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_739),
.B(n_531),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_734),
.B(n_542),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_SL g839 ( 
.A(n_748),
.B(n_480),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_740),
.B(n_531),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_673),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_810),
.B(n_744),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_757),
.Y(n_843)
);

AND2x6_ASAP7_75t_L g844 ( 
.A(n_795),
.B(n_723),
.Y(n_844)
);

NAND2x1_ASAP7_75t_L g845 ( 
.A(n_805),
.B(n_486),
.Y(n_845)
);

INVx6_ASAP7_75t_SL g846 ( 
.A(n_772),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_757),
.Y(n_847)
);

INVx4_ASAP7_75t_L g848 ( 
.A(n_755),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_787),
.B(n_712),
.Y(n_849)
);

OR2x2_ASAP7_75t_L g850 ( 
.A(n_813),
.B(n_746),
.Y(n_850)
);

NAND2x1p5_ASAP7_75t_L g851 ( 
.A(n_755),
.B(n_695),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_765),
.B(n_712),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_759),
.B(n_732),
.Y(n_853)
);

BUFx3_ASAP7_75t_L g854 ( 
.A(n_807),
.Y(n_854)
);

OR2x6_ASAP7_75t_L g855 ( 
.A(n_772),
.B(n_620),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_759),
.B(n_733),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_773),
.B(n_738),
.Y(n_857)
);

NAND2x1p5_ASAP7_75t_L g858 ( 
.A(n_755),
.B(n_593),
.Y(n_858)
);

INVx4_ASAP7_75t_L g859 ( 
.A(n_755),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_765),
.B(n_712),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_790),
.B(n_712),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_769),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_769),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_822),
.B(n_563),
.Y(n_864)
);

AND2x6_ASAP7_75t_L g865 ( 
.A(n_795),
.B(n_737),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_810),
.B(n_670),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_755),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_764),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_771),
.Y(n_869)
);

NOR2xp67_ASAP7_75t_L g870 ( 
.A(n_751),
.B(n_737),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_773),
.B(n_634),
.Y(n_871)
);

NOR2x1_ASAP7_75t_SL g872 ( 
.A(n_805),
.B(n_634),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_790),
.B(n_740),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_760),
.B(n_692),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_780),
.B(n_691),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_815),
.B(n_669),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_750),
.Y(n_877)
);

AND2x4_ASAP7_75t_L g878 ( 
.A(n_776),
.B(n_598),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_812),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_799),
.Y(n_880)
);

OR2x2_ASAP7_75t_L g881 ( 
.A(n_815),
.B(n_613),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_780),
.B(n_552),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_750),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_776),
.B(n_705),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_762),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_774),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_786),
.B(n_552),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_754),
.Y(n_888)
);

INVxp67_ASAP7_75t_L g889 ( 
.A(n_754),
.Y(n_889)
);

NOR2xp67_ASAP7_75t_L g890 ( 
.A(n_822),
.B(n_438),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_784),
.B(n_64),
.Y(n_891)
);

AND2x4_ASAP7_75t_L g892 ( 
.A(n_784),
.B(n_68),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_797),
.B(n_680),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_785),
.B(n_440),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_786),
.B(n_552),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_795),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_816),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_775),
.B(n_551),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_775),
.B(n_551),
.Y(n_899)
);

OR2x2_ASAP7_75t_L g900 ( 
.A(n_785),
.B(n_442),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_795),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_797),
.B(n_562),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_816),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_756),
.B(n_70),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_817),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_818),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_778),
.B(n_554),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_846),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_885),
.B(n_788),
.Y(n_909)
);

INVx6_ASAP7_75t_SL g910 ( 
.A(n_855),
.Y(n_910)
);

INVx8_ASAP7_75t_L g911 ( 
.A(n_844),
.Y(n_911)
);

BUFx12f_ASAP7_75t_L g912 ( 
.A(n_855),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_893),
.B(n_819),
.Y(n_913)
);

INVx6_ASAP7_75t_SL g914 ( 
.A(n_871),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_889),
.B(n_828),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_868),
.Y(n_916)
);

INVx5_ASAP7_75t_L g917 ( 
.A(n_867),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_869),
.Y(n_918)
);

BUFx2_ASAP7_75t_L g919 ( 
.A(n_846),
.Y(n_919)
);

BUFx2_ASAP7_75t_SL g920 ( 
.A(n_854),
.Y(n_920)
);

AOI22xp33_ASAP7_75t_L g921 ( 
.A1(n_852),
.A2(n_779),
.B1(n_800),
.B2(n_795),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_862),
.Y(n_922)
);

BUFx12f_ASAP7_75t_L g923 ( 
.A(n_871),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_867),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_853),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_886),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_905),
.Y(n_927)
);

BUFx12f_ASAP7_75t_L g928 ( 
.A(n_884),
.Y(n_928)
);

BUFx2_ASAP7_75t_L g929 ( 
.A(n_884),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_874),
.Y(n_930)
);

BUFx2_ASAP7_75t_L g931 ( 
.A(n_853),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_906),
.Y(n_932)
);

INVx4_ASAP7_75t_L g933 ( 
.A(n_867),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_843),
.Y(n_934)
);

NAND2x1p5_ASAP7_75t_L g935 ( 
.A(n_848),
.B(n_824),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_856),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_856),
.B(n_779),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_875),
.B(n_788),
.Y(n_938)
);

INVx1_ASAP7_75t_SL g939 ( 
.A(n_842),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_860),
.A2(n_824),
.B1(n_762),
.B2(n_800),
.Y(n_940)
);

OR2x2_ASAP7_75t_L g941 ( 
.A(n_894),
.B(n_778),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_847),
.Y(n_942)
);

BUFx3_ASAP7_75t_L g943 ( 
.A(n_857),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_877),
.B(n_792),
.Y(n_944)
);

INVx1_ASAP7_75t_SL g945 ( 
.A(n_850),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_863),
.Y(n_946)
);

BUFx12f_ASAP7_75t_L g947 ( 
.A(n_857),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_861),
.B(n_800),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_864),
.Y(n_949)
);

NAND2x1p5_ASAP7_75t_L g950 ( 
.A(n_848),
.B(n_800),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_866),
.Y(n_951)
);

INVx3_ASAP7_75t_SL g952 ( 
.A(n_876),
.Y(n_952)
);

NAND2x1p5_ASAP7_75t_L g953 ( 
.A(n_859),
.B(n_772),
.Y(n_953)
);

NAND2x1p5_ASAP7_75t_L g954 ( 
.A(n_859),
.B(n_802),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_897),
.Y(n_955)
);

BUFx12f_ASAP7_75t_L g956 ( 
.A(n_904),
.Y(n_956)
);

INVx4_ASAP7_75t_L g957 ( 
.A(n_896),
.Y(n_957)
);

INVx6_ASAP7_75t_L g958 ( 
.A(n_904),
.Y(n_958)
);

INVx1_ASAP7_75t_SL g959 ( 
.A(n_849),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_881),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_873),
.B(n_800),
.Y(n_961)
);

BUFx4f_ASAP7_75t_SL g962 ( 
.A(n_878),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_896),
.Y(n_963)
);

INVx1_ASAP7_75t_SL g964 ( 
.A(n_945),
.Y(n_964)
);

AOI22xp33_ASAP7_75t_L g965 ( 
.A1(n_913),
.A2(n_938),
.B1(n_939),
.B2(n_814),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_916),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_938),
.B(n_883),
.Y(n_967)
);

BUFx12f_ASAP7_75t_L g968 ( 
.A(n_923),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_909),
.B(n_888),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_909),
.B(n_801),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_SL g971 ( 
.A1(n_960),
.A2(n_865),
.B1(n_839),
.B2(n_814),
.Y(n_971)
);

AOI22xp33_ASAP7_75t_L g972 ( 
.A1(n_939),
.A2(n_781),
.B1(n_777),
.B2(n_865),
.Y(n_972)
);

BUFx4f_ASAP7_75t_L g973 ( 
.A(n_956),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_SL g974 ( 
.A1(n_945),
.A2(n_789),
.B(n_831),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_918),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_926),
.Y(n_976)
);

BUFx2_ASAP7_75t_L g977 ( 
.A(n_914),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_921),
.A2(n_896),
.B1(n_901),
.B2(n_870),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_947),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_912),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_941),
.A2(n_781),
.B1(n_865),
.B2(n_796),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_928),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_L g983 ( 
.A1(n_937),
.A2(n_865),
.B1(n_796),
.B2(n_792),
.Y(n_983)
);

INVx6_ASAP7_75t_L g984 ( 
.A(n_917),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_927),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_951),
.A2(n_890),
.B1(n_878),
.B2(n_833),
.Y(n_986)
);

BUFx8_ASAP7_75t_SL g987 ( 
.A(n_929),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_932),
.Y(n_988)
);

BUFx4f_ASAP7_75t_SL g989 ( 
.A(n_914),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_931),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_934),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_942),
.Y(n_992)
);

AO22x1_ASAP7_75t_L g993 ( 
.A1(n_949),
.A2(n_844),
.B1(n_892),
.B2(n_891),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_946),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_955),
.Y(n_995)
);

CKINVDCx11_ASAP7_75t_R g996 ( 
.A(n_952),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_L g997 ( 
.A1(n_944),
.A2(n_801),
.B1(n_827),
.B2(n_903),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_961),
.B(n_902),
.Y(n_998)
);

INVx6_ASAP7_75t_L g999 ( 
.A(n_917),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_922),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_961),
.Y(n_1001)
);

INVx6_ASAP7_75t_L g1002 ( 
.A(n_917),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_908),
.Y(n_1003)
);

INVxp67_ASAP7_75t_L g1004 ( 
.A(n_920),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_959),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_959),
.Y(n_1006)
);

OAI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_962),
.A2(n_900),
.B1(n_826),
.B2(n_749),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_919),
.Y(n_1008)
);

CKINVDCx20_ASAP7_75t_R g1009 ( 
.A(n_930),
.Y(n_1009)
);

INVx6_ASAP7_75t_L g1010 ( 
.A(n_963),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_915),
.A2(n_827),
.B1(n_838),
.B2(n_880),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_958),
.Y(n_1012)
);

CKINVDCx11_ASAP7_75t_R g1013 ( 
.A(n_943),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_958),
.Y(n_1014)
);

INVx6_ASAP7_75t_L g1015 ( 
.A(n_963),
.Y(n_1015)
);

OAI21xp5_ASAP7_75t_SL g1016 ( 
.A1(n_971),
.A2(n_789),
.B(n_833),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_975),
.Y(n_1017)
);

INVx2_ASAP7_75t_SL g1018 ( 
.A(n_973),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_976),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_971),
.A2(n_1007),
.B1(n_981),
.B2(n_983),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_969),
.B(n_925),
.Y(n_1021)
);

AOI222xp33_ASAP7_75t_L g1022 ( 
.A1(n_970),
.A2(n_936),
.B1(n_838),
.B2(n_832),
.C1(n_823),
.C2(n_802),
.Y(n_1022)
);

INVx4_ASAP7_75t_L g1023 ( 
.A(n_984),
.Y(n_1023)
);

OAI222xp33_ASAP7_75t_L g1024 ( 
.A1(n_965),
.A2(n_940),
.B1(n_948),
.B2(n_768),
.C1(n_899),
.C2(n_898),
.Y(n_1024)
);

AOI222xp33_ASAP7_75t_L g1025 ( 
.A1(n_1007),
.A2(n_872),
.B1(n_798),
.B2(n_820),
.C1(n_516),
.C2(n_782),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_985),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_966),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_991),
.Y(n_1028)
);

CKINVDCx6p67_ASAP7_75t_R g1029 ( 
.A(n_968),
.Y(n_1029)
);

AOI22xp33_ASAP7_75t_L g1030 ( 
.A1(n_981),
.A2(n_844),
.B1(n_821),
.B2(n_891),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_988),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_992),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_1000),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_965),
.A2(n_940),
.B1(n_851),
.B2(n_901),
.Y(n_1034)
);

NAND2x1p5_ASAP7_75t_L g1035 ( 
.A(n_1005),
.B(n_901),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_1006),
.B(n_830),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_994),
.Y(n_1037)
);

OAI222xp33_ASAP7_75t_L g1038 ( 
.A1(n_964),
.A2(n_948),
.B1(n_954),
.B2(n_950),
.C1(n_935),
.C2(n_907),
.Y(n_1038)
);

OAI222xp33_ASAP7_75t_L g1039 ( 
.A1(n_986),
.A2(n_935),
.B1(n_953),
.B2(n_858),
.C1(n_752),
.C2(n_770),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_995),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_SL g1041 ( 
.A1(n_974),
.A2(n_783),
.B(n_829),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_997),
.A2(n_911),
.B1(n_879),
.B2(n_766),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_998),
.A2(n_808),
.B1(n_809),
.B2(n_763),
.Y(n_1043)
);

AOI22xp33_ASAP7_75t_SL g1044 ( 
.A1(n_1009),
.A2(n_911),
.B1(n_756),
.B2(n_879),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_967),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1001),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1011),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1011),
.Y(n_1048)
);

OR2x2_ASAP7_75t_L g1049 ( 
.A(n_990),
.B(n_791),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_984),
.Y(n_1050)
);

OR2x2_ASAP7_75t_SL g1051 ( 
.A(n_1012),
.B(n_910),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_972),
.A2(n_911),
.B1(n_766),
.B2(n_910),
.Y(n_1052)
);

INVx2_ASAP7_75t_SL g1053 ( 
.A(n_973),
.Y(n_1053)
);

INVxp67_ASAP7_75t_L g1054 ( 
.A(n_987),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_996),
.A2(n_982),
.B1(n_1013),
.B2(n_980),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_1013),
.A2(n_753),
.B1(n_812),
.B2(n_803),
.Y(n_1056)
);

INVx5_ASAP7_75t_L g1057 ( 
.A(n_984),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_1004),
.B(n_1008),
.Y(n_1058)
);

INVx3_ASAP7_75t_L g1059 ( 
.A(n_999),
.Y(n_1059)
);

OAI21xp33_ASAP7_75t_L g1060 ( 
.A1(n_1003),
.A2(n_794),
.B(n_758),
.Y(n_1060)
);

AOI22xp33_ASAP7_75t_L g1061 ( 
.A1(n_979),
.A2(n_812),
.B1(n_806),
.B2(n_761),
.Y(n_1061)
);

INVx1_ASAP7_75t_SL g1062 ( 
.A(n_1010),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_1014),
.B(n_804),
.Y(n_1063)
);

CKINVDCx20_ASAP7_75t_R g1064 ( 
.A(n_989),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_978),
.A2(n_806),
.B1(n_761),
.B2(n_804),
.Y(n_1065)
);

AOI221xp5_ASAP7_75t_L g1066 ( 
.A1(n_1020),
.A2(n_487),
.B1(n_993),
.B2(n_835),
.C(n_837),
.Y(n_1066)
);

NAND3xp33_ASAP7_75t_L g1067 ( 
.A(n_1041),
.B(n_840),
.C(n_806),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_1044),
.A2(n_999),
.B1(n_1002),
.B2(n_989),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_1022),
.A2(n_499),
.B1(n_486),
.B2(n_882),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1045),
.B(n_887),
.Y(n_1070)
);

AOI22xp33_ASAP7_75t_L g1071 ( 
.A1(n_1047),
.A2(n_499),
.B1(n_486),
.B2(n_761),
.Y(n_1071)
);

AOI22xp33_ASAP7_75t_L g1072 ( 
.A1(n_1048),
.A2(n_499),
.B1(n_977),
.B2(n_895),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_SL g1073 ( 
.A1(n_1016),
.A2(n_829),
.B(n_793),
.Y(n_1073)
);

AOI22xp33_ASAP7_75t_L g1074 ( 
.A1(n_1060),
.A2(n_499),
.B1(n_829),
.B2(n_793),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_SL g1075 ( 
.A1(n_1052),
.A2(n_1002),
.B1(n_999),
.B2(n_1015),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_1041),
.A2(n_1002),
.B1(n_1010),
.B2(n_1015),
.Y(n_1076)
);

AOI22xp33_ASAP7_75t_L g1077 ( 
.A1(n_1056),
.A2(n_793),
.B1(n_1010),
.B2(n_1015),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_1016),
.A2(n_957),
.B1(n_933),
.B2(n_924),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_1021),
.B(n_924),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_1034),
.A2(n_957),
.B1(n_767),
.B2(n_933),
.Y(n_1080)
);

AOI22xp33_ASAP7_75t_L g1081 ( 
.A1(n_1025),
.A2(n_767),
.B1(n_841),
.B2(n_834),
.Y(n_1081)
);

OAI22xp33_ASAP7_75t_L g1082 ( 
.A1(n_1049),
.A2(n_558),
.B1(n_554),
.B2(n_845),
.Y(n_1082)
);

AOI22xp33_ASAP7_75t_SL g1083 ( 
.A1(n_1042),
.A2(n_558),
.B1(n_554),
.B2(n_562),
.Y(n_1083)
);

AOI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_1030),
.A2(n_544),
.B1(n_836),
.B2(n_558),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1027),
.Y(n_1085)
);

OAI221xp5_ASAP7_75t_L g1086 ( 
.A1(n_1055),
.A2(n_836),
.B1(n_512),
.B2(n_509),
.C(n_506),
.Y(n_1086)
);

OAI22x1_ASAP7_75t_L g1087 ( 
.A1(n_1046),
.A2(n_1032),
.B1(n_1037),
.B2(n_1031),
.Y(n_1087)
);

AOI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_1018),
.A2(n_825),
.B1(n_811),
.B2(n_805),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1040),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_1043),
.A2(n_825),
.B1(n_512),
.B2(n_509),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_1051),
.A2(n_811),
.B1(n_513),
.B2(n_512),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_1029),
.A2(n_506),
.B1(n_495),
.B2(n_513),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_1061),
.A2(n_513),
.B1(n_29),
.B2(n_30),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1028),
.B(n_28),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1017),
.B(n_30),
.Y(n_1095)
);

AOI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_1063),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_1053),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1019),
.B(n_37),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_1035),
.Y(n_1099)
);

OAI221xp5_ASAP7_75t_L g1100 ( 
.A1(n_1058),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.C(n_42),
.Y(n_1100)
);

AOI221xp5_ASAP7_75t_L g1101 ( 
.A1(n_1024),
.A2(n_42),
.B1(n_43),
.B2(n_46),
.C(n_47),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1035),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_1064),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_1103)
);

OAI222xp33_ASAP7_75t_L g1104 ( 
.A1(n_1026),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.C1(n_53),
.C2(n_54),
.Y(n_1104)
);

AOI22xp33_ASAP7_75t_L g1105 ( 
.A1(n_1033),
.A2(n_56),
.B1(n_73),
.B2(n_74),
.Y(n_1105)
);

AOI221xp5_ASAP7_75t_L g1106 ( 
.A1(n_1036),
.A2(n_56),
.B1(n_75),
.B2(n_78),
.C(n_81),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1050),
.A2(n_289),
.B1(n_90),
.B2(n_91),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1062),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_1054),
.A2(n_89),
.B1(n_93),
.B2(n_95),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_1050),
.A2(n_288),
.B1(n_98),
.B2(n_101),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1101),
.A2(n_1039),
.B(n_1038),
.Y(n_1111)
);

NAND2xp33_ASAP7_75t_L g1112 ( 
.A(n_1107),
.B(n_1057),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1108),
.B(n_1079),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1085),
.B(n_1062),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_1075),
.B(n_1023),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1100),
.A2(n_1059),
.B1(n_1023),
.B2(n_1065),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_1067),
.B(n_113),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1089),
.B(n_114),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1087),
.B(n_117),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1070),
.B(n_1095),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1073),
.B(n_121),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_1099),
.B(n_122),
.Y(n_1122)
);

OAI21xp33_ASAP7_75t_L g1123 ( 
.A1(n_1096),
.A2(n_132),
.B(n_133),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1098),
.B(n_134),
.Y(n_1124)
);

OAI21xp5_ASAP7_75t_SL g1125 ( 
.A1(n_1103),
.A2(n_135),
.B(n_137),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1094),
.B(n_1077),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_1083),
.B(n_139),
.Y(n_1127)
);

NAND3xp33_ASAP7_75t_L g1128 ( 
.A(n_1106),
.B(n_140),
.C(n_141),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_1076),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1069),
.B(n_144),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1068),
.B(n_145),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1069),
.B(n_146),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1107),
.B(n_153),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1102),
.B(n_155),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1066),
.B(n_156),
.Y(n_1135)
);

OAI31xp33_ASAP7_75t_L g1136 ( 
.A1(n_1104),
.A2(n_1097),
.A3(n_1093),
.B(n_1091),
.Y(n_1136)
);

NAND3xp33_ASAP7_75t_SL g1137 ( 
.A(n_1110),
.B(n_158),
.C(n_159),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1080),
.B(n_161),
.Y(n_1138)
);

NAND3xp33_ASAP7_75t_L g1139 ( 
.A(n_1105),
.B(n_162),
.C(n_163),
.Y(n_1139)
);

NAND3xp33_ASAP7_75t_L g1140 ( 
.A(n_1109),
.B(n_164),
.C(n_165),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_1082),
.B(n_1078),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1084),
.B(n_166),
.Y(n_1142)
);

OAI221xp5_ASAP7_75t_SL g1143 ( 
.A1(n_1086),
.A2(n_170),
.B1(n_176),
.B2(n_177),
.C(n_180),
.Y(n_1143)
);

OAI221xp5_ASAP7_75t_SL g1144 ( 
.A1(n_1092),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.C(n_188),
.Y(n_1144)
);

NAND4xp25_ASAP7_75t_L g1145 ( 
.A(n_1072),
.B(n_190),
.C(n_193),
.D(n_196),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_1114),
.B(n_1113),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1114),
.B(n_1081),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1120),
.Y(n_1148)
);

NAND3xp33_ASAP7_75t_L g1149 ( 
.A(n_1135),
.B(n_1074),
.C(n_1090),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1118),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1118),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1119),
.Y(n_1152)
);

NOR3xp33_ASAP7_75t_L g1153 ( 
.A(n_1125),
.B(n_1088),
.C(n_1071),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1129),
.B(n_1126),
.Y(n_1154)
);

OAI211xp5_ASAP7_75t_SL g1155 ( 
.A1(n_1124),
.A2(n_1136),
.B(n_1111),
.C(n_1141),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1119),
.B(n_199),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1141),
.B(n_201),
.Y(n_1157)
);

NAND3xp33_ASAP7_75t_L g1158 ( 
.A(n_1128),
.B(n_203),
.C(n_206),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1121),
.B(n_208),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_1122),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1122),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1121),
.B(n_215),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_L g1163 ( 
.A(n_1115),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1117),
.B(n_217),
.Y(n_1164)
);

NOR3xp33_ASAP7_75t_L g1165 ( 
.A(n_1137),
.B(n_222),
.C(n_226),
.Y(n_1165)
);

NOR3xp33_ASAP7_75t_L g1166 ( 
.A(n_1140),
.B(n_228),
.C(n_229),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_1146),
.Y(n_1167)
);

NAND4xp25_ASAP7_75t_L g1168 ( 
.A(n_1155),
.B(n_1116),
.C(n_1143),
.D(n_1123),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1152),
.B(n_1112),
.Y(n_1169)
);

OA22x2_ASAP7_75t_L g1170 ( 
.A1(n_1163),
.A2(n_1133),
.B1(n_1127),
.B2(n_1131),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1146),
.B(n_1112),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1146),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1148),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_1160),
.Y(n_1174)
);

OR2x2_ASAP7_75t_L g1175 ( 
.A(n_1154),
.B(n_1134),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_1150),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1150),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_1160),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1151),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1160),
.B(n_1132),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1151),
.Y(n_1181)
);

NAND4xp75_ASAP7_75t_SL g1182 ( 
.A(n_1157),
.B(n_1130),
.C(n_1132),
.D(n_1138),
.Y(n_1182)
);

INVx2_ASAP7_75t_SL g1183 ( 
.A(n_1161),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1176),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1167),
.B(n_1147),
.Y(n_1185)
);

INVx2_ASAP7_75t_SL g1186 ( 
.A(n_1167),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1173),
.B(n_1147),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1176),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1177),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1179),
.Y(n_1190)
);

XNOR2xp5_ASAP7_75t_L g1191 ( 
.A(n_1182),
.B(n_1156),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1181),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1172),
.Y(n_1193)
);

INVx2_ASAP7_75t_SL g1194 ( 
.A(n_1185),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_1186),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1189),
.Y(n_1196)
);

OA22x2_ASAP7_75t_L g1197 ( 
.A1(n_1191),
.A2(n_1171),
.B1(n_1169),
.B2(n_1178),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1190),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1192),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_1187),
.Y(n_1200)
);

OA22x2_ASAP7_75t_L g1201 ( 
.A1(n_1193),
.A2(n_1171),
.B1(n_1169),
.B2(n_1180),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1184),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_1188),
.B(n_1175),
.Y(n_1203)
);

OAI22x1_ASAP7_75t_SL g1204 ( 
.A1(n_1184),
.A2(n_1183),
.B1(n_1170),
.B2(n_1168),
.Y(n_1204)
);

INVx2_ASAP7_75t_SL g1205 ( 
.A(n_1195),
.Y(n_1205)
);

INVxp67_ASAP7_75t_L g1206 ( 
.A(n_1204),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1196),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1194),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1196),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1199),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_1202),
.Y(n_1211)
);

INVx1_ASAP7_75t_SL g1212 ( 
.A(n_1197),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1206),
.A2(n_1201),
.B1(n_1200),
.B2(n_1203),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1211),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1207),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1212),
.A2(n_1198),
.B1(n_1174),
.B2(n_1159),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1205),
.A2(n_1208),
.B1(n_1210),
.B2(n_1209),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1214),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1213),
.A2(n_1174),
.B1(n_1158),
.B2(n_1149),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1215),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1216),
.A2(n_1159),
.B1(n_1162),
.B2(n_1164),
.Y(n_1221)
);

NAND4xp25_ASAP7_75t_SL g1222 ( 
.A(n_1217),
.B(n_1166),
.C(n_1153),
.D(n_1165),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1218),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1220),
.Y(n_1224)
);

OA22x2_ASAP7_75t_L g1225 ( 
.A1(n_1219),
.A2(n_1142),
.B1(n_1144),
.B2(n_1145),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1221),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_1222),
.B(n_1139),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1224),
.B(n_231),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1225),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1226),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1227),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1223),
.Y(n_1232)
);

NOR2x1_ASAP7_75t_L g1233 ( 
.A(n_1228),
.B(n_1231),
.Y(n_1233)
);

NOR3xp33_ASAP7_75t_SL g1234 ( 
.A(n_1230),
.B(n_238),
.C(n_239),
.Y(n_1234)
);

OAI22x1_ASAP7_75t_L g1235 ( 
.A1(n_1229),
.A2(n_241),
.B1(n_243),
.B2(n_244),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_SL g1236 ( 
.A1(n_1232),
.A2(n_245),
.B(n_249),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1233),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1235),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1234),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1236),
.Y(n_1240)
);

INVx1_ASAP7_75t_SL g1241 ( 
.A(n_1237),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1238),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1239),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_1240),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1242),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1243),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1244),
.Y(n_1247)
);

AOI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1247),
.A2(n_1241),
.B1(n_1228),
.B2(n_255),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1246),
.A2(n_252),
.B1(n_254),
.B2(n_257),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1245),
.A2(n_258),
.B1(n_262),
.B2(n_267),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1248),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_SL g1252 ( 
.A1(n_1251),
.A2(n_1249),
.B1(n_1250),
.B2(n_273),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1252),
.Y(n_1253)
);

AOI221x1_ASAP7_75t_L g1254 ( 
.A1(n_1253),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.C(n_279),
.Y(n_1254)
);

AOI211xp5_ASAP7_75t_L g1255 ( 
.A1(n_1254),
.A2(n_280),
.B(n_283),
.C(n_285),
.Y(n_1255)
);


endmodule