module fake_jpeg_13554_n_520 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_520);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_520;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_8),
.B(n_4),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_20),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_52),
.B(n_60),
.Y(n_105)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_55),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_20),
.B(n_17),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_61),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_63),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_31),
.B(n_17),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_70),
.Y(n_109)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_65),
.Y(n_116)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_67),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_68),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_69),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_72),
.Y(n_152)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

BUFx24_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_40),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_80),
.Y(n_114)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

BUFx4f_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_78),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_44),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g120 ( 
.A(n_81),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_40),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_89),
.B(n_96),
.Y(n_127)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_0),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_30),
.Y(n_128)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_31),
.B(n_0),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_32),
.B(n_0),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_97),
.B(n_99),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_40),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_40),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_100),
.B(n_33),
.Y(n_143)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_26),
.Y(n_101)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_L g102 ( 
.A1(n_94),
.A2(n_37),
.B1(n_41),
.B2(n_36),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_102),
.A2(n_124),
.B1(n_56),
.B2(n_63),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_30),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_103),
.B(n_141),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_67),
.A2(n_21),
.B1(n_45),
.B2(n_43),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_113),
.A2(n_154),
.B1(n_37),
.B2(n_45),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_49),
.B1(n_45),
.B2(n_21),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_65),
.B(n_30),
.C(n_43),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_126),
.B(n_39),
.C(n_28),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_143),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_93),
.B(n_33),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_58),
.B(n_32),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_151),
.B(n_50),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_51),
.A2(n_45),
.B1(n_21),
.B2(n_48),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_61),
.Y(n_156)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_75),
.Y(n_157)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_73),
.Y(n_159)
);

INVx11_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_112),
.Y(n_161)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_161),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_48),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_162),
.Y(n_244)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_163),
.Y(n_238)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_164),
.Y(n_233)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_117),
.Y(n_165)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_165),
.Y(n_234)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_167),
.Y(n_243)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_112),
.Y(n_168)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_168),
.Y(n_219)
);

NAND2xp33_ASAP7_75t_SL g170 ( 
.A(n_103),
.B(n_69),
.Y(n_170)
);

AND2x4_ASAP7_75t_SL g217 ( 
.A(n_170),
.B(n_104),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_127),
.B(n_48),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_171),
.B(n_172),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_114),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_173),
.A2(n_196),
.B1(n_142),
.B2(n_139),
.Y(n_251)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_116),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_174),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_175),
.B(n_179),
.C(n_204),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_106),
.A2(n_59),
.B1(n_77),
.B2(n_85),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_176),
.A2(n_190),
.B1(n_191),
.B2(n_202),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_137),
.B(n_101),
.C(n_76),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_180),
.Y(n_220)
);

CKINVDCx12_ASAP7_75t_R g181 ( 
.A(n_108),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_181),
.Y(n_258)
);

BUFx12f_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_182),
.Y(n_230)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_183),
.Y(n_221)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_184),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g185 ( 
.A(n_118),
.Y(n_185)
);

BUFx16f_ASAP7_75t_L g256 ( 
.A(n_185),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_109),
.B(n_38),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_210),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_187),
.A2(n_209),
.B1(n_139),
.B2(n_152),
.Y(n_227)
);

CKINVDCx12_ASAP7_75t_R g188 ( 
.A(n_111),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_188),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_122),
.B(n_90),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_189),
.B(n_197),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_106),
.A2(n_37),
.B1(n_33),
.B2(n_58),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_133),
.A2(n_34),
.B1(n_39),
.B2(n_28),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_114),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_192),
.Y(n_250)
);

INVx11_ASAP7_75t_L g193 ( 
.A(n_130),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_193),
.Y(n_225)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_125),
.Y(n_194)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_138),
.Y(n_195)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_L g196 ( 
.A1(n_102),
.A2(n_86),
.B1(n_72),
.B2(n_71),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_141),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_148),
.A2(n_134),
.B1(n_115),
.B2(n_120),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_198),
.A2(n_205),
.B1(n_152),
.B2(n_145),
.Y(n_246)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_138),
.Y(n_199)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_199),
.Y(n_235)
);

CKINVDCx12_ASAP7_75t_R g200 ( 
.A(n_138),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_200),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_129),
.A2(n_18),
.B1(n_34),
.B2(n_38),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_109),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_203),
.B(n_207),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_136),
.B(n_55),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_120),
.A2(n_62),
.B1(n_83),
.B2(n_81),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_118),
.Y(n_206)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_206),
.Y(n_240)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_150),
.Y(n_208)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_208),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_135),
.A2(n_68),
.B1(n_79),
.B2(n_18),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_105),
.B(n_50),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_116),
.Y(n_211)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_211),
.Y(n_255)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_132),
.Y(n_212)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_212),
.Y(n_261)
);

BUFx12f_ASAP7_75t_L g213 ( 
.A(n_132),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_214),
.Y(n_252)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_110),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_105),
.B(n_47),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_215),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_110),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_216),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_217),
.B(n_204),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_227),
.A2(n_246),
.B1(n_263),
.B2(n_212),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_192),
.A2(n_130),
.B1(n_131),
.B2(n_119),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_229),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_160),
.B(n_121),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_232),
.B(n_239),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_175),
.B(n_144),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_196),
.A2(n_135),
.B1(n_145),
.B2(n_142),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_249),
.A2(n_251),
.B1(n_254),
.B2(n_260),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_187),
.A2(n_153),
.B1(n_47),
.B2(n_129),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_201),
.B(n_130),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_194),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_201),
.A2(n_123),
.B1(n_107),
.B2(n_41),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_186),
.B(n_0),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_264),
.Y(n_288)
);

OAI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_189),
.A2(n_21),
.B1(n_41),
.B2(n_36),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_179),
.B(n_1),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_221),
.Y(n_265)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_265),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_242),
.B(n_210),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_266),
.B(n_268),
.Y(n_344)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_221),
.Y(n_267)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_267),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_228),
.B(n_183),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_252),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_269),
.B(n_270),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_250),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_224),
.Y(n_271)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_271),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_273),
.A2(n_193),
.B(n_241),
.Y(n_317)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_222),
.Y(n_274)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_274),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_245),
.B(n_177),
.Y(n_277)
);

OAI21xp33_ASAP7_75t_L g327 ( 
.A1(n_277),
.A2(n_305),
.B(n_287),
.Y(n_327)
);

A2O1A1Ixp33_ASAP7_75t_L g278 ( 
.A1(n_239),
.A2(n_201),
.B(n_170),
.C(n_204),
.Y(n_278)
);

O2A1O1Ixp33_ASAP7_75t_L g311 ( 
.A1(n_278),
.A2(n_299),
.B(n_217),
.C(n_257),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_279),
.B(n_98),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_231),
.Y(n_280)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_280),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_218),
.B(n_166),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_281),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_218),
.B(n_169),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_282),
.Y(n_335)
);

INVx8_ASAP7_75t_L g283 ( 
.A(n_224),
.Y(n_283)
);

INVx5_ASAP7_75t_L g323 ( 
.A(n_283),
.Y(n_323)
);

INVx8_ASAP7_75t_L g284 ( 
.A(n_238),
.Y(n_284)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_284),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_247),
.A2(n_165),
.B(n_164),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_285),
.A2(n_167),
.B(n_178),
.Y(n_332)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_222),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_286),
.B(n_287),
.Y(n_316)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_255),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_229),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g319 ( 
.A1(n_289),
.A2(n_292),
.B1(n_234),
.B2(n_214),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_290),
.A2(n_244),
.B1(n_240),
.B2(n_225),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_264),
.B(n_180),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_291),
.B(n_295),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_217),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_255),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_293),
.A2(n_297),
.B1(n_301),
.B2(n_234),
.Y(n_331)
);

INVx13_ASAP7_75t_L g294 ( 
.A(n_259),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_294),
.Y(n_347)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_220),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_253),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_296),
.B(n_298),
.Y(n_340)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_231),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_253),
.Y(n_298)
);

AO22x2_ASAP7_75t_SL g299 ( 
.A1(n_251),
.A2(n_198),
.B1(n_178),
.B2(n_205),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_220),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_300),
.B(n_302),
.Y(n_341)
);

BUFx12f_ASAP7_75t_L g301 ( 
.A(n_241),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_261),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_248),
.B(n_236),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_303),
.B(n_304),
.Y(n_342)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_261),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_248),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_238),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_306),
.B(n_307),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_232),
.B(n_163),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_237),
.A2(n_161),
.B1(n_168),
.B2(n_206),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_240),
.B1(n_225),
.B2(n_219),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_290),
.A2(n_236),
.B1(n_260),
.B2(n_246),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_310),
.A2(n_314),
.B1(n_325),
.B2(n_329),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g363 ( 
.A(n_311),
.B(n_319),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_312),
.A2(n_333),
.B1(n_334),
.B2(n_284),
.Y(n_356)
);

OA21x2_ASAP7_75t_L g313 ( 
.A1(n_276),
.A2(n_235),
.B(n_226),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_313),
.B(n_337),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_317),
.B(n_346),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_273),
.A2(n_244),
.B(n_223),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_322),
.A2(n_328),
.B(n_332),
.Y(n_374)
);

AOI32xp33_ASAP7_75t_L g324 ( 
.A1(n_303),
.A2(n_275),
.A3(n_276),
.B1(n_278),
.B2(n_273),
.Y(n_324)
);

FAx1_ASAP7_75t_SL g382 ( 
.A(n_324),
.B(n_256),
.CI(n_78),
.CON(n_382),
.SN(n_382)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_275),
.A2(n_223),
.B1(n_262),
.B2(n_219),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_327),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_285),
.A2(n_235),
.B(n_226),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_299),
.A2(n_184),
.B1(n_185),
.B2(n_213),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_331),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_299),
.A2(n_233),
.B1(n_243),
.B2(n_230),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_272),
.A2(n_233),
.B1(n_243),
.B2(n_195),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_291),
.A2(n_288),
.B1(n_279),
.B2(n_267),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_288),
.A2(n_185),
.B1(n_213),
.B2(n_41),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_338),
.B(n_343),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_286),
.A2(n_182),
.B1(n_199),
.B2(n_230),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_296),
.B(n_258),
.C(n_174),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_345),
.B(n_295),
.C(n_294),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_326),
.Y(n_349)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_349),
.Y(n_408)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_316),
.Y(n_350)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_350),
.Y(n_387)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_316),
.Y(n_351)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_351),
.Y(n_395)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_340),
.Y(n_352)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_352),
.Y(n_401)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_340),
.Y(n_354)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_354),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_318),
.B(n_301),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_355),
.B(n_362),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_356),
.A2(n_371),
.B1(n_378),
.B2(n_381),
.Y(n_411)
);

BUFx12_ASAP7_75t_L g357 ( 
.A(n_347),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_357),
.Y(n_385)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_341),
.Y(n_360)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_360),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_318),
.B(n_301),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_361),
.B(n_367),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_344),
.B(n_335),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_341),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_364),
.B(n_370),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_324),
.B(n_298),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_365),
.B(n_375),
.C(n_346),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_335),
.B(n_300),
.Y(n_367)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_315),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_342),
.A2(n_265),
.B1(n_274),
.B2(n_302),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_321),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_372),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_339),
.B(n_304),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_373),
.B(n_377),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_325),
.B(n_283),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_376),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_339),
.B(n_280),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_342),
.A2(n_271),
.B1(n_297),
.B2(n_306),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_315),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_379),
.B(n_380),
.Y(n_391)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_326),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_334),
.A2(n_182),
.B1(n_256),
.B2(n_78),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_382),
.A2(n_313),
.B(n_345),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_369),
.B(n_309),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_383),
.B(n_397),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_384),
.B(n_378),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_368),
.A2(n_328),
.B1(n_312),
.B2(n_332),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_388),
.A2(n_389),
.B1(n_390),
.B2(n_407),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_368),
.A2(n_311),
.B1(n_310),
.B2(n_314),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_359),
.A2(n_329),
.B1(n_348),
.B2(n_337),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_371),
.B(n_350),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_394),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_396),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_374),
.A2(n_348),
.B(n_317),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_358),
.B(n_322),
.C(n_313),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_398),
.B(n_403),
.C(n_384),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_374),
.A2(n_347),
.B(n_336),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_400),
.B(n_406),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_358),
.B(n_320),
.C(n_321),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_359),
.B(n_323),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_351),
.A2(n_336),
.B1(n_323),
.B2(n_320),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_352),
.B(n_338),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_409),
.B(n_2),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_354),
.A2(n_330),
.B1(n_343),
.B2(n_256),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_410),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_392),
.A2(n_363),
.B1(n_353),
.B2(n_360),
.Y(n_413)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_413),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_415),
.B(n_419),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_403),
.B(n_365),
.C(n_375),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_416),
.B(n_417),
.C(n_431),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_398),
.B(n_364),
.C(n_363),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_396),
.B(n_382),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_420),
.B(n_424),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_392),
.A2(n_366),
.B1(n_373),
.B2(n_379),
.Y(n_422)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_422),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_402),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_423),
.B(n_426),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_397),
.B(n_382),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_402),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_389),
.B(n_377),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_427),
.B(n_388),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_399),
.A2(n_366),
.B1(n_370),
.B2(n_380),
.Y(n_428)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_428),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_411),
.A2(n_349),
.B1(n_357),
.B2(n_372),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_430),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_387),
.B(n_349),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_412),
.B(n_330),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_432),
.B(n_434),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_387),
.B(n_357),
.C(n_381),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_433),
.B(n_436),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_412),
.B(n_2),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_435),
.A2(n_401),
.B1(n_395),
.B2(n_404),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_395),
.B(n_401),
.C(n_404),
.Y(n_436)
);

CKINVDCx14_ASAP7_75t_R g446 ( 
.A(n_437),
.Y(n_446)
);

XNOR2x2_ASAP7_75t_SL g439 ( 
.A(n_419),
.B(n_394),
.Y(n_439)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_439),
.Y(n_469)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_442),
.Y(n_473)
);

AOI21xp33_ASAP7_75t_L g445 ( 
.A1(n_414),
.A2(n_385),
.B(n_405),
.Y(n_445)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_445),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_448),
.B(n_424),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_431),
.B(n_400),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_451),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_421),
.A2(n_390),
.B1(n_405),
.B2(n_407),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_453),
.A2(n_425),
.B1(n_429),
.B2(n_411),
.Y(n_461)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_427),
.Y(n_454)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_454),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_436),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_455),
.B(n_457),
.Y(n_474)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_420),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_418),
.A2(n_386),
.B1(n_410),
.B2(n_391),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_458),
.A2(n_453),
.B1(n_425),
.B2(n_438),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_459),
.B(n_467),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_461),
.A2(n_452),
.B1(n_442),
.B2(n_446),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_462),
.A2(n_466),
.B1(n_437),
.B2(n_408),
.Y(n_483)
);

BUFx24_ASAP7_75t_SL g463 ( 
.A(n_444),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_463),
.B(n_470),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_451),
.A2(n_417),
.B(n_433),
.Y(n_464)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_464),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_449),
.A2(n_435),
.B1(n_409),
.B2(n_385),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_451),
.A2(n_386),
.B(n_391),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_441),
.B(n_415),
.C(n_416),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_468),
.B(n_471),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_458),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_441),
.B(n_408),
.C(n_393),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_471),
.Y(n_476)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_476),
.Y(n_494)
);

AOI22x1_ASAP7_75t_SL g477 ( 
.A1(n_469),
.A2(n_448),
.B1(n_450),
.B2(n_439),
.Y(n_477)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_477),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_468),
.B(n_447),
.C(n_456),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_479),
.B(n_481),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_480),
.B(n_483),
.Y(n_493)
);

FAx1_ASAP7_75t_SL g481 ( 
.A(n_467),
.B(n_464),
.CI(n_460),
.CON(n_481),
.SN(n_481)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_474),
.B(n_456),
.C(n_457),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_482),
.B(n_484),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_472),
.B(n_440),
.C(n_443),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_472),
.B(n_440),
.C(n_473),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_487),
.B(n_488),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_461),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_488)
);

NOR2xp67_ASAP7_75t_R g490 ( 
.A(n_484),
.B(n_469),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_490),
.B(n_8),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_485),
.A2(n_473),
.B1(n_465),
.B2(n_459),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_491),
.B(n_492),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_486),
.B(n_465),
.C(n_7),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_479),
.A2(n_5),
.B(n_7),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_497),
.A2(n_477),
.B(n_475),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g499 ( 
.A1(n_478),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g503 ( 
.A(n_499),
.Y(n_503)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_500),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_495),
.A2(n_482),
.B(n_487),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_501),
.B(n_505),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_489),
.B(n_481),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_502),
.B(n_493),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_494),
.A2(n_496),
.B(n_498),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_506),
.B(n_499),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_508),
.B(n_510),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_509),
.B(n_504),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_512),
.A2(n_513),
.B1(n_511),
.B2(n_503),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_507),
.A2(n_493),
.B(n_492),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_514),
.B(n_515),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_511),
.B(n_10),
.Y(n_515)
);

AOI322xp5_ASAP7_75t_L g517 ( 
.A1(n_516),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_515),
.C2(n_514),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_517),
.B(n_11),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_518),
.B(n_13),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_519),
.A2(n_13),
.B(n_11),
.Y(n_520)
);


endmodule