module fake_jpeg_18006_n_347 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_347);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_347;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx8_ASAP7_75t_SL g20 ( 
.A(n_8),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_37),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_49),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_30),
.Y(n_49)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_62),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_30),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_33),
.Y(n_76)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx5_ASAP7_75t_SL g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_31),
.Y(n_63)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_47),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_48),
.B1(n_43),
.B2(n_38),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_69),
.A2(n_74),
.B1(n_86),
.B2(n_100),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_40),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_70),
.B(n_98),
.Y(n_114)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_48),
.B1(n_43),
.B2(n_40),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_45),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_75),
.B(n_77),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_76),
.B(n_90),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_49),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_80),
.B(n_82),
.Y(n_129)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

OAI32xp33_ASAP7_75t_L g83 ( 
.A1(n_58),
.A2(n_23),
.A3(n_19),
.B1(n_31),
.B2(n_24),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_83),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_58),
.B(n_23),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_85),
.B(n_88),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_67),
.A2(n_48),
.B1(n_43),
.B2(n_39),
.Y(n_86)
);

AND2x4_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_42),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_87),
.A2(n_26),
.B(n_25),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_61),
.B(n_19),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_68),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_56),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVxp33_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVxp33_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_65),
.B(n_34),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_97),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_42),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_51),
.A2(n_18),
.B1(n_33),
.B2(n_37),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_99),
.A2(n_109),
.B1(n_32),
.B2(n_29),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_66),
.A2(n_18),
.B1(n_24),
.B2(n_25),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_101),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_59),
.B(n_42),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_103),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_55),
.B(n_26),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_53),
.A2(n_41),
.B1(n_47),
.B2(n_44),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_105),
.A2(n_35),
.B1(n_32),
.B2(n_29),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_63),
.B(n_36),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_21),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_54),
.A2(n_41),
.B1(n_18),
.B2(n_47),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_107),
.A2(n_108),
.B1(n_34),
.B2(n_28),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_54),
.A2(n_41),
.B1(n_37),
.B2(n_34),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g110 ( 
.A1(n_53),
.A2(n_44),
.B1(n_28),
.B2(n_46),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_111),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_53),
.A2(n_44),
.B1(n_28),
.B2(n_35),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_112),
.A2(n_120),
.B1(n_132),
.B2(n_109),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_17),
.B1(n_35),
.B2(n_32),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_70),
.B(n_36),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_131),
.C(n_87),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_77),
.Y(n_153)
);

AO21x1_ASAP7_75t_L g164 ( 
.A1(n_130),
.A2(n_138),
.B(n_110),
.Y(n_164)
);

AND2x2_ASAP7_75t_SL g131 ( 
.A(n_87),
.B(n_84),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_76),
.B(n_35),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_110),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_76),
.A2(n_20),
.B(n_1),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_140),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_87),
.B(n_0),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_141),
.A2(n_104),
.B1(n_75),
.B2(n_96),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_144),
.B(n_145),
.Y(n_200)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_114),
.B(n_84),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_158),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_136),
.Y(n_147)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_148),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_149),
.B(n_156),
.Y(n_176)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_150),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_151),
.A2(n_155),
.B(n_121),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_152),
.Y(n_196)
);

NAND3xp33_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_113),
.C(n_137),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_154),
.A2(n_160),
.B1(n_169),
.B2(n_125),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_119),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_98),
.C(n_102),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_162),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_83),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_79),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_159),
.B(n_164),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_118),
.A2(n_104),
.B1(n_71),
.B2(n_69),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_72),
.C(n_81),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_78),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_166),
.Y(n_190)
);

AO21x1_ASAP7_75t_L g165 ( 
.A1(n_135),
.A2(n_110),
.B(n_111),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_165),
.A2(n_170),
.B(n_141),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_122),
.B(n_131),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_89),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_138),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_135),
.A2(n_91),
.B1(n_92),
.B2(n_95),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_168),
.A2(n_120),
.B1(n_112),
.B2(n_123),
.Y(n_177)
);

AO21x2_ASAP7_75t_L g169 ( 
.A1(n_140),
.A2(n_118),
.B(n_69),
.Y(n_169)
);

O2A1O1Ixp33_ASAP7_75t_SL g170 ( 
.A1(n_118),
.A2(n_111),
.B(n_69),
.C(n_73),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_115),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_171),
.B(n_117),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_172),
.A2(n_202),
.B1(n_203),
.B2(n_168),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_118),
.B(n_141),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_173),
.A2(n_175),
.B(n_184),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_177),
.A2(n_179),
.B1(n_182),
.B2(n_195),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_161),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_178),
.B(n_194),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_169),
.A2(n_140),
.B1(n_125),
.B2(n_134),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_169),
.A2(n_141),
.B1(n_126),
.B2(n_113),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_166),
.A2(n_126),
.B(n_124),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_124),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_162),
.C(n_155),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_187),
.A2(n_197),
.B(n_199),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_145),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_192),
.B(n_147),
.Y(n_225)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_148),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_169),
.A2(n_123),
.B1(n_121),
.B2(n_132),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_169),
.A2(n_130),
.B(n_142),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_159),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_169),
.A2(n_111),
.B1(n_117),
.B2(n_80),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_158),
.A2(n_128),
.B(n_139),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_201),
.A2(n_193),
.B(n_173),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_154),
.A2(n_133),
.B1(n_105),
.B2(n_94),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_149),
.A2(n_133),
.B1(n_136),
.B2(n_139),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_157),
.Y(n_204)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_204),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_207),
.A2(n_209),
.B1(n_216),
.B2(n_218),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_172),
.A2(n_163),
.B1(n_167),
.B2(n_165),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_191),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_210),
.B(n_211),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_191),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_217),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_230),
.C(n_232),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_176),
.A2(n_165),
.B1(n_170),
.B2(n_146),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_189),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_202),
.A2(n_170),
.B1(n_164),
.B2(n_160),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_183),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_219),
.B(n_227),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_196),
.A2(n_164),
.B1(n_153),
.B2(n_156),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_220),
.A2(n_233),
.B1(n_178),
.B2(n_29),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_221),
.B(n_222),
.Y(n_239)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_180),
.Y(n_223)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_223),
.Y(n_246)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_183),
.Y(n_224)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_226),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_174),
.B(n_150),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_231),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_185),
.B(n_145),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_185),
.B(n_136),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_179),
.A2(n_147),
.B1(n_116),
.B2(n_3),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_174),
.B(n_32),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_192),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_186),
.C(n_198),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_237),
.B(n_250),
.C(n_214),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_215),
.A2(n_190),
.B1(n_197),
.B2(n_199),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_238),
.A2(n_242),
.B1(n_255),
.B2(n_233),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_229),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_240),
.B(n_231),
.Y(n_261)
);

OA21x2_ASAP7_75t_L g241 ( 
.A1(n_205),
.A2(n_190),
.B(n_188),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_241),
.B(n_248),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_208),
.A2(n_188),
.B1(n_195),
.B2(n_175),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_206),
.B(n_182),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_249),
.Y(n_265)
);

OA21x2_ASAP7_75t_L g248 ( 
.A1(n_205),
.A2(n_184),
.B(n_177),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_206),
.B(n_201),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_181),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_181),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_216),
.Y(n_267)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_213),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_256),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_280),
.Y(n_292)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_261),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_236),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_270),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_247),
.A2(n_213),
.B1(n_207),
.B2(n_209),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_263),
.A2(n_274),
.B1(n_279),
.B2(n_270),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_267),
.C(n_268),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_222),
.C(n_204),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_269),
.B(n_278),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_208),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_224),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_246),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_235),
.B(n_220),
.C(n_218),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_275),
.C(n_251),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_247),
.A2(n_234),
.B1(n_211),
.B2(n_223),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_237),
.B(n_29),
.C(n_17),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_238),
.A2(n_0),
.B(n_1),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_276),
.A2(n_248),
.B(n_258),
.Y(n_293)
);

NOR4xp25_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_17),
.C(n_10),
.D(n_12),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_277),
.B(n_255),
.Y(n_286)
);

AOI21xp33_ASAP7_75t_L g278 ( 
.A1(n_243),
.A2(n_9),
.B(n_16),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_280),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_281),
.B(n_282),
.Y(n_312)
);

O2A1O1Ixp33_ASAP7_75t_R g282 ( 
.A1(n_272),
.A2(n_248),
.B(n_242),
.C(n_241),
.Y(n_282)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_286),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_289),
.C(n_290),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_250),
.C(n_239),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_239),
.C(n_244),
.Y(n_290)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_291),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_293),
.A2(n_297),
.B(n_274),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_294),
.Y(n_309)
);

A2O1A1O1Ixp25_ASAP7_75t_L g295 ( 
.A1(n_267),
.A2(n_241),
.B(n_249),
.C(n_245),
.D(n_253),
.Y(n_295)
);

OAI221xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_17),
.B1(n_9),
.B2(n_10),
.C(n_7),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_271),
.B(n_245),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_292),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_263),
.A2(n_3),
.B(n_4),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_265),
.B(n_275),
.C(n_273),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_4),
.C(n_5),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_283),
.B(n_285),
.Y(n_299)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_299),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_288),
.B(n_260),
.Y(n_301)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_301),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_265),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_313),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_282),
.A2(n_266),
.B1(n_279),
.B2(n_269),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_306),
.Y(n_318)
);

OAI21xp33_ASAP7_75t_L g304 ( 
.A1(n_295),
.A2(n_266),
.B(n_276),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_304),
.A2(n_297),
.B(n_284),
.Y(n_324)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_305),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_292),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_293),
.C(n_287),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_9),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_311),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_303),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_322),
.C(n_300),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_323),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_300),
.B(n_284),
.C(n_289),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_312),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_324),
.B(n_13),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_319),
.A2(n_321),
.B(n_314),
.Y(n_325)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_325),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_326),
.B(n_331),
.C(n_316),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_317),
.A2(n_307),
.B1(n_310),
.B2(n_304),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_327),
.B(n_329),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_333),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_318),
.A2(n_305),
.B1(n_313),
.B2(n_302),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_8),
.Y(n_330)
);

AOI21xp33_ASAP7_75t_L g334 ( 
.A1(n_330),
.A2(n_13),
.B(n_14),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_322),
.B(n_13),
.C(n_14),
.Y(n_333)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_334),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_332),
.A2(n_316),
.B(n_14),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_336),
.B(n_338),
.C(n_331),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_330),
.B(n_328),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_340),
.A2(n_341),
.B(n_335),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_343),
.A2(n_337),
.B(n_338),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_344),
.A2(n_342),
.B(n_15),
.Y(n_345)
);

BUFx24_ASAP7_75t_SL g346 ( 
.A(n_345),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_15),
.Y(n_347)
);


endmodule