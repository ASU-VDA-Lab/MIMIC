module real_jpeg_5387_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_0),
.A2(n_36),
.B1(n_41),
.B2(n_46),
.Y(n_35)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_0),
.A2(n_46),
.B1(n_108),
.B2(n_110),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_0),
.A2(n_46),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_0),
.A2(n_46),
.B1(n_232),
.B2(n_234),
.Y(n_231)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_2),
.A2(n_50),
.B1(n_51),
.B2(n_55),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_2),
.A2(n_50),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_2),
.A2(n_50),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_2),
.A2(n_37),
.B1(n_50),
.B2(n_276),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_3),
.A2(n_250),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_3),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_3),
.A2(n_295),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_3),
.A2(n_295),
.B1(n_391),
.B2(n_392),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_L g408 ( 
.A1(n_3),
.A2(n_295),
.B1(n_403),
.B2(n_409),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_4),
.B(n_260),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_4),
.A2(n_259),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_4),
.B(n_190),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_4),
.B(n_369),
.C(n_371),
.Y(n_368)
);

OAI22xp33_ASAP7_75t_L g373 ( 
.A1(n_4),
.A2(n_374),
.B1(n_375),
.B2(n_377),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_4),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_4),
.B(n_146),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_4),
.A2(n_25),
.B1(n_314),
.B2(n_420),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_5),
.A2(n_288),
.B1(n_290),
.B2(n_291),
.Y(n_287)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_5),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_5),
.A2(n_280),
.B1(n_290),
.B2(n_306),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_5),
.A2(n_290),
.B1(n_377),
.B2(n_381),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_5),
.A2(n_290),
.B1(n_409),
.B2(n_421),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_6),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_7),
.A2(n_122),
.B1(n_125),
.B2(n_126),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_7),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_7),
.A2(n_61),
.B1(n_125),
.B2(n_182),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_7),
.A2(n_125),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_7),
.A2(n_125),
.B1(n_265),
.B2(n_268),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_8),
.A2(n_109),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_8),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_8),
.A2(n_187),
.B1(n_280),
.B2(n_282),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g396 ( 
.A1(n_8),
.A2(n_187),
.B1(n_397),
.B2(n_400),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_8),
.A2(n_187),
.B1(n_377),
.B2(n_460),
.Y(n_459)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_9),
.Y(n_134)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_10),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_10),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_10),
.Y(n_315)
);

BUFx5_ASAP7_75t_L g337 ( 
.A(n_10),
.Y(n_337)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_11),
.Y(n_93)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_11),
.Y(n_97)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_11),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_11),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g257 ( 
.A(n_11),
.Y(n_257)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_12),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_13),
.Y(n_91)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_13),
.Y(n_94)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_13),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_13),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_13),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_13),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_13),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_13),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_13),
.Y(n_261)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_13),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_14),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_14),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_14),
.A2(n_81),
.B1(n_109),
.B2(n_115),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_14),
.A2(n_81),
.B1(n_168),
.B2(n_171),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_14),
.A2(n_81),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_15),
.Y(n_75)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_506),
.C(n_510),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_504),
.B(n_508),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_494),
.B(n_503),
.Y(n_18)
);

OAI31xp33_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_219),
.A3(n_240),
.B(n_491),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_199),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_21),
.B(n_199),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_118),
.C(n_162),
.Y(n_21)
);

FAx1_ASAP7_75t_SL g359 ( 
.A(n_22),
.B(n_118),
.CI(n_162),
.CON(n_359),
.SN(n_359)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_85),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g218 ( 
.A1(n_23),
.A2(n_24),
.B(n_87),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_47),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_24),
.A2(n_86),
.B1(n_87),
.B2(n_117),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_24),
.A2(n_47),
.B1(n_86),
.B2(n_351),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_33),
.B(n_35),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_25),
.B(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_25),
.A2(n_263),
.B1(n_271),
.B2(n_275),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_25),
.A2(n_275),
.B(n_312),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_25),
.A2(n_174),
.B(n_396),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_25),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_25),
.A2(n_314),
.B1(n_408),
.B2(n_420),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_25),
.A2(n_35),
.B(n_312),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_28),
.Y(n_270)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_28),
.Y(n_403)
);

BUFx5_ASAP7_75t_L g409 ( 
.A(n_28),
.Y(n_409)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_32),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_32),
.Y(n_429)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_35),
.Y(n_175)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_38),
.A2(n_71),
.B1(n_72),
.B2(n_74),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_44),
.Y(n_422)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_45),
.Y(n_399)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_45),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_47),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_58),
.B(n_76),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_49),
.A2(n_59),
.B1(n_77),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g131 ( 
.A1(n_52),
.A2(n_84),
.B1(n_132),
.B2(n_135),
.Y(n_131)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_53),
.Y(n_158)
);

INVx5_ASAP7_75t_L g379 ( 
.A(n_53),
.Y(n_379)
);

INVx6_ASAP7_75t_L g384 ( 
.A(n_53),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_53),
.Y(n_444)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_54),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g376 ( 
.A(n_54),
.Y(n_376)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_58),
.B(n_160),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_58),
.A2(n_154),
.B(n_155),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_58),
.A2(n_76),
.B(n_155),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_58),
.A2(n_154),
.B1(n_160),
.B2(n_181),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_58),
.A2(n_475),
.B(n_476),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_59),
.A2(n_77),
.B1(n_373),
.B2(n_380),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_59),
.A2(n_77),
.B1(n_380),
.B2(n_390),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_59),
.A2(n_77),
.B1(n_390),
.B2(n_459),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_70),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_69),
.Y(n_60)
);

INVx5_ASAP7_75t_L g367 ( 
.A(n_61),
.Y(n_367)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_68),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_69),
.Y(n_391)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_73),
.Y(n_267)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_77),
.Y(n_154)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_78),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_84),
.Y(n_183)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_107),
.B(n_113),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_88),
.B(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_88),
.A2(n_190),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_88),
.A2(n_190),
.B1(n_287),
.B2(n_293),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_88),
.A2(n_107),
.B(n_190),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_89),
.A2(n_186),
.B(n_189),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_89),
.A2(n_116),
.B1(n_301),
.B2(n_303),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_89),
.A2(n_116),
.B1(n_186),
.B2(n_294),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_89),
.A2(n_500),
.B(n_501),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_98),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_99),
.Y(n_306)
);

INVx6_ASAP7_75t_SL g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_106),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_107),
.B(n_190),
.Y(n_189)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_109),
.Y(n_292)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_112),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_113),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_114),
.Y(n_216)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_115),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_116),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_116),
.A2(n_210),
.B(n_215),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_152),
.B(n_161),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_119),
.B(n_152),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_130),
.B1(n_146),
.B2(n_147),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_121),
.A2(n_131),
.B(n_193),
.Y(n_192)
);

OAI32xp33_ASAP7_75t_L g441 ( 
.A1(n_122),
.A2(n_442),
.A3(n_445),
.B1(n_448),
.B2(n_449),
.Y(n_441)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_SL g457 ( 
.A1(n_123),
.A2(n_374),
.B(n_448),
.Y(n_457)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_124),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_124),
.Y(n_285)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_129),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_130),
.B(n_194),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_130),
.A2(n_147),
.B(n_205),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_130),
.A2(n_230),
.B(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_130),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_130),
.A2(n_146),
.B1(n_342),
.B2(n_457),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_130),
.A2(n_146),
.B(n_498),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_136),
.Y(n_130)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_131),
.B(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_131),
.A2(n_305),
.B1(n_308),
.B2(n_309),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_131),
.A2(n_305),
.B1(n_308),
.B2(n_341),
.Y(n_340)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_133),
.Y(n_451)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_140),
.B1(n_143),
.B2(n_144),
.Y(n_136)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_137),
.Y(n_195)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_139),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_139),
.Y(n_255)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_139),
.Y(n_307)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx6_ASAP7_75t_L g447 ( 
.A(n_141),
.Y(n_447)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_142),
.Y(n_145)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_146),
.B(n_194),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_149),
.Y(n_198)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_159),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_153),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_154),
.B(n_374),
.Y(n_418)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_157),
.Y(n_453)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_158),
.Y(n_463)
);

FAx1_ASAP7_75t_SL g199 ( 
.A(n_161),
.B(n_200),
.CI(n_218),
.CON(n_199),
.SN(n_199)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_184),
.C(n_191),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_163),
.B(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_178),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_164),
.A2(n_178),
.B1(n_179),
.B2(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_164),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_174),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_166),
.A2(n_264),
.B(n_337),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_167),
.Y(n_316)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_169),
.Y(n_276)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_170),
.Y(n_173)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_184),
.A2(n_185),
.B1(n_191),
.B2(n_192),
.Y(n_353)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_189),
.B(n_215),
.Y(n_506)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_229),
.Y(n_228)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_197),
.B(n_374),
.Y(n_448)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_199),
.B(n_221),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_209),
.B2(n_217),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_207),
.B2(n_208),
.Y(n_202)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_203),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_203),
.A2(n_208),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_203),
.B(n_227),
.C(n_235),
.Y(n_502)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_204),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_208),
.C(n_209),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_206),
.A2(n_231),
.B(n_308),
.Y(n_326)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_209),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_209),
.A2(n_217),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_209),
.B(n_222),
.C(n_225),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_220),
.A2(n_492),
.B(n_493),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_235),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_231),
.Y(n_498)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_234),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g500 ( 
.A(n_237),
.Y(n_500)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OA21x2_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_360),
.B(n_485),
.Y(n_240)
);

NAND3xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_345),
.C(n_357),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_330),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_243),
.A2(n_487),
.B(n_488),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_318),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_244),
.B(n_318),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_298),
.C(n_310),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_245),
.B(n_344),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_277),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_246),
.B(n_278),
.C(n_286),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_262),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_247),
.B(n_262),
.Y(n_333)
);

OAI32xp33_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_250),
.A3(n_252),
.B1(n_254),
.B2(n_258),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVxp33_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_272),
.Y(n_271)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g371 ( 
.A(n_276),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_286),
.Y(n_277)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_279),
.Y(n_309)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx4_ASAP7_75t_SL g283 ( 
.A(n_284),
.Y(n_283)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_287),
.Y(n_303)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_288),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_298),
.B(n_310),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.C(n_304),
.Y(n_298)
);

FAx1_ASAP7_75t_SL g332 ( 
.A(n_299),
.B(n_300),
.CI(n_304),
.CON(n_332),
.SN(n_332)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_317),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_311),
.B(n_317),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_316),
.Y(n_312)
);

INVx3_ASAP7_75t_SL g313 ( 
.A(n_314),
.Y(n_313)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_319),
.B(n_321),
.C(n_323),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_323),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_329),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_325),
.A2(n_326),
.B1(n_327),
.B2(n_328),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_325),
.B(n_328),
.C(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_327),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_329),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_343),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_331),
.B(n_343),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.C(n_334),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_332),
.B(n_483),
.Y(n_482)
);

BUFx24_ASAP7_75t_SL g511 ( 
.A(n_332),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_333),
.B(n_334),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_338),
.C(n_340),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_335),
.A2(n_336),
.B1(n_338),
.B2(n_339),
.Y(n_470)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g469 ( 
.A(n_340),
.B(n_470),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

A2O1A1O1Ixp25_ASAP7_75t_L g485 ( 
.A1(n_345),
.A2(n_357),
.B(n_486),
.C(n_489),
.D(n_490),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_346),
.B(n_356),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_346),
.B(n_356),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_349),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_347),
.B(n_350),
.C(n_355),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_352),
.B1(n_354),
.B2(n_355),
.Y(n_349)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_350),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_352),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_358),
.B(n_359),
.Y(n_490)
);

BUFx24_ASAP7_75t_SL g512 ( 
.A(n_359),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_480),
.B(n_484),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_362),
.A2(n_465),
.B(n_479),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_363),
.A2(n_437),
.B(n_464),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_364),
.A2(n_404),
.B(n_436),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_385),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_365),
.B(n_385),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_372),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_366),
.B(n_372),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_368),
.Y(n_366)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_374),
.B(n_427),
.Y(n_426)
);

INVx3_ASAP7_75t_SL g375 ( 
.A(n_376),
.Y(n_375)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_384),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_395),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_387),
.A2(n_388),
.B1(n_389),
.B2(n_394),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_387),
.B(n_394),
.C(n_395),
.Y(n_438)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_389),
.Y(n_394)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_396),
.Y(n_411)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx6_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx6_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_416),
.B(n_435),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_415),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_406),
.B(n_415),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_407),
.A2(n_410),
.B1(n_411),
.B2(n_412),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_417),
.A2(n_423),
.B(n_434),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_419),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_418),
.B(n_419),
.Y(n_434)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_424),
.B(n_425),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_426),
.B(n_430),
.Y(n_425)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx8_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx4_ASAP7_75t_SL g431 ( 
.A(n_432),
.Y(n_431)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_439),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_438),
.B(n_439),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_455),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_440),
.B(n_456),
.C(n_458),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_441),
.B(n_454),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_441),
.B(n_454),
.Y(n_473)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx11_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_452),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_458),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_459),
.Y(n_475)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_467),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_466),
.B(n_467),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_468),
.A2(n_469),
.B1(n_471),
.B2(n_472),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_468),
.B(n_474),
.C(n_477),
.Y(n_481)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_473),
.A2(n_474),
.B1(n_477),
.B2(n_478),
.Y(n_472)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_473),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_474),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_482),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_481),
.B(n_482),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_495),
.B(n_496),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_495),
.B(n_496),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_496),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_496),
.B(n_506),
.Y(n_509)
);

FAx1_ASAP7_75t_SL g496 ( 
.A(n_497),
.B(n_499),
.CI(n_502),
.CON(n_496),
.SN(n_496)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_507),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_506),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);


endmodule