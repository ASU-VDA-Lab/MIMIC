module real_aes_8925_n_286 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_286);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_286;
wire n_480;
wire n_476;
wire n_758;
wire n_887;
wire n_436;
wire n_599;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_635;
wire n_792;
wire n_386;
wire n_503;
wire n_673;
wire n_518;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_815;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_289;
wire n_462;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_656;
wire n_316;
wire n_532;
wire n_755;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_527;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_749;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_741;
wire n_314;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
wire n_862;
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_0), .A2(n_241), .B1(n_329), .B2(n_334), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_1), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_2), .A2(n_224), .B1(n_658), .B2(n_762), .Y(n_761) );
XOR2x2_ASAP7_75t_L g796 ( .A(n_3), .B(n_797), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_4), .A2(n_173), .B1(n_433), .B2(n_436), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_5), .A2(n_55), .B1(n_427), .B2(n_600), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_6), .Y(n_455) );
INVx1_ASAP7_75t_L g640 ( .A(n_7), .Y(n_640) );
AOI222xp33_ASAP7_75t_L g809 ( .A1(n_8), .A2(n_25), .B1(n_231), .B2(n_384), .C1(n_496), .C2(n_502), .Y(n_809) );
AOI22xp33_ASAP7_75t_SL g701 ( .A1(n_9), .A2(n_175), .B1(n_357), .B2(n_547), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_10), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_11), .B(n_644), .Y(n_643) );
CKINVDCx20_ASAP7_75t_R g789 ( .A(n_12), .Y(n_789) );
AOI22xp33_ASAP7_75t_SL g675 ( .A1(n_13), .A2(n_98), .B1(n_436), .B2(n_676), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_14), .A2(n_153), .B1(n_676), .B2(n_717), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_15), .A2(n_74), .B1(n_481), .B2(n_804), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_16), .A2(n_204), .B1(n_323), .B2(n_474), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_17), .Y(n_625) );
AOI22xp33_ASAP7_75t_SL g541 ( .A1(n_18), .A2(n_63), .B1(n_329), .B2(n_334), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g301 ( .A1(n_19), .A2(n_302), .B1(n_407), .B2(n_408), .Y(n_301) );
INVx1_ASAP7_75t_L g407 ( .A(n_19), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_20), .A2(n_281), .B1(n_435), .B2(n_535), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_21), .A2(n_87), .B1(n_431), .B2(n_502), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_22), .A2(n_76), .B1(n_414), .B2(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g605 ( .A(n_23), .Y(n_605) );
AO22x2_ASAP7_75t_L g318 ( .A1(n_24), .A2(n_81), .B1(n_310), .B2(n_315), .Y(n_318) );
INVx1_ASAP7_75t_L g828 ( .A(n_24), .Y(n_828) );
AOI222xp33_ASAP7_75t_L g681 ( .A1(n_26), .A2(n_97), .B1(n_122), .B2(n_376), .C1(n_496), .C2(n_523), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g659 ( .A(n_27), .Y(n_659) );
AOI22xp33_ASAP7_75t_SL g730 ( .A1(n_28), .A2(n_194), .B1(n_703), .B2(n_731), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_29), .A2(n_239), .B1(n_505), .B2(n_579), .Y(n_678) );
CKINVDCx20_ASAP7_75t_R g393 ( .A(n_30), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_31), .A2(n_184), .B1(n_449), .B2(n_607), .Y(n_606) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_32), .Y(n_709) );
CKINVDCx20_ASAP7_75t_R g690 ( .A(n_33), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_34), .A2(n_49), .B1(n_544), .B2(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_35), .A2(n_36), .B1(n_600), .B2(n_644), .Y(n_799) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_37), .A2(n_214), .B1(n_362), .B2(n_547), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_38), .A2(n_155), .B1(n_441), .B2(n_572), .Y(n_669) );
AO22x2_ASAP7_75t_L g320 ( .A1(n_39), .A2(n_83), .B1(n_310), .B2(n_311), .Y(n_320) );
INVx1_ASAP7_75t_L g829 ( .A(n_39), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_40), .A2(n_130), .B1(n_656), .B2(n_658), .Y(n_655) );
AOI211xp5_ASAP7_75t_L g286 ( .A1(n_41), .A2(n_287), .B(n_296), .C(n_830), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g365 ( .A(n_42), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_43), .A2(n_73), .B1(n_441), .B2(n_758), .Y(n_757) );
AOI22xp33_ASAP7_75t_SL g508 ( .A1(n_44), .A2(n_47), .B1(n_509), .B2(n_510), .Y(n_508) );
AOI22xp33_ASAP7_75t_SL g504 ( .A1(n_45), .A2(n_112), .B1(n_481), .B2(n_505), .Y(n_504) );
AOI22xp33_ASAP7_75t_SL g881 ( .A1(n_46), .A2(n_216), .B1(n_439), .B2(n_656), .Y(n_881) );
AOI22xp33_ASAP7_75t_SL g495 ( .A1(n_48), .A2(n_273), .B1(n_376), .B2(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_50), .B(n_600), .Y(n_693) );
INVx1_ASAP7_75t_L g581 ( .A(n_51), .Y(n_581) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_52), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_53), .A2(n_86), .B1(n_356), .B2(n_359), .Y(n_355) );
AOI22xp5_ASAP7_75t_SL g590 ( .A1(n_54), .A2(n_270), .B1(n_591), .B2(n_593), .Y(n_590) );
AOI22xp33_ASAP7_75t_SL g506 ( .A1(n_56), .A2(n_199), .B1(n_334), .B2(n_419), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_57), .Y(n_777) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_58), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_59), .A2(n_240), .B1(n_351), .B2(n_420), .Y(n_856) );
CKINVDCx20_ASAP7_75t_R g873 ( .A(n_60), .Y(n_873) );
XOR2x2_ASAP7_75t_L g490 ( .A(n_61), .B(n_491), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_62), .A2(n_261), .B1(n_376), .B2(n_496), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_64), .B(n_846), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_65), .A2(n_238), .B1(n_550), .B2(n_633), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_66), .A2(n_262), .B1(n_535), .B2(n_602), .Y(n_601) );
AOI22xp33_ASAP7_75t_SL g641 ( .A1(n_67), .A2(n_272), .B1(n_447), .B2(n_449), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_68), .B(n_646), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_69), .A2(n_213), .B1(n_357), .B2(n_574), .Y(n_808) );
CKINVDCx20_ASAP7_75t_R g788 ( .A(n_70), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_71), .B(n_427), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_72), .A2(n_159), .B1(n_540), .B2(n_680), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_75), .A2(n_185), .B1(n_414), .B2(n_415), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_77), .A2(n_154), .B1(n_340), .B2(n_577), .Y(n_576) );
AOI22xp33_ASAP7_75t_SL g691 ( .A1(n_78), .A2(n_145), .B1(n_390), .B2(n_435), .Y(n_691) );
AOI22xp33_ASAP7_75t_SL g715 ( .A1(n_79), .A2(n_121), .B1(n_716), .B2(n_717), .Y(n_715) );
AOI22xp33_ASAP7_75t_SL g537 ( .A1(n_80), .A2(n_111), .B1(n_417), .B2(n_538), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_82), .A2(n_139), .B1(n_335), .B2(n_574), .Y(n_573) );
AOI22xp33_ASAP7_75t_SL g698 ( .A1(n_84), .A2(n_222), .B1(n_330), .B2(n_477), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_85), .A2(n_211), .B1(n_415), .B2(n_550), .Y(n_597) );
INVx1_ASAP7_75t_L g294 ( .A(n_88), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_89), .B(n_844), .Y(n_843) );
CKINVDCx20_ASAP7_75t_R g348 ( .A(n_90), .Y(n_348) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_91), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_92), .B(n_465), .Y(n_464) );
AOI22xp33_ASAP7_75t_SL g702 ( .A1(n_93), .A2(n_187), .B1(n_323), .B2(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_94), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g292 ( .A(n_95), .Y(n_292) );
INVx1_ASAP7_75t_L g608 ( .A(n_96), .Y(n_608) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_99), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_100), .A2(n_207), .B1(n_359), .B2(n_477), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_101), .A2(n_141), .B1(n_477), .B2(n_577), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_102), .A2(n_243), .B1(n_335), .B2(n_547), .Y(n_802) );
CKINVDCx20_ASAP7_75t_R g838 ( .A(n_103), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_104), .A2(n_193), .B1(n_540), .B2(n_633), .Y(n_851) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_105), .Y(n_561) );
CKINVDCx20_ASAP7_75t_R g616 ( .A(n_106), .Y(n_616) );
CKINVDCx20_ASAP7_75t_R g556 ( .A(n_107), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_108), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_109), .A2(n_162), .B1(n_377), .B2(n_449), .Y(n_564) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_110), .Y(n_711) );
INVx1_ASAP7_75t_L g866 ( .A(n_113), .Y(n_866) );
OA22x2_ASAP7_75t_L g869 ( .A1(n_113), .A2(n_866), .B1(n_870), .B2(n_887), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_114), .A2(n_129), .B1(n_505), .B2(n_579), .Y(n_628) );
AOI22xp33_ASAP7_75t_SL g878 ( .A1(n_115), .A2(n_116), .B1(n_502), .B2(n_676), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_117), .A2(n_126), .B1(n_377), .B2(n_676), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_118), .B(n_424), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_119), .A2(n_225), .B1(n_359), .B2(n_545), .Y(n_763) );
OAI22xp5_ASAP7_75t_SL g739 ( .A1(n_120), .A2(n_740), .B1(n_741), .B2(n_764), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_120), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_123), .A2(n_258), .B1(n_356), .B2(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_124), .B(n_466), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_125), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_127), .A2(n_276), .B1(n_477), .B2(n_703), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g354 ( .A(n_128), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_131), .A2(n_203), .B1(n_335), .B2(n_574), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_132), .A2(n_167), .B1(n_419), .B2(n_420), .Y(n_418) );
AOI222xp33_ASAP7_75t_L g446 ( .A1(n_133), .A2(n_170), .B1(n_218), .B2(n_385), .C1(n_447), .C2(n_448), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_134), .A2(n_257), .B1(n_535), .B2(n_848), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_135), .A2(n_202), .B1(n_734), .B2(n_781), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_136), .A2(n_245), .B1(n_329), .B2(n_593), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_137), .A2(n_198), .B1(n_734), .B2(n_853), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_138), .A2(n_283), .B1(n_423), .B2(n_719), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_140), .A2(n_268), .B1(n_733), .B2(n_734), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g382 ( .A(n_142), .Y(n_382) );
INVx2_ASAP7_75t_L g295 ( .A(n_143), .Y(n_295) );
AOI22xp33_ASAP7_75t_SL g548 ( .A1(n_144), .A2(n_186), .B1(n_549), .B2(n_550), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_146), .Y(n_454) );
AOI22xp33_ASAP7_75t_SL g725 ( .A1(n_147), .A2(n_210), .B1(n_726), .B2(n_728), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_148), .Y(n_749) );
AOI222xp33_ASAP7_75t_L g791 ( .A1(n_149), .A2(n_163), .B1(n_227), .B2(n_385), .C1(n_607), .C2(n_792), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_150), .A2(n_254), .B1(n_390), .B2(n_840), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_151), .B(n_427), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_152), .A2(n_265), .B1(n_630), .B2(n_671), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_156), .A2(n_247), .B1(n_431), .B2(n_435), .Y(n_430) );
AOI22xp33_ASAP7_75t_SL g629 ( .A1(n_157), .A2(n_172), .B1(n_419), .B2(n_630), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g855 ( .A1(n_158), .A2(n_229), .B1(n_444), .B2(n_726), .Y(n_855) );
AND2x6_ASAP7_75t_L g291 ( .A(n_160), .B(n_292), .Y(n_291) );
HB1xp67_ASAP7_75t_L g822 ( .A(n_160), .Y(n_822) );
AO22x2_ASAP7_75t_L g309 ( .A1(n_161), .A2(n_236), .B1(n_310), .B2(n_311), .Y(n_309) );
AOI22xp33_ASAP7_75t_SL g526 ( .A1(n_164), .A2(n_205), .B1(n_466), .B2(n_527), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g327 ( .A(n_165), .Y(n_327) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_166), .Y(n_400) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_168), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_169), .A2(n_235), .B1(n_579), .B2(n_580), .Y(n_578) );
AOI22xp33_ASAP7_75t_SL g543 ( .A1(n_171), .A2(n_264), .B1(n_544), .B2(n_545), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_174), .B(n_424), .Y(n_674) );
XNOR2xp5_ASAP7_75t_L g705 ( .A(n_176), .B(n_706), .Y(n_705) );
AOI22xp33_ASAP7_75t_SL g722 ( .A1(n_177), .A2(n_178), .B1(n_538), .B2(n_723), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_179), .A2(n_275), .B1(n_439), .B2(n_441), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_180), .A2(n_612), .B1(n_613), .B2(n_635), .Y(n_611) );
CKINVDCx14_ASAP7_75t_R g635 ( .A(n_180), .Y(n_635) );
CKINVDCx20_ASAP7_75t_R g395 ( .A(n_181), .Y(n_395) );
AOI22xp33_ASAP7_75t_SL g886 ( .A1(n_182), .A2(n_269), .B1(n_352), .B2(n_580), .Y(n_886) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_183), .Y(n_682) );
AOI22xp33_ASAP7_75t_SL g885 ( .A1(n_188), .A2(n_259), .B1(n_477), .B2(n_577), .Y(n_885) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_189), .Y(n_461) );
AOI22xp33_ASAP7_75t_SL g699 ( .A1(n_190), .A2(n_232), .B1(n_481), .B2(n_652), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_191), .B(n_644), .Y(n_694) );
AO22x2_ASAP7_75t_L g314 ( .A1(n_192), .A2(n_248), .B1(n_310), .B2(n_315), .Y(n_314) );
AOI22xp33_ASAP7_75t_SL g650 ( .A1(n_195), .A2(n_253), .B1(n_439), .B2(n_580), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_196), .B(n_427), .Y(n_499) );
XOR2x2_ASAP7_75t_L g410 ( .A(n_197), .B(n_411), .Y(n_410) );
CKINVDCx20_ASAP7_75t_R g621 ( .A(n_200), .Y(n_621) );
AOI22xp33_ASAP7_75t_SL g651 ( .A1(n_201), .A2(n_206), .B1(n_574), .B2(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g568 ( .A(n_208), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_209), .Y(n_566) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_212), .Y(n_748) );
AOI22xp33_ASAP7_75t_SL g874 ( .A1(n_215), .A2(n_255), .B1(n_447), .B2(n_449), .Y(n_874) );
AOI22xp33_ASAP7_75t_SL g882 ( .A1(n_217), .A2(n_237), .B1(n_592), .B2(n_883), .Y(n_882) );
CKINVDCx20_ASAP7_75t_R g387 ( .A(n_219), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g370 ( .A(n_220), .Y(n_370) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_221), .A2(n_451), .B1(n_484), .B2(n_485), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_221), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g618 ( .A(n_223), .Y(n_618) );
AOI22xp33_ASAP7_75t_SL g695 ( .A1(n_226), .A2(n_279), .B1(n_433), .B2(n_447), .Y(n_695) );
AOI22xp33_ASAP7_75t_SL g511 ( .A1(n_228), .A2(n_274), .B1(n_361), .B2(n_512), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g624 ( .A(n_230), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_233), .A2(n_278), .B1(n_329), .B2(n_334), .Y(n_328) );
XOR2x2_ASAP7_75t_L g518 ( .A(n_234), .B(n_519), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_236), .B(n_827), .Y(n_826) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_242), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_244), .A2(n_251), .B1(n_443), .B2(n_444), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_246), .Y(n_772) );
INVx1_ASAP7_75t_L g825 ( .A(n_248), .Y(n_825) );
CKINVDCx20_ASAP7_75t_R g321 ( .A(n_249), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_250), .A2(n_280), .B1(n_423), .B2(n_427), .Y(n_422) );
INVx1_ASAP7_75t_L g525 ( .A(n_252), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g831 ( .A1(n_256), .A2(n_832), .B1(n_833), .B2(n_857), .Y(n_831) );
CKINVDCx20_ASAP7_75t_R g857 ( .A(n_256), .Y(n_857) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_260), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_263), .A2(n_266), .B1(n_342), .B2(n_577), .Y(n_634) );
INVx1_ASAP7_75t_L g704 ( .A(n_267), .Y(n_704) );
INVx1_ASAP7_75t_L g310 ( .A(n_271), .Y(n_310) );
INVx1_ASAP7_75t_L g312 ( .A(n_271), .Y(n_312) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_277), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g558 ( .A(n_282), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_284), .B(n_424), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g766 ( .A1(n_285), .A2(n_767), .B1(n_793), .B2(n_794), .Y(n_766) );
CKINVDCx16_ASAP7_75t_R g793 ( .A(n_285), .Y(n_793) );
CKINVDCx20_ASAP7_75t_R g287 ( .A(n_288), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_289), .Y(n_288) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
HB1xp67_ASAP7_75t_L g821 ( .A(n_292), .Y(n_821) );
OAI21xp5_ASAP7_75t_L g864 ( .A1(n_293), .A2(n_820), .B(n_865), .Y(n_864) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
AOI221xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_514), .B1(n_815), .B2(n_816), .C(n_817), .Y(n_296) );
INVx1_ASAP7_75t_L g816 ( .A(n_297), .Y(n_816) );
AOI22xp5_ASAP7_75t_SL g297 ( .A1(n_298), .A2(n_489), .B1(n_490), .B2(n_513), .Y(n_297) );
INVx1_ASAP7_75t_L g513 ( .A(n_298), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_300), .B1(n_409), .B2(n_488), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g408 ( .A(n_302), .Y(n_408) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_363), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g303 ( .A(n_304), .B(n_338), .Y(n_303) );
OAI221xp5_ASAP7_75t_SL g304 ( .A1(n_305), .A2(n_321), .B1(n_322), .B2(n_327), .C(n_328), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g773 ( .A(n_306), .Y(n_773) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_316), .Y(n_307) );
AND2x2_ASAP7_75t_L g332 ( .A(n_308), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g440 ( .A(n_308), .B(n_316), .Y(n_440) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_313), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_309), .B(n_314), .Y(n_326) );
INVx2_ASAP7_75t_L g346 ( .A(n_309), .Y(n_346) );
AND2x2_ASAP7_75t_L g381 ( .A(n_309), .B(n_318), .Y(n_381) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g315 ( .A(n_312), .Y(n_315) );
INVx1_ASAP7_75t_L g406 ( .A(n_313), .Y(n_406) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g347 ( .A(n_314), .Y(n_347) );
AND2x2_ASAP7_75t_L g353 ( .A(n_314), .B(n_346), .Y(n_353) );
INVx1_ASAP7_75t_L g380 ( .A(n_314), .Y(n_380) );
AND2x4_ASAP7_75t_L g324 ( .A(n_316), .B(n_325), .Y(n_324) );
AND2x4_ASAP7_75t_L g352 ( .A(n_316), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g358 ( .A(n_316), .B(n_345), .Y(n_358) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
AND2x2_ASAP7_75t_L g333 ( .A(n_317), .B(n_320), .Y(n_333) );
OR2x2_ASAP7_75t_L g344 ( .A(n_317), .B(n_320), .Y(n_344) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g386 ( .A(n_318), .B(n_320), .Y(n_386) );
AND2x2_ASAP7_75t_L g379 ( .A(n_319), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g399 ( .A(n_319), .Y(n_399) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g337 ( .A(n_320), .Y(n_337) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
BUFx3_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
BUFx3_ASAP7_75t_L g441 ( .A(n_324), .Y(n_441) );
BUFx2_ASAP7_75t_SL g510 ( .A(n_324), .Y(n_510) );
BUFx2_ASAP7_75t_SL g550 ( .A(n_324), .Y(n_550) );
BUFx2_ASAP7_75t_L g580 ( .A(n_324), .Y(n_580) );
BUFx3_ASAP7_75t_L g734 ( .A(n_324), .Y(n_734) );
INVx1_ASAP7_75t_L g805 ( .A(n_324), .Y(n_805) );
AND2x2_ASAP7_75t_L g652 ( .A(n_325), .B(n_399), .Y(n_652) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x6_ASAP7_75t_L g336 ( .A(n_326), .B(n_337), .Y(n_336) );
BUFx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_330), .Y(n_419) );
INVx5_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g574 ( .A(n_331), .Y(n_574) );
INVx4_ASAP7_75t_L g592 ( .A(n_331), .Y(n_592) );
INVx3_ASAP7_75t_L g671 ( .A(n_331), .Y(n_671) );
BUFx3_ASAP7_75t_L g727 ( .A(n_331), .Y(n_727) );
INVx8_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_L g362 ( .A(n_333), .B(n_345), .Y(n_362) );
NAND2x1p5_ASAP7_75t_L g373 ( .A(n_333), .B(n_353), .Y(n_373) );
AND2x6_ASAP7_75t_L g429 ( .A(n_333), .B(n_353), .Y(n_429) );
BUFx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx2_ASAP7_75t_L g420 ( .A(n_335), .Y(n_420) );
BUFx2_ASAP7_75t_L g593 ( .A(n_335), .Y(n_593) );
BUFx2_ASAP7_75t_L g630 ( .A(n_335), .Y(n_630) );
INVx6_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g728 ( .A(n_336), .Y(n_728) );
INVx1_ASAP7_75t_SL g883 ( .A(n_336), .Y(n_883) );
INVx1_ASAP7_75t_L g434 ( .A(n_337), .Y(n_434) );
OAI221xp5_ASAP7_75t_SL g338 ( .A1(n_339), .A2(n_348), .B1(n_349), .B2(n_354), .C(n_355), .Y(n_338) );
INVx1_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
INVx4_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g443 ( .A(n_341), .Y(n_443) );
INVx2_ASAP7_75t_SL g540 ( .A(n_341), .Y(n_540) );
INVx2_ASAP7_75t_L g596 ( .A(n_341), .Y(n_596) );
INVx5_ASAP7_75t_SL g783 ( .A(n_341), .Y(n_783) );
INVx11_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx11_ASAP7_75t_L g478 ( .A(n_342), .Y(n_478) );
AND2x6_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
AND2x4_ASAP7_75t_L g426 ( .A(n_343), .B(n_353), .Y(n_426) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g368 ( .A(n_344), .B(n_369), .Y(n_368) );
AND2x6_ASAP7_75t_L g385 ( .A(n_345), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx3_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_352), .Y(n_417) );
INVx2_ASAP7_75t_L g482 ( .A(n_352), .Y(n_482) );
BUFx3_ASAP7_75t_L g579 ( .A(n_352), .Y(n_579) );
BUFx3_ASAP7_75t_L g658 ( .A(n_352), .Y(n_658) );
INVx1_ASAP7_75t_L g369 ( .A(n_353), .Y(n_369) );
BUFx3_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_357), .Y(n_544) );
INVx3_ASAP7_75t_L g724 ( .A(n_357), .Y(n_724) );
BUFx3_ASAP7_75t_L g762 ( .A(n_357), .Y(n_762) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
BUFx2_ASAP7_75t_SL g414 ( .A(n_358), .Y(n_414) );
BUFx2_ASAP7_75t_SL g505 ( .A(n_358), .Y(n_505) );
INVx2_ASAP7_75t_L g657 ( .A(n_358), .Y(n_657) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx3_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx3_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx6_ASAP7_75t_L g445 ( .A(n_362), .Y(n_445) );
BUFx3_ASAP7_75t_L g680 ( .A(n_362), .Y(n_680) );
BUFx3_ASAP7_75t_L g703 ( .A(n_362), .Y(n_703) );
NOR3xp33_ASAP7_75t_L g363 ( .A(n_364), .B(n_374), .C(n_394), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_366), .B1(n_370), .B2(n_371), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g453 ( .A1(n_366), .A2(n_454), .B1(n_455), .B2(n_456), .Y(n_453) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g617 ( .A(n_367), .Y(n_617) );
INVx1_ASAP7_75t_SL g745 ( .A(n_367), .Y(n_745) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx3_ASAP7_75t_L g557 ( .A(n_368), .Y(n_557) );
BUFx6f_ASAP7_75t_L g787 ( .A(n_368), .Y(n_787) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g559 ( .A(n_372), .Y(n_559) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx3_ASAP7_75t_L g458 ( .A(n_373), .Y(n_458) );
OAI222xp33_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_382), .B1(n_383), .B2(n_387), .C1(n_388), .C2(n_393), .Y(n_374) );
OAI221xp5_ASAP7_75t_SL g747 ( .A1(n_375), .A2(n_522), .B1(n_748), .B2(n_749), .C(n_750), .Y(n_747) );
INVx2_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx4f_ASAP7_75t_SL g447 ( .A(n_378), .Y(n_447) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_378), .Y(n_529) );
BUFx2_ASAP7_75t_L g607 ( .A(n_378), .Y(n_607) );
BUFx6f_ASAP7_75t_L g848 ( .A(n_378), .Y(n_848) );
AND2x4_ASAP7_75t_L g378 ( .A(n_379), .B(n_381), .Y(n_378) );
INVx1_ASAP7_75t_L g392 ( .A(n_380), .Y(n_392) );
AND2x4_ASAP7_75t_L g391 ( .A(n_381), .B(n_392), .Y(n_391) );
NAND2x1p5_ASAP7_75t_L g398 ( .A(n_381), .B(n_399), .Y(n_398) );
AND2x4_ASAP7_75t_L g433 ( .A(n_381), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_SL g460 ( .A(n_384), .Y(n_460) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx4_ASAP7_75t_L g524 ( .A(n_385), .Y(n_524) );
BUFx3_ASAP7_75t_L g563 ( .A(n_385), .Y(n_563) );
INVx2_ASAP7_75t_L g689 ( .A(n_385), .Y(n_689) );
INVx2_ASAP7_75t_SL g837 ( .A(n_385), .Y(n_837) );
INVx1_ASAP7_75t_L g404 ( .A(n_386), .Y(n_404) );
AND2x4_ASAP7_75t_L g436 ( .A(n_386), .B(n_406), .Y(n_436) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx2_ASAP7_75t_L g792 ( .A(n_390), .Y(n_792) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
BUFx12f_ASAP7_75t_L g449 ( .A(n_391), .Y(n_449) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_391), .Y(n_466) );
INVx1_ASAP7_75t_L g712 ( .A(n_391), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B1(n_400), .B2(n_401), .Y(n_394) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx4_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_398), .Y(n_469) );
BUFx3_ASAP7_75t_L g567 ( .A(n_398), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_401), .A2(n_468), .B1(n_469), .B2(n_470), .Y(n_467) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g754 ( .A(n_402), .Y(n_754) );
CKINVDCx16_ASAP7_75t_R g402 ( .A(n_403), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_403), .A2(n_566), .B1(n_567), .B2(n_568), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_403), .A2(n_469), .B1(n_624), .B2(n_625), .Y(n_623) );
OR2x6_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx3_ASAP7_75t_L g488 ( .A(n_409), .Y(n_488) );
OA22x2_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_450), .B1(n_486), .B2(n_487), .Y(n_409) );
INVx1_ASAP7_75t_L g487 ( .A(n_410), .Y(n_487) );
NAND4xp75_ASAP7_75t_L g411 ( .A(n_412), .B(n_421), .C(n_437), .D(n_446), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_418), .Y(n_412) );
INVx4_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx3_ASAP7_75t_L g733 ( .A(n_416), .Y(n_733) );
INVx4_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_SL g421 ( .A(n_422), .B(n_430), .Y(n_421) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_424), .Y(n_844) );
INVx5_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g533 ( .A(n_425), .Y(n_533) );
INVx2_ASAP7_75t_L g600 ( .A(n_425), .Y(n_600) );
INVx2_ASAP7_75t_L g646 ( .A(n_425), .Y(n_646) );
INVx4_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_SL g719 ( .A(n_428), .Y(n_719) );
INVx1_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
BUFx4f_ASAP7_75t_L g644 ( .A(n_429), .Y(n_644) );
BUFx2_ASAP7_75t_L g846 ( .A(n_429), .Y(n_846) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx2_ASAP7_75t_L g535 ( .A(n_433), .Y(n_535) );
BUFx3_ASAP7_75t_L g676 ( .A(n_433), .Y(n_676) );
BUFx2_ASAP7_75t_L g716 ( .A(n_433), .Y(n_716) );
BUFx2_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
BUFx2_ASAP7_75t_SL g502 ( .A(n_436), .Y(n_502) );
BUFx6f_ASAP7_75t_L g602 ( .A(n_436), .Y(n_602) );
BUFx3_ASAP7_75t_L g717 ( .A(n_436), .Y(n_717) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_442), .Y(n_437) );
INVx1_ASAP7_75t_L g475 ( .A(n_439), .Y(n_475) );
BUFx2_ASAP7_75t_L g731 ( .A(n_439), .Y(n_731) );
BUFx3_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx3_ASAP7_75t_L g509 ( .A(n_440), .Y(n_509) );
BUFx3_ASAP7_75t_L g547 ( .A(n_440), .Y(n_547) );
BUFx3_ASAP7_75t_L g572 ( .A(n_440), .Y(n_572) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g549 ( .A(n_445), .Y(n_549) );
INVx3_ASAP7_75t_L g577 ( .A(n_445), .Y(n_577) );
INVx1_ASAP7_75t_L g462 ( .A(n_447), .Y(n_462) );
BUFx4f_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g497 ( .A(n_449), .Y(n_497) );
INVx1_ASAP7_75t_L g486 ( .A(n_450), .Y(n_486) );
INVx2_ASAP7_75t_L g485 ( .A(n_451), .Y(n_485) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_471), .Y(n_451) );
NOR3xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_459), .C(n_467), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_456), .A2(n_744), .B1(n_745), .B2(n_746), .Y(n_743) );
OAI221xp5_ASAP7_75t_SL g786 ( .A1(n_456), .A2(n_787), .B1(n_788), .B2(n_789), .C(n_790), .Y(n_786) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx3_ASAP7_75t_L g619 ( .A(n_458), .Y(n_619) );
OAI221xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B1(n_462), .B2(n_463), .C(n_464), .Y(n_459) );
OAI21xp5_ASAP7_75t_SL g493 ( .A1(n_460), .A2(n_494), .B(n_495), .Y(n_493) );
OAI222xp33_ASAP7_75t_L g708 ( .A1(n_460), .A2(n_709), .B1(n_710), .B2(n_711), .C1(n_712), .C2(n_713), .Y(n_708) );
BUFx4f_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_479), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_476), .Y(n_472) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx4_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_SL g512 ( .A(n_478), .Y(n_512) );
INVx3_ASAP7_75t_L g758 ( .A(n_478), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_483), .Y(n_479) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NAND3xp33_ASAP7_75t_L g491 ( .A(n_492), .B(n_503), .C(n_507), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_498), .Y(n_492) );
INVx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
NAND3xp33_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .C(n_501), .Y(n_498) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_506), .Y(n_503) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_511), .Y(n_507) );
BUFx4f_ASAP7_75t_SL g633 ( .A(n_509), .Y(n_633) );
INVx1_ASAP7_75t_L g815 ( .A(n_514), .Y(n_815) );
XNOR2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_583), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_551), .B1(n_552), .B2(n_582), .Y(n_517) );
INVx2_ASAP7_75t_L g582 ( .A(n_518), .Y(n_582) );
NAND3x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_536), .C(n_542), .Y(n_519) );
NOR2x1_ASAP7_75t_SL g520 ( .A(n_521), .B(n_530), .Y(n_520) );
OAI21xp5_ASAP7_75t_SL g521 ( .A1(n_522), .A2(n_525), .B(n_526), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx4_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx2_ASAP7_75t_L g604 ( .A(n_524), .Y(n_604) );
INVx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx4_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g710 ( .A(n_529), .Y(n_710) );
NAND3xp33_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .C(n_534), .Y(n_530) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_541), .Y(n_536) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_548), .Y(n_542) );
INVx1_ASAP7_75t_SL g776 ( .A(n_544), .Y(n_776) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g771 ( .A(n_549), .Y(n_771) );
INVx2_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
XOR2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_581), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_569), .Y(n_553) );
NOR3xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_560), .C(n_565), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B1(n_558), .B2(n_559), .Y(n_555) );
OAI21xp33_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_562), .B(n_564), .Y(n_560) );
OAI21xp5_ASAP7_75t_SL g639 ( .A1(n_562), .A2(n_640), .B(n_641), .Y(n_639) );
OAI21xp5_ASAP7_75t_SL g872 ( .A1(n_562), .A2(n_873), .B(n_874), .Y(n_872) );
INVx3_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_567), .A2(n_752), .B1(n_753), .B2(n_754), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_575), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_578), .Y(n_575) );
INVxp67_ASAP7_75t_L g778 ( .A(n_579), .Y(n_778) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_585), .B1(n_663), .B2(n_814), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_609), .B1(n_610), .B2(n_662), .Y(n_585) );
INVx2_ASAP7_75t_SL g662 ( .A(n_586), .Y(n_662) );
XOR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_608), .Y(n_586) );
NOR4xp75_ASAP7_75t_L g587 ( .A(n_588), .B(n_594), .C(n_598), .D(n_603), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_589), .B(n_590), .Y(n_588) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND2x1_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_599), .B(n_601), .Y(n_598) );
INVx1_ASAP7_75t_SL g841 ( .A(n_602), .Y(n_841) );
OAI21xp5_ASAP7_75t_SL g603 ( .A1(n_604), .A2(n_605), .B(n_606), .Y(n_603) );
OAI21xp5_ASAP7_75t_SL g620 ( .A1(n_604), .A2(n_621), .B(n_622), .Y(n_620) );
INVx2_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
AO22x1_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_636), .B1(n_660), .B2(n_661), .Y(n_610) );
INVx1_ASAP7_75t_L g661 ( .A(n_611), .Y(n_661) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_626), .Y(n_613) );
NOR3xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_620), .C(n_623), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_617), .B1(n_618), .B2(n_619), .Y(n_615) );
OA211x2_ASAP7_75t_L g672 ( .A1(n_619), .A2(n_673), .B(n_674), .C(n_675), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_627), .B(n_631), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_634), .Y(n_631) );
INVx3_ASAP7_75t_SL g660 ( .A(n_636), .Y(n_660) );
XOR2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_659), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_638), .B(n_648), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_639), .B(n_642), .Y(n_638) );
NAND3xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .C(n_647), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_649), .B(n_653), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
INVx3_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx3_ASAP7_75t_L g853 ( .A(n_657), .Y(n_853) );
INVx1_ASAP7_75t_L g814 ( .A(n_663), .Y(n_814) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_737), .B1(n_812), .B2(n_813), .Y(n_663) );
INVx1_ASAP7_75t_L g812 ( .A(n_664), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_666), .B1(n_683), .B2(n_736), .Y(n_664) );
INVx3_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
XOR2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_682), .Y(n_666) );
NAND4xp75_ASAP7_75t_L g667 ( .A(n_668), .B(n_672), .C(n_677), .D(n_681), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
AND2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
INVx2_ASAP7_75t_L g736 ( .A(n_683), .Y(n_736) );
OA22x2_ASAP7_75t_SL g683 ( .A1(n_684), .A2(n_685), .B1(n_705), .B2(n_735), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
XOR2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_704), .Y(n_685) );
NAND2x1_ASAP7_75t_L g686 ( .A(n_687), .B(n_696), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_688), .B(n_692), .Y(n_687) );
OAI21xp5_ASAP7_75t_SL g688 ( .A1(n_689), .A2(n_690), .B(n_691), .Y(n_688) );
NAND3xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .C(n_695), .Y(n_692) );
NOR2x1_ASAP7_75t_L g696 ( .A(n_697), .B(n_700), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
INVx1_ASAP7_75t_L g735 ( .A(n_705), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_707), .B(n_720), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_714), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_715), .B(n_718), .Y(n_714) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_729), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_725), .Y(n_721) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx3_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_732), .Y(n_729) );
INVx1_ASAP7_75t_L g813 ( .A(n_737), .Y(n_813) );
XNOR2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_765), .Y(n_737) );
BUFx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_742), .B(n_755), .Y(n_741) );
NOR3xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_747), .C(n_751), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_756), .B(n_760), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_757), .B(n_759), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_763), .Y(n_760) );
AOI22xp5_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_795), .B1(n_810), .B2(n_811), .Y(n_765) );
INVx1_ASAP7_75t_L g810 ( .A(n_766), .Y(n_810) );
INVx2_ASAP7_75t_SL g794 ( .A(n_767), .Y(n_794) );
AND4x1_ASAP7_75t_L g767 ( .A(n_768), .B(n_779), .C(n_785), .D(n_791), .Y(n_767) );
NOR2xp33_ASAP7_75t_L g768 ( .A(n_769), .B(n_774), .Y(n_768) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_771), .B1(n_772), .B2(n_773), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_776), .B1(n_777), .B2(n_778), .Y(n_774) );
AND2x2_ASAP7_75t_L g779 ( .A(n_780), .B(n_784), .Y(n_779) );
INVx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVxp67_ASAP7_75t_L g811 ( .A(n_795), .Y(n_811) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
NAND4xp75_ASAP7_75t_L g797 ( .A(n_798), .B(n_801), .C(n_806), .D(n_809), .Y(n_797) );
AND2x2_ASAP7_75t_SL g798 ( .A(n_799), .B(n_800), .Y(n_798) );
AND2x2_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .Y(n_801) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
AND2x2_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
INVx1_ASAP7_75t_SL g817 ( .A(n_818), .Y(n_817) );
NOR2x1_ASAP7_75t_L g818 ( .A(n_819), .B(n_823), .Y(n_818) );
OR2x2_ASAP7_75t_SL g888 ( .A(n_819), .B(n_824), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_820), .B(n_822), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g859 ( .A(n_820), .Y(n_859) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_821), .B(n_862), .Y(n_865) );
CKINVDCx16_ASAP7_75t_R g862 ( .A(n_822), .Y(n_862) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_824), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_825), .B(n_826), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_828), .B(n_829), .Y(n_827) );
OAI322xp33_ASAP7_75t_L g830 ( .A1(n_831), .A2(n_858), .A3(n_860), .B1(n_863), .B2(n_866), .C1(n_867), .C2(n_888), .Y(n_830) );
CKINVDCx20_ASAP7_75t_R g832 ( .A(n_833), .Y(n_832) );
HB1xp67_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
NAND2xp5_ASAP7_75t_SL g834 ( .A(n_835), .B(n_849), .Y(n_834) );
NOR2xp33_ASAP7_75t_SL g835 ( .A(n_836), .B(n_842), .Y(n_835) );
OAI21xp5_ASAP7_75t_SL g836 ( .A1(n_837), .A2(n_838), .B(n_839), .Y(n_836) );
INVx2_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
NAND3xp33_ASAP7_75t_L g842 ( .A(n_843), .B(n_845), .C(n_847), .Y(n_842) );
NOR2x1_ASAP7_75t_L g849 ( .A(n_850), .B(n_854), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_851), .B(n_852), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_855), .B(n_856), .Y(n_854) );
BUFx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
HB1xp67_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
CKINVDCx20_ASAP7_75t_R g863 ( .A(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g887 ( .A(n_870), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_871), .B(n_879), .Y(n_870) );
NOR2xp67_ASAP7_75t_L g871 ( .A(n_872), .B(n_875), .Y(n_871) );
NAND3xp33_ASAP7_75t_L g875 ( .A(n_876), .B(n_877), .C(n_878), .Y(n_875) );
NOR2x1_ASAP7_75t_L g879 ( .A(n_880), .B(n_884), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_881), .B(n_882), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_885), .B(n_886), .Y(n_884) );
endmodule