module fake_jpeg_20257_n_319 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_319);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_145;
wire n_18;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_28),
.Y(n_39)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_31),
.Y(n_38)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_32),
.B(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_13),
.Y(n_59)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_32),
.Y(n_41)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_30),
.A2(n_14),
.B1(n_13),
.B2(n_17),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_47),
.Y(n_62)
);

INVxp33_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_56),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_49),
.Y(n_68)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_29),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_25),
.Y(n_73)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_59),
.B(n_36),
.Y(n_77)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_61),
.Y(n_79)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_53),
.A2(n_41),
.B(n_39),
.C(n_38),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_35),
.B1(n_40),
.B2(n_45),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_53),
.A2(n_43),
.B1(n_41),
.B2(n_39),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_52),
.B1(n_35),
.B2(n_55),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_SL g69 ( 
.A(n_54),
.B(n_36),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_69),
.B(n_52),
.Y(n_82)
);

AOI32xp33_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_38),
.A3(n_37),
.B1(n_28),
.B2(n_26),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_73),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_47),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_77),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_80),
.A2(n_93),
.B1(n_95),
.B2(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_15),
.Y(n_121)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_66),
.Y(n_122)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

NOR2x1_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_65),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_87),
.A2(n_88),
.B(n_82),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_65),
.A2(n_52),
.B(n_15),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_71),
.B1(n_67),
.B2(n_73),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_64),
.B(n_19),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_35),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_97),
.Y(n_102)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_91),
.B(n_78),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_92),
.A2(n_68),
.B(n_75),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_63),
.A2(n_40),
.B1(n_45),
.B2(n_58),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_63),
.A2(n_45),
.B1(n_51),
.B2(n_55),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_68),
.A2(n_45),
.B1(n_27),
.B2(n_49),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_44),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_97),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_101),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_86),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_91),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_106),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_116),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_83),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_64),
.C(n_75),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_25),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_60),
.B1(n_68),
.B2(n_49),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_109),
.A2(n_57),
.B1(n_72),
.B2(n_56),
.Y(n_146)
);

BUFx12_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_112),
.A2(n_113),
.B(n_101),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_115),
.A2(n_118),
.B(n_120),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_81),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_89),
.A2(n_80),
.B1(n_92),
.B2(n_88),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_87),
.B1(n_94),
.B2(n_90),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_11),
.B(n_21),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_85),
.A2(n_72),
.B1(n_46),
.B2(n_62),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_119),
.A2(n_124),
.B1(n_66),
.B2(n_62),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_87),
.A2(n_21),
.B(n_19),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_93),
.Y(n_141)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_62),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_123),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_84),
.A2(n_72),
.B1(n_62),
.B2(n_50),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_126),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_103),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_131),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_92),
.Y(n_128)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_116),
.B(n_98),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_103),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_134),
.B(n_136),
.Y(n_185)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_138),
.A2(n_157),
.B1(n_110),
.B2(n_31),
.Y(n_177)
);

AOI22x1_ASAP7_75t_SL g140 ( 
.A1(n_113),
.A2(n_88),
.B1(n_94),
.B2(n_98),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_140),
.A2(n_144),
.B1(n_153),
.B2(n_110),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_141),
.B(n_23),
.Y(n_184)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_95),
.B(n_93),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_143),
.A2(n_156),
.B(n_112),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_95),
.B1(n_98),
.B2(n_96),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_108),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_149),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_154),
.B1(n_155),
.B2(n_111),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_42),
.Y(n_147)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_29),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_152),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_114),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_151),
.B(n_114),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_106),
.A2(n_14),
.B1(n_18),
.B2(n_15),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_100),
.A2(n_61),
.B1(n_42),
.B2(n_14),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_102),
.A2(n_34),
.B1(n_33),
.B2(n_24),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_111),
.A2(n_34),
.B1(n_33),
.B2(n_24),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_158),
.A2(n_128),
.B(n_137),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_104),
.Y(n_161)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_161),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_162),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_133),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_164),
.B(n_166),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_130),
.Y(n_166)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_169),
.A2(n_174),
.B1(n_157),
.B2(n_129),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_139),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_171),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_132),
.B(n_121),
.Y(n_171)
);

AOI21x1_ASAP7_75t_SL g172 ( 
.A1(n_125),
.A2(n_120),
.B(n_113),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_172),
.A2(n_143),
.B(n_148),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_173),
.A2(n_177),
.B1(n_182),
.B2(n_155),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_149),
.A2(n_110),
.B1(n_78),
.B2(n_70),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_152),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_178),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_78),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_183),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_142),
.A2(n_18),
.B1(n_20),
.B2(n_16),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_154),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_147),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_141),
.B(n_23),
.C(n_20),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_146),
.C(n_135),
.Y(n_202)
);

INVx13_ASAP7_75t_L g188 ( 
.A(n_185),
.Y(n_188)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_176),
.B(n_125),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_184),
.Y(n_215)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_194),
.A2(n_6),
.B(n_10),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_195),
.B(n_22),
.Y(n_233)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_186),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_196),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_129),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_199),
.Y(n_231)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_206),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_201),
.A2(n_204),
.B(n_147),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_202),
.B(n_0),
.C(n_1),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_128),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_163),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_205),
.B(n_207),
.Y(n_218)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_168),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_178),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_158),
.B(n_127),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_211),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_136),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_179),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_6),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_213),
.A2(n_180),
.B1(n_183),
.B2(n_169),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_175),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_225),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_223),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_216),
.A2(n_234),
.B1(n_204),
.B2(n_196),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_190),
.A2(n_180),
.B1(n_160),
.B2(n_174),
.Y(n_217)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_202),
.A2(n_187),
.B1(n_172),
.B2(n_162),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_222),
.A2(n_226),
.B1(n_209),
.B2(n_193),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_176),
.Y(n_225)
);

AOI21xp33_ASAP7_75t_L g226 ( 
.A1(n_203),
.A2(n_177),
.B(n_7),
.Y(n_226)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_227),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_6),
.Y(n_228)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_228),
.Y(n_255)
);

FAx1_ASAP7_75t_SL g229 ( 
.A(n_191),
.B(n_20),
.CI(n_22),
.CON(n_229),
.SN(n_229)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_234),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_232),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_194),
.B(n_22),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_195),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_210),
.A2(n_20),
.B1(n_1),
.B2(n_2),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_233),
.C(n_200),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_235),
.Y(n_238)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_238),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_240),
.A2(n_223),
.B1(n_206),
.B2(n_204),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_222),
.A2(n_210),
.B1(n_209),
.B2(n_213),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_241),
.A2(n_253),
.B1(n_189),
.B2(n_229),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_246),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_201),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_220),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_250),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_231),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_214),
.B(n_232),
.C(n_221),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_240),
.C(n_246),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_224),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_252),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_219),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_211),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_192),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_218),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_261),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_260),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_263),
.B(n_269),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_237),
.B(n_215),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_270),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_192),
.C(n_229),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_268),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_248),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_230),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_241),
.A2(n_10),
.B1(n_9),
.B2(n_8),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_9),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_259),
.B(n_243),
.Y(n_273)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_237),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_276),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_262),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_239),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_278),
.B(n_283),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_265),
.A2(n_264),
.B1(n_257),
.B2(n_261),
.Y(n_279)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_279),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_280),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_282),
.A2(n_6),
.B1(n_8),
.B2(n_7),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_242),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_242),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_284),
.B(n_9),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_272),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_297),
.Y(n_299)
);

INVx11_ASAP7_75t_L g287 ( 
.A(n_280),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_288),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_255),
.C(n_1),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_0),
.C(n_1),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_293),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_0),
.C(n_1),
.Y(n_293)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_294),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_293),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_282),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_291),
.A2(n_281),
.B1(n_3),
.B2(n_4),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_305),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_303),
.Y(n_308)
);

AOI21x1_ASAP7_75t_L g304 ( 
.A1(n_285),
.A2(n_281),
.B(n_3),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_304),
.A2(n_297),
.B(n_4),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_2),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_2),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_292),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_310),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_298),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_298),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_308),
.C(n_288),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_289),
.Y(n_315)
);

MAJx2_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_287),
.C(n_299),
.Y(n_316)
);

A2O1A1Ixp33_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_313),
.B(n_307),
.C(n_301),
.Y(n_317)
);

OAI21x1_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_295),
.B(n_4),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_3),
.B(n_5),
.Y(n_319)
);


endmodule