module fake_jpeg_18674_n_168 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_168);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_20),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_33),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_32),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_22),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_3),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_26),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_12),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_10),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_0),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_9),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_48),
.Y(n_74)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_2),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_3),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_11),
.Y(n_77)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_49),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_84),
.Y(n_93)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_86),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_81),
.A2(n_50),
.B1(n_75),
.B2(n_65),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_95),
.B1(n_60),
.B2(n_76),
.Y(n_108)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_84),
.A2(n_68),
.B1(n_53),
.B2(n_52),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_79),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_82),
.A2(n_54),
.B1(n_58),
.B2(n_59),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_89),
.A2(n_86),
.B1(n_83),
.B2(n_79),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_56),
.B1(n_73),
.B2(n_62),
.Y(n_117)
);

OR2x2_ASAP7_75t_SL g100 ( 
.A(n_95),
.B(n_71),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_100),
.A2(n_56),
.B(n_74),
.Y(n_115)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_105),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_71),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_72),
.Y(n_113)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_107),
.Y(n_126)
);

OAI22x1_ASAP7_75t_L g123 ( 
.A1(n_108),
.A2(n_64),
.B1(n_57),
.B2(n_77),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_63),
.B1(n_61),
.B2(n_64),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_106),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_113),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_108),
.A2(n_88),
.B1(n_97),
.B2(n_67),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_117),
.B1(n_118),
.B2(n_125),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_98),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_120),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_123),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_99),
.A2(n_77),
.B1(n_69),
.B2(n_66),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_70),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_124),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_123),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_69),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_66),
.B1(n_21),
.B2(n_23),
.Y(n_125)
);

AOI21xp33_ASAP7_75t_L g127 ( 
.A1(n_100),
.A2(n_18),
.B(n_45),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_127),
.A2(n_119),
.B1(n_8),
.B2(n_9),
.Y(n_142)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_117),
.B(n_0),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_133),
.A2(n_138),
.B(n_7),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_1),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_136),
.Y(n_144)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_139),
.A2(n_141),
.B1(n_127),
.B2(n_112),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_142),
.B(n_24),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_146),
.Y(n_153)
);

OAI32xp33_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_29),
.A3(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_148)
);

XOR2x2_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_141),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_138),
.A2(n_8),
.B(n_17),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_151),
.C(n_137),
.Y(n_155)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_152),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_153),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_157),
.B(n_144),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_155),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_154),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

BUFx24_ASAP7_75t_SL g162 ( 
.A(n_161),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_140),
.B(n_145),
.Y(n_163)
);

A2O1A1O1Ixp25_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_154),
.B(n_150),
.C(n_129),
.D(n_143),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_164),
.Y(n_165)
);

AOI21xp33_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_25),
.B(n_30),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_166),
.A2(n_36),
.B(n_40),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_41),
.B(n_42),
.Y(n_168)
);


endmodule