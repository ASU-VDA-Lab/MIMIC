module fake_jpeg_2002_n_229 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_229);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_25),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_33),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_21),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_23),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_25),
.Y(n_72)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

BUFx16f_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

BUFx6f_ASAP7_75t_SL g77 ( 
.A(n_45),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_12),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_11),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_3),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_86),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_88),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_89),
.B(n_55),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_82),
.A2(n_65),
.B1(n_58),
.B2(n_72),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_102),
.B1(n_58),
.B2(n_77),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_101),
.Y(n_107)
);

NAND3xp33_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_69),
.C(n_64),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_64),
.B1(n_79),
.B2(n_55),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_79),
.B1(n_63),
.B2(n_74),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_89),
.A2(n_77),
.B1(n_72),
.B2(n_80),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_62),
.B1(n_71),
.B2(n_60),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_86),
.B(n_68),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_82),
.A2(n_58),
.B1(n_69),
.B2(n_80),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_76),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_63),
.Y(n_113)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_76),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_106),
.B(n_108),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_61),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_SL g126 ( 
.A1(n_109),
.A2(n_113),
.B(n_67),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_110),
.A2(n_111),
.B1(n_122),
.B2(n_78),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_93),
.B1(n_91),
.B2(n_98),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_92),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_112),
.Y(n_129)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_119),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_118),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_60),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_70),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_0),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_62),
.B1(n_75),
.B2(n_57),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_121),
.A2(n_85),
.B1(n_59),
.B2(n_54),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_96),
.A2(n_78),
.B1(n_70),
.B2(n_67),
.Y(n_122)
);

INVxp67_ASAP7_75t_SL g123 ( 
.A(n_100),
.Y(n_123)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

OAI22x1_ASAP7_75t_L g125 ( 
.A1(n_111),
.A2(n_100),
.B1(n_85),
.B2(n_59),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_125),
.A2(n_141),
.B1(n_128),
.B2(n_142),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_127),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_128),
.A2(n_132),
.B1(n_144),
.B2(n_130),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_54),
.B1(n_66),
.B2(n_2),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_66),
.B(n_1),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_133),
.A2(n_121),
.B(n_114),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_138),
.B(n_139),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_116),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_53),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_133),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_110),
.A2(n_66),
.B1(n_1),
.B2(n_2),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_115),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_143),
.B(n_5),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_104),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_145),
.B(n_13),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_105),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_153),
.C(n_157),
.Y(n_171)
);

NAND3xp33_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_156),
.C(n_169),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_152),
.A2(n_165),
.B1(n_167),
.B2(n_17),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_52),
.C(n_51),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_4),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_154),
.B(n_162),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_160),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_6),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_50),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_49),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_15),
.C(n_17),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_6),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_144),
.A2(n_7),
.B(n_9),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_163),
.A2(n_18),
.B(n_19),
.Y(n_185)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_170),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_131),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_166),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_14),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_26),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_179),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_168),
.A2(n_15),
.B(n_16),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_177),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_180),
.A2(n_181),
.B1(n_42),
.B2(n_47),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_168),
.A2(n_152),
.B1(n_146),
.B2(n_165),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_161),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_182),
.A2(n_189),
.B1(n_39),
.B2(n_40),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_150),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_186),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_166),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_20),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_188),
.Y(n_194)
);

OAI32xp33_ASAP7_75t_L g193 ( 
.A1(n_191),
.A2(n_24),
.A3(n_27),
.B1(n_29),
.B2(n_36),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_193),
.A2(n_202),
.B1(n_189),
.B2(n_186),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_37),
.C(n_38),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_203),
.C(n_179),
.Y(n_205)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_190),
.Y(n_197)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_197),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_199),
.B(n_201),
.Y(n_206)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_176),
.C(n_191),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_178),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_195),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_205),
.B(n_211),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_181),
.Y(n_207)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_210),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_202),
.A2(n_177),
.B1(n_173),
.B2(n_187),
.Y(n_210)
);

BUFx24_ASAP7_75t_SL g211 ( 
.A(n_194),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_196),
.A2(n_172),
.B(n_174),
.Y(n_212)
);

AO21x1_ASAP7_75t_L g215 ( 
.A1(n_212),
.A2(n_192),
.B(n_185),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_207),
.A2(n_192),
.B1(n_196),
.B2(n_174),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_213),
.A2(n_209),
.B1(n_206),
.B2(n_193),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_205),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_215),
.Y(n_220)
);

NOR3xp33_ASAP7_75t_SL g223 ( 
.A(n_219),
.B(n_217),
.C(n_214),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_221),
.A2(n_218),
.B1(n_216),
.B2(n_213),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_223),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_220),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_215),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_219),
.C(n_198),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_227),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_184),
.Y(n_229)
);


endmodule