module real_jpeg_5457_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_173;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_1),
.B(n_45),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_1),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_2),
.B(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_2),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_2),
.B(n_101),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_3),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_4),
.B(n_34),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_4),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_4),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_4),
.B(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_4),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_5),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_5),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_5),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_5),
.B(n_148),
.Y(n_147)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_7),
.Y(n_93)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_7),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_7),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_8),
.Y(n_112)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_9),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_10),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_10),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_10),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_10),
.B(n_126),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_10),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_11),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_11),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_11),
.B(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_11),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_11),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_11),
.B(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_12),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_13),
.B(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_120),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_119),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_81),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_18),
.B(n_81),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_49),
.C(n_62),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_19),
.A2(n_20),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_30),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_21),
.B(n_31),
.C(n_37),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_27),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_22),
.B(n_27),
.Y(n_163)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_37),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_36),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_43),
.B1(n_44),
.B2(n_48),
.Y(n_37)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_42),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_43),
.B(n_48),
.Y(n_117)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_49),
.A2(n_62),
.B1(n_63),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_49),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_54),
.C(n_56),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_50),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_166)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_56),
.B(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_60),
.Y(n_140)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_69),
.Y(n_63)
);

MAJx2_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_70),
.C(n_80),
.Y(n_95)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_75),
.B2(n_80),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_106),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_96),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_94),
.B2(n_95),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_93),
.Y(n_157)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx24_ASAP7_75t_SL g178 ( 
.A(n_96),
.Y(n_178)
);

FAx1_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_100),
.CI(n_103),
.CON(n_96),
.SN(n_96)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_118),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_117),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OA21x2_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_169),
.B(n_176),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_160),
.B(n_168),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_149),
.B(n_159),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_131),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_131),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_128),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_141),
.B2(n_142),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_136),
.C(n_141),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_147),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_147),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_154),
.B(n_158),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_152),
.Y(n_158)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_167),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_167),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_164),
.C(n_171),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_165),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_172),
.Y(n_176)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);


endmodule