module fake_jpeg_7309_n_176 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_6),
.B(n_14),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_15),
.B(n_0),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_17),
.C(n_28),
.Y(n_45)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_40),
.Y(n_48)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_30),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_44),
.B(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_30),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_17),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_41),
.B(n_40),
.C(n_38),
.Y(n_63)
);

CKINVDCx6p67_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_18),
.B1(n_28),
.B2(n_31),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_55),
.A2(n_57),
.B1(n_18),
.B2(n_22),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_33),
.A2(n_15),
.B1(n_22),
.B2(n_31),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_40),
.B(n_25),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_23),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_64),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_75),
.B1(n_78),
.B2(n_41),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_74),
.Y(n_88)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_23),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_66),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_20),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_20),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_27),
.Y(n_70)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_71),
.Y(n_92)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_46),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_52),
.Y(n_83)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_79),
.B(n_27),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_73),
.Y(n_104)
);

AOI22x1_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_62),
.B1(n_36),
.B2(n_56),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_95),
.B1(n_98),
.B2(n_47),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_83),
.B(n_84),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_52),
.B1(n_33),
.B2(n_42),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_86),
.A2(n_72),
.B1(n_68),
.B2(n_75),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_36),
.C(n_51),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_35),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_51),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_90),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_36),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_60),
.A2(n_42),
.B1(n_37),
.B2(n_34),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_32),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_71),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_78),
.A2(n_42),
.B1(n_37),
.B2(n_34),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_100),
.A2(n_107),
.B1(n_82),
.B2(n_53),
.Y(n_118)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_35),
.B(n_58),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_82),
.B(n_93),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_106),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_74),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_74),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_109),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_90),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_115),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_53),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_84),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_SL g113 ( 
.A1(n_84),
.A2(n_13),
.A3(n_11),
.B1(n_9),
.B2(n_8),
.C1(n_5),
.C2(n_7),
.Y(n_113)
);

AOI322xp5_ASAP7_75t_SL g128 ( 
.A1(n_113),
.A2(n_13),
.A3(n_9),
.B1(n_95),
.B2(n_91),
.C1(n_5),
.C2(n_7),
.Y(n_128)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_116),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_35),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_127),
.B1(n_100),
.B2(n_123),
.Y(n_135)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_125),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_112),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_124),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_127)
);

NAND3xp33_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_1),
.C(n_2),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_111),
.B(n_83),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_129),
.B(n_83),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_101),
.Y(n_131)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_130),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_137),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_135),
.A2(n_142),
.B1(n_123),
.B2(n_126),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_136),
.A2(n_141),
.B(n_99),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_121),
.B(n_94),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_101),
.B(n_107),
.C(n_81),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_115),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_117),
.C(n_129),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_148),
.C(n_150),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_146),
.A2(n_149),
.B(n_151),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_140),
.A2(n_131),
.B1(n_117),
.B2(n_120),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_152),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_143),
.B(n_110),
.Y(n_148)
);

NOR2xp67_ASAP7_75t_SL g149 ( 
.A(n_136),
.B(n_121),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_142),
.A2(n_119),
.B1(n_127),
.B2(n_116),
.Y(n_151)
);

NAND3xp33_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_139),
.C(n_135),
.Y(n_153)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_138),
.B(n_134),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_159),
.B(n_96),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_132),
.C(n_105),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_148),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_145),
.A2(n_99),
.B(n_92),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_160),
.B(n_162),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_161),
.B(n_1),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_158),
.A2(n_96),
.B1(n_47),
.B2(n_24),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_68),
.B1(n_24),
.B2(n_19),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_163),
.A2(n_19),
.B1(n_24),
.B2(n_32),
.Y(n_168)
);

O2A1O1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_156),
.A2(n_32),
.B(n_58),
.C(n_4),
.Y(n_165)
);

AO22x1_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_1),
.B1(n_3),
.B2(n_74),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_168),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_160),
.C(n_161),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_167),
.A2(n_164),
.B(n_165),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_171),
.A2(n_172),
.B(n_166),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_173),
.A2(n_174),
.B(n_3),
.Y(n_175)
);

MAJx2_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_168),
.C(n_3),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_19),
.Y(n_176)
);


endmodule