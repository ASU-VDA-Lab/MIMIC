module fake_jpeg_15178_n_304 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_304);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_304;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

INVx8_ASAP7_75t_SL g42 ( 
.A(n_12),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_43),
.B(n_71),
.Y(n_83)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx5_ASAP7_75t_SL g112 ( 
.A(n_46),
.Y(n_112)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_49),
.B(n_61),
.Y(n_130)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx5_ASAP7_75t_SL g114 ( 
.A(n_51),
.Y(n_114)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_63),
.Y(n_82)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_65),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_28),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_67),
.Y(n_100)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_70),
.Y(n_101)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_0),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_17),
.B(n_1),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_39),
.Y(n_84)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_75),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_16),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_80),
.Y(n_115)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_17),
.B(n_1),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_79),
.B(n_32),
.Y(n_109)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_84),
.B(n_92),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_68),
.A2(n_21),
.B1(n_35),
.B2(n_34),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_85),
.A2(n_86),
.B1(n_112),
.B2(n_81),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_55),
.A2(n_25),
.B1(n_35),
.B2(n_34),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_60),
.A2(n_31),
.B1(n_38),
.B2(n_33),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_89),
.A2(n_96),
.B1(n_122),
.B2(n_123),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_30),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_52),
.A2(n_38),
.B1(n_31),
.B2(n_19),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_43),
.B(n_30),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_97),
.B(n_105),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g99 ( 
.A(n_46),
.B(n_19),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_99),
.A2(n_107),
.B1(n_112),
.B2(n_93),
.Y(n_152)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_103),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_39),
.Y(n_105)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

NOR2x1_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_63),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_78),
.A2(n_33),
.B(n_32),
.C(n_26),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_86),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_109),
.B(n_121),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_65),
.B(n_26),
.Y(n_116)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_59),
.B(n_25),
.Y(n_117)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_117),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_48),
.B(n_3),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_50),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_56),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_74),
.B(n_14),
.Y(n_124)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_124),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_57),
.B(n_15),
.Y(n_127)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_43),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_85),
.B1(n_102),
.B2(n_118),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_9),
.Y(n_131)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_131),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_11),
.C(n_107),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_145),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_83),
.B(n_96),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_135),
.B(n_149),
.Y(n_176)
);

NAND2xp33_ASAP7_75t_SL g136 ( 
.A(n_99),
.B(n_128),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_SL g179 ( 
.A(n_136),
.B(n_139),
.C(n_146),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_140),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_147),
.Y(n_183)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_142),
.Y(n_193)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_143),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_82),
.C(n_115),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_81),
.A2(n_102),
.B1(n_108),
.B2(n_106),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_148),
.A2(n_163),
.B1(n_160),
.B2(n_143),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_101),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_88),
.Y(n_151)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_111),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_89),
.B(n_95),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_153),
.B(n_154),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_130),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_93),
.B(n_113),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_155),
.B(n_158),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_162),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_90),
.B(n_126),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_114),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

BUFx24_ASAP7_75t_L g164 ( 
.A(n_114),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_164),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_87),
.B(n_118),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_167),
.B(n_169),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_87),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_88),
.Y(n_170)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_120),
.Y(n_172)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_111),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_170),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_194),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_178),
.A2(n_190),
.B(n_177),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_138),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_191),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_185),
.A2(n_188),
.B1(n_204),
.B2(n_200),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_152),
.A2(n_138),
.B1(n_136),
.B2(n_134),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_145),
.B(n_172),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_132),
.B(n_144),
.Y(n_191)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_198),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_205),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_133),
.A2(n_173),
.B1(n_161),
.B2(n_151),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_142),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_206),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_187),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_216),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_176),
.B(n_159),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_208),
.B(n_191),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_178),
.A2(n_164),
.B(n_147),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_209),
.A2(n_175),
.B(n_196),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_181),
.A2(n_178),
.B1(n_189),
.B2(n_190),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_212),
.A2(n_194),
.B1(n_204),
.B2(n_200),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_165),
.C(n_157),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_224),
.C(n_193),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_174),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_214),
.Y(n_247)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_215),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_195),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_201),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_217),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_168),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_227),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_184),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_221),
.A2(n_192),
.B1(n_177),
.B2(n_185),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_201),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_223),
.Y(n_243)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_179),
.B(n_166),
.Y(n_224)
);

O2A1O1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_179),
.A2(n_164),
.B(n_137),
.C(n_150),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_225),
.A2(n_228),
.B(n_205),
.Y(n_231)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_203),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_184),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_188),
.B(n_133),
.Y(n_227)
);

NOR2x1_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_140),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_177),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_231),
.A2(n_242),
.B(n_209),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_232),
.B(n_241),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_234),
.B(n_249),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_236),
.A2(n_227),
.B1(n_212),
.B2(n_218),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_244),
.C(n_246),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_230),
.A2(n_183),
.B(n_180),
.Y(n_242)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_245),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_175),
.C(n_199),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_248),
.A2(n_228),
.B(n_225),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_196),
.Y(n_249)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_251),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_234),
.B(n_219),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_253),
.B(n_262),
.Y(n_274)
);

AOI322xp5_ASAP7_75t_L g269 ( 
.A1(n_255),
.A2(n_235),
.A3(n_241),
.B1(n_243),
.B2(n_237),
.C1(n_238),
.C2(n_233),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_256),
.B(n_258),
.Y(n_272)
);

BUFx24_ASAP7_75t_SL g257 ( 
.A(n_247),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_259),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_236),
.A2(n_228),
.B1(n_221),
.B2(n_218),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_250),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_213),
.C(n_223),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_264),
.C(n_246),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_211),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_217),
.C(n_226),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_239),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_222),
.C(n_216),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_273),
.C(n_261),
.Y(n_278)
);

NOR3xp33_ASAP7_75t_SL g267 ( 
.A(n_252),
.B(n_242),
.C(n_231),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_268),
.Y(n_282)
);

A2O1A1Ixp33_ASAP7_75t_L g268 ( 
.A1(n_256),
.A2(n_235),
.B(n_248),
.C(n_238),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_269),
.B(n_275),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_233),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_254),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_237),
.C(n_220),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_270),
.A2(n_251),
.B1(n_264),
.B2(n_265),
.Y(n_277)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_280),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_272),
.A2(n_254),
.B1(n_259),
.B2(n_207),
.Y(n_279)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_279),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_267),
.A2(n_263),
.B(n_215),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_281),
.B(n_284),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_271),
.C(n_266),
.Y(n_284)
);

AOI21x1_ASAP7_75t_L g285 ( 
.A1(n_268),
.A2(n_206),
.B(n_250),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_274),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_286),
.A2(n_290),
.B(n_292),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_220),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_291),
.Y(n_296)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_285),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_289),
.A2(n_282),
.B(n_283),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_293),
.A2(n_294),
.B(n_287),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_288),
.A2(n_277),
.B1(n_281),
.B2(n_280),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_297),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_276),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_296),
.B(n_294),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_300),
.C(n_284),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_298),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_301),
.B(n_302),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_278),
.Y(n_304)
);


endmodule