module fake_jpeg_32120_n_529 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_529);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_529;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_57),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_61),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_63),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_64),
.Y(n_144)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_65),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_29),
.B(n_7),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_66),
.B(n_79),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_67),
.Y(n_151)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g122 ( 
.A(n_70),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_73),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_17),
.B(n_7),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_74),
.B(n_75),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_17),
.B(n_7),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_76),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_77),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_78),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_19),
.B(n_9),
.C(n_2),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_22),
.B(n_9),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_85),
.Y(n_110)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_81),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_83),
.Y(n_148)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_22),
.B(n_9),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_6),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_100),
.Y(n_136)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_88),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_93),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

BUFx24_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_99),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_24),
.B(n_30),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_47),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_24),
.B(n_30),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_103),
.B(n_37),
.Y(n_124)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_104),
.Y(n_153)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_105),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_106),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_36),
.Y(n_107)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_107),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_108),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_109),
.A2(n_68),
.B1(n_58),
.B2(n_71),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_86),
.A2(n_56),
.B1(n_106),
.B2(n_101),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_112),
.A2(n_130),
.B1(n_155),
.B2(n_168),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_124),
.B(n_157),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_62),
.A2(n_45),
.B1(n_44),
.B2(n_34),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_L g134 ( 
.A1(n_57),
.A2(n_25),
.B(n_47),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_140),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_64),
.A2(n_21),
.B1(n_43),
.B2(n_32),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_156),
.A2(n_164),
.B1(n_82),
.B2(n_39),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_78),
.B(n_26),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_78),
.B(n_37),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_166),
.Y(n_206)
);

OA22x2_ASAP7_75t_L g164 ( 
.A1(n_72),
.A2(n_44),
.B1(n_45),
.B2(n_50),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_73),
.B(n_26),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_96),
.A2(n_36),
.B1(n_45),
.B2(n_44),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_59),
.B(n_18),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_27),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_96),
.A2(n_100),
.B1(n_67),
.B2(n_76),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_170),
.A2(n_89),
.B1(n_97),
.B2(n_94),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_100),
.B(n_18),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_34),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_175),
.Y(n_236)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_127),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_176),
.Y(n_226)
);

INVx11_ASAP7_75t_L g177 ( 
.A(n_128),
.Y(n_177)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_177),
.Y(n_246)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_118),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_179),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_L g180 ( 
.A1(n_117),
.A2(n_99),
.B1(n_77),
.B2(n_83),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_180),
.A2(n_188),
.B1(n_192),
.B2(n_132),
.Y(n_238)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_125),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_181),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_182),
.B(n_189),
.Y(n_234)
);

BUFx16f_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_183),
.Y(n_263)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_184),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_125),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_185),
.Y(n_233)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_114),
.Y(n_186)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_186),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_187),
.A2(n_221),
.B1(n_122),
.B2(n_138),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_126),
.B(n_21),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_111),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_190),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_191),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_161),
.A2(n_88),
.B1(n_25),
.B2(n_50),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_136),
.A2(n_20),
.B1(n_43),
.B2(n_27),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_193),
.A2(n_156),
.B1(n_170),
.B2(n_168),
.Y(n_227)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_121),
.Y(n_194)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_194),
.Y(n_240)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_113),
.Y(n_195)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_195),
.Y(n_243)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_143),
.Y(n_196)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_196),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_110),
.B(n_32),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_197),
.Y(n_260)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_198),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_150),
.Y(n_199)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_199),
.Y(n_259)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_127),
.Y(n_200)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_200),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_133),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_201),
.B(n_202),
.Y(n_250)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_116),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_131),
.Y(n_203)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_203),
.Y(n_255)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_153),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_204),
.Y(n_261)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_142),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_205),
.Y(n_232)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_129),
.Y(n_207)
);

BUFx4f_ASAP7_75t_L g251 ( 
.A(n_207),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_208),
.Y(n_249)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_149),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_241)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_135),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_146),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_115),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_133),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_214),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_161),
.B(n_45),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_164),
.B(n_11),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_216),
.Y(n_237)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_120),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_129),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_217),
.A2(n_224),
.B1(n_165),
.B2(n_148),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_160),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_219),
.Y(n_247)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_139),
.Y(n_219)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_128),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_222),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_137),
.B(n_109),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_119),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_152),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_225),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_144),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_159),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_227),
.A2(n_262),
.B1(n_180),
.B2(n_220),
.Y(n_275)
);

A2O1A1Ixp33_ASAP7_75t_L g231 ( 
.A1(n_173),
.A2(n_164),
.B(n_130),
.C(n_39),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_231),
.B(n_195),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_235),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_238),
.B(n_239),
.Y(n_276)
);

NAND2x1_ASAP7_75t_L g239 ( 
.A(n_178),
.B(n_39),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_215),
.A2(n_148),
.B1(n_165),
.B2(n_138),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_245),
.A2(n_181),
.B1(n_207),
.B2(n_185),
.Y(n_289)
);

NOR2xp67_ASAP7_75t_L g254 ( 
.A(n_174),
.B(n_132),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_187),
.A2(n_119),
.B(n_139),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_257),
.A2(n_200),
.B(n_176),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_237),
.A2(n_206),
.B(n_191),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_266),
.A2(n_278),
.B(n_288),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_267),
.A2(n_286),
.B(n_241),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_250),
.Y(n_268)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_268),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_250),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_269),
.B(n_272),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_256),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_273),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_237),
.B(n_229),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_274),
.B(n_285),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_275),
.A2(n_277),
.B1(n_283),
.B2(n_251),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_239),
.A2(n_184),
.B1(n_167),
.B2(n_151),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_229),
.A2(n_186),
.B(n_177),
.Y(n_278)
);

FAx1_ASAP7_75t_SL g279 ( 
.A(n_245),
.B(n_183),
.CI(n_223),
.CON(n_279),
.SN(n_279)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_279),
.B(n_289),
.Y(n_313)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_256),
.Y(n_280)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_280),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_233),
.Y(n_281)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_281),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_226),
.A2(n_141),
.B1(n_175),
.B2(n_199),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_282),
.A2(n_287),
.B1(n_291),
.B2(n_295),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_239),
.A2(n_144),
.B1(n_151),
.B2(n_167),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_247),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_284),
.B(n_290),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_253),
.B(n_225),
.Y(n_285)
);

A2O1A1Ixp33_ASAP7_75t_SL g286 ( 
.A1(n_257),
.A2(n_183),
.B(n_122),
.C(n_224),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_226),
.A2(n_141),
.B1(n_219),
.B2(n_212),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_253),
.A2(n_218),
.B(n_123),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_247),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_264),
.A2(n_216),
.B1(n_162),
.B2(n_147),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_249),
.B(n_209),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_292),
.B(n_293),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_238),
.A2(n_205),
.B1(n_203),
.B2(n_217),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_246),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_294),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_264),
.A2(n_246),
.B1(n_227),
.B2(n_258),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_236),
.A2(n_145),
.B1(n_115),
.B2(n_108),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_296),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_234),
.B(n_0),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_297),
.B(n_298),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_252),
.B(n_0),
.Y(n_298)
);

INVxp33_ASAP7_75t_L g299 ( 
.A(n_267),
.Y(n_299)
);

INVxp33_ASAP7_75t_L g351 ( 
.A(n_299),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_244),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_301),
.B(n_297),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_298),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_302),
.B(n_304),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_268),
.B(n_260),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_280),
.B(n_231),
.C(n_240),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_306),
.B(n_325),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_276),
.A2(n_236),
.B(n_259),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_310),
.A2(n_311),
.B(n_317),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_276),
.A2(n_259),
.B(n_261),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_272),
.B(n_252),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_314),
.B(n_329),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_315),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_276),
.A2(n_261),
.B(n_232),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_285),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_318),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_322),
.A2(n_327),
.B1(n_293),
.B2(n_289),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_276),
.A2(n_232),
.B(n_244),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_323),
.A2(n_286),
.B(n_279),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_266),
.B(n_240),
.C(n_242),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_292),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_326),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_275),
.A2(n_232),
.B1(n_265),
.B2(n_248),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_273),
.B(n_243),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_314),
.Y(n_330)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_330),
.Y(n_363)
);

MAJx2_ASAP7_75t_L g334 ( 
.A(n_312),
.B(n_268),
.C(n_269),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_334),
.B(n_344),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_301),
.B(n_278),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_335),
.B(n_306),
.C(n_325),
.Y(n_370)
);

OAI22xp33_ASAP7_75t_L g336 ( 
.A1(n_315),
.A2(n_286),
.B1(n_295),
.B2(n_279),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_336),
.A2(n_357),
.B1(n_311),
.B2(n_310),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_313),
.A2(n_271),
.B1(n_283),
.B2(n_277),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g381 ( 
.A1(n_337),
.A2(n_359),
.B1(n_309),
.B2(n_322),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_303),
.A2(n_288),
.B(n_286),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_338),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_339),
.A2(n_324),
.B1(n_308),
.B2(n_329),
.Y(n_371)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_307),
.Y(n_340)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_340),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_341),
.B(n_343),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_304),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_342),
.B(n_350),
.Y(n_375)
);

AO22x1_ASAP7_75t_SL g343 ( 
.A1(n_307),
.A2(n_286),
.B1(n_279),
.B2(n_270),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_303),
.B(n_286),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_346),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_303),
.B(n_287),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_348),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_300),
.A2(n_327),
.B1(n_322),
.B2(n_308),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_349),
.A2(n_316),
.B1(n_310),
.B2(n_317),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_317),
.A2(n_294),
.B(n_282),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_312),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_352),
.B(n_356),
.Y(n_369)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_307),
.Y(n_354)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_354),
.Y(n_377)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_324),
.Y(n_355)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_355),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_321),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_313),
.A2(n_296),
.B1(n_294),
.B2(n_228),
.Y(n_357)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_305),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_319),
.B(n_294),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_360),
.B(n_329),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_358),
.B(n_325),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_361),
.B(n_370),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_347),
.B(n_321),
.Y(n_362)
);

CKINVDCx14_ASAP7_75t_R g413 ( 
.A(n_362),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_354),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_368),
.B(n_378),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_371),
.A2(n_373),
.B1(n_376),
.B2(n_348),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_355),
.A2(n_326),
.B1(n_318),
.B2(n_324),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_332),
.B(n_302),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_374),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_358),
.B(n_301),
.C(n_306),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_379),
.A2(n_386),
.B1(n_350),
.B2(n_349),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_330),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_380),
.B(n_391),
.Y(n_411)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_381),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_331),
.B(n_320),
.Y(n_382)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_382),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_335),
.B(n_319),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g400 ( 
.A(n_384),
.B(n_390),
.Y(n_400)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_385),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_336),
.A2(n_327),
.B1(n_323),
.B2(n_311),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_344),
.B(n_319),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_387),
.B(n_341),
.Y(n_401)
);

INVx13_ASAP7_75t_L g389 ( 
.A(n_351),
.Y(n_389)
);

INVx13_ASAP7_75t_L g393 ( 
.A(n_389),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_334),
.B(n_345),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_360),
.B(n_323),
.C(n_328),
.Y(n_391)
);

INVxp33_ASAP7_75t_L g394 ( 
.A(n_369),
.Y(n_394)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_394),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_366),
.A2(n_353),
.B(n_338),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_395),
.A2(n_333),
.B(n_315),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_396),
.A2(n_408),
.B1(n_379),
.B2(n_386),
.Y(n_426)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_374),
.Y(n_398)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_398),
.Y(n_425)
);

NOR3xp33_ASAP7_75t_L g399 ( 
.A(n_375),
.B(n_320),
.C(n_345),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_399),
.B(n_402),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_401),
.B(n_409),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_364),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_362),
.B(n_343),
.Y(n_404)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_404),
.Y(n_431)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_377),
.Y(n_405)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_405),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_390),
.B(n_328),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_406),
.B(n_410),
.Y(n_441)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_377),
.Y(n_407)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_407),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_371),
.A2(n_348),
.B1(n_357),
.B2(n_353),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_370),
.B(n_346),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_363),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_363),
.B(n_328),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_414),
.B(n_415),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_378),
.B(n_387),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_373),
.B(n_343),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_416),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_417),
.A2(n_366),
.B1(n_388),
.B2(n_346),
.Y(n_428)
);

BUFx24_ASAP7_75t_SL g419 ( 
.A(n_365),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_419),
.A2(n_365),
.B1(n_230),
.B2(n_243),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_423),
.B(n_437),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_426),
.A2(n_435),
.B1(n_436),
.B2(n_398),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_409),
.B(n_401),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_427),
.B(n_434),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_428),
.B(n_430),
.Y(n_444)
);

FAx1_ASAP7_75t_SL g433 ( 
.A(n_404),
.B(n_372),
.CI(n_364),
.CON(n_433),
.SN(n_433)
);

OR2x2_ASAP7_75t_L g460 ( 
.A(n_433),
.B(n_416),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_400),
.B(n_372),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_413),
.A2(n_339),
.B1(n_316),
.B2(n_383),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_420),
.A2(n_383),
.B1(n_385),
.B2(n_391),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_392),
.A2(n_388),
.B1(n_367),
.B2(n_384),
.Y(n_437)
);

XOR2x2_ASAP7_75t_SL g438 ( 
.A(n_402),
.B(n_367),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_438),
.B(n_395),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_392),
.A2(n_361),
.B1(n_351),
.B2(n_333),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_440),
.B(n_443),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_400),
.B(n_389),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_429),
.B(n_397),
.C(n_427),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_446),
.B(n_447),
.C(n_450),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_429),
.B(n_397),
.C(n_403),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_448),
.B(n_437),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_425),
.A2(n_412),
.B1(n_418),
.B2(n_405),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_449),
.B(n_454),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_451),
.B(n_428),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_SL g452 ( 
.A1(n_438),
.A2(n_410),
.B1(n_407),
.B2(n_408),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_452),
.A2(n_430),
.B(n_426),
.Y(n_463)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_439),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_432),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_455),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_443),
.B(n_411),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_456),
.B(n_458),
.Y(n_464)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_424),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_457),
.A2(n_459),
.B1(n_462),
.B2(n_309),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_441),
.B(n_396),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_442),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_460),
.A2(n_440),
.B(n_421),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_431),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_461),
.B(n_433),
.Y(n_474)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_422),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g492 ( 
.A(n_463),
.B(n_465),
.Y(n_492)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_467),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_445),
.A2(n_394),
.B1(n_433),
.B2(n_393),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_468),
.B(n_474),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_444),
.A2(n_453),
.B1(n_451),
.B2(n_452),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_469),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_470),
.B(n_475),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_471),
.B(n_472),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_SL g473 ( 
.A(n_453),
.B(n_434),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_473),
.B(n_263),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_447),
.B(n_446),
.C(n_444),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_450),
.B(n_393),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_476),
.B(n_263),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_460),
.B(n_359),
.C(n_305),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_477),
.A2(n_255),
.B(n_233),
.Y(n_489)
);

FAx1_ASAP7_75t_SL g479 ( 
.A(n_451),
.B(n_251),
.CI(n_305),
.CON(n_479),
.SN(n_479)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_479),
.B(n_228),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_464),
.B(n_281),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_484),
.B(n_485),
.Y(n_502)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_478),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_474),
.B(n_281),
.Y(n_486)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_486),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_469),
.A2(n_251),
.B1(n_242),
.B2(n_230),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_488),
.B(n_490),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_489),
.B(n_494),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_491),
.B(n_493),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_472),
.B(n_255),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_483),
.A2(n_475),
.B(n_470),
.Y(n_495)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_495),
.B(n_480),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_487),
.B(n_471),
.C(n_477),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_496),
.B(n_504),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_SL g498 ( 
.A(n_492),
.B(n_473),
.Y(n_498)
);

OA21x2_ASAP7_75t_L g510 ( 
.A1(n_498),
.A2(n_499),
.B(n_491),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_487),
.A2(n_466),
.B(n_476),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_492),
.B(n_479),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_501),
.B(n_505),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_482),
.B(n_2),
.C(n_3),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_481),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_496),
.B(n_482),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_507),
.B(n_509),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_510),
.B(n_512),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_502),
.B(n_3),
.Y(n_511)
);

O2A1O1Ixp33_ASAP7_75t_SL g519 ( 
.A1(n_511),
.A2(n_503),
.B(n_10),
.C(n_11),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_506),
.B(n_3),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_504),
.B(n_5),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_513),
.B(n_5),
.Y(n_515)
);

A2O1A1Ixp33_ASAP7_75t_SL g520 ( 
.A1(n_515),
.A2(n_519),
.B(n_5),
.C(n_10),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_514),
.A2(n_500),
.B(n_498),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_518),
.A2(n_508),
.B(n_503),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_520),
.B(n_521),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_516),
.A2(n_497),
.B(n_511),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_522),
.B(n_517),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_524),
.A2(n_497),
.B(n_12),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_523),
.C(n_14),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_526),
.B(n_11),
.C(n_14),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_527),
.B(n_11),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_528),
.B(n_14),
.C(n_16),
.Y(n_529)
);


endmodule