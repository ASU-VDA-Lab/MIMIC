module fake_jpeg_47_n_88 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_88);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_88;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx2_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_23),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_2),
.B(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_19),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_22),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_37),
.Y(n_41)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_28),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_35),
.B1(n_31),
.B2(n_26),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_28),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_30),
.Y(n_44)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_32),
.B(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_42),
.Y(n_53)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_45),
.B1(n_31),
.B2(n_25),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_37),
.B(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

AO22x2_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_50),
.Y(n_55)
);

AND2x6_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_12),
.Y(n_47)
);

NOR3xp33_ASAP7_75t_SL g59 ( 
.A(n_47),
.B(n_52),
.C(n_4),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_27),
.C(n_20),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_4),
.Y(n_58)
);

AND2x6_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_18),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_56),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_43),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_57),
.B(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_58),
.B(n_60),
.Y(n_63)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_43),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_15),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_46),
.B1(n_45),
.B2(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_46),
.B1(n_45),
.B2(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_59),
.C(n_17),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_6),
.C(n_7),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_13),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_69),
.B(n_5),
.Y(n_72)
);

OAI32xp33_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_74),
.C(n_76),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_72),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_65),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_73),
.A2(n_66),
.B1(n_63),
.B2(n_68),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_71),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_81),
.A2(n_82),
.B(n_77),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_80),
.B(n_75),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_79),
.B(n_67),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

NOR3xp33_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_76),
.C(n_9),
.Y(n_86)
);

MAJx2_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_8),
.C(n_9),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_10),
.Y(n_88)
);


endmodule