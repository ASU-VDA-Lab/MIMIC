module real_aes_4524_n_375 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_1285, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_1286, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_375);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_1285;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_1286;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_375;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_830;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_592;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_400;
wire n_1160;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_417;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_527;
wire n_552;
wire n_590;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1250;
wire n_1095;
wire n_859;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_749;
wire n_914;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1161;
wire n_686;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_837;
wire n_829;
wire n_1030;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_1004;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1129;
wire n_742;
wire n_1014;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_510;
wire n_550;
wire n_966;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_807;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1194;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1120;
wire n_689;
wire n_946;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_739;
wire n_1162;
wire n_762;
wire n_442;
wire n_740;
wire n_639;
wire n_1186;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_414;
wire n_776;
wire n_1138;
wire n_890;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_577;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_937;
wire n_773;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_816;
wire n_625;
wire n_953;
wire n_716;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_443;
wire n_1029;
wire n_1207;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_1167;
wire n_609;
wire n_1006;
wire n_1259;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1054;
wire n_1050;
wire n_426;
wire n_1134;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1060;
wire n_1154;
wire n_632;
wire n_714;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1033;
wire n_1028;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1127;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1015;
wire n_863;
wire n_1226;
wire n_525;
wire n_644;
wire n_1150;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1240;
wire n_987;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_555;
wire n_974;
wire n_857;
wire n_376;
wire n_491;
wire n_1110;
wire n_1137;
wire n_460;
wire n_666;
wire n_660;
wire n_886;
wire n_767;
wire n_889;
wire n_379;
wire n_1021;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1198;
wire n_993;
wire n_819;
wire n_737;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_449;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1252;
wire n_430;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1273;
wire n_959;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_1183;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_698;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_483;
wire n_394;
wire n_1280;
wire n_729;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_603;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_0), .A2(n_259), .B1(n_517), .B2(n_526), .Y(n_873) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1), .Y(n_1227) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_2), .A2(n_357), .B1(n_520), .B2(n_521), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_3), .A2(n_8), .B1(n_950), .B2(n_951), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_4), .A2(n_86), .B1(n_454), .B2(n_592), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_5), .A2(n_193), .B1(n_518), .B2(n_524), .Y(n_872) );
AOI22xp5_ASAP7_75t_L g810 ( .A1(n_6), .A2(n_200), .B1(n_551), .B2(n_590), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_7), .A2(n_152), .B1(n_520), .B2(n_521), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_9), .A2(n_166), .B1(n_445), .B2(n_450), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_10), .A2(n_321), .B1(n_518), .B2(n_524), .Y(n_633) );
AOI22xp33_ASAP7_75t_SL g916 ( .A1(n_11), .A2(n_256), .B1(n_760), .B2(n_917), .Y(n_916) );
INVx1_ASAP7_75t_L g735 ( .A(n_12), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g1235 ( .A1(n_13), .A2(n_153), .B1(n_773), .B2(n_1236), .Y(n_1235) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_14), .A2(n_335), .B1(n_445), .B2(n_702), .Y(n_831) );
AOI22xp5_ASAP7_75t_L g839 ( .A1(n_15), .A2(n_304), .B1(n_461), .B2(n_477), .Y(n_839) );
AOI221xp5_ASAP7_75t_L g1223 ( .A1(n_16), .A2(n_286), .B1(n_541), .B2(n_1224), .C(n_1226), .Y(n_1223) );
AOI22xp33_ASAP7_75t_L g1261 ( .A1(n_17), .A2(n_32), .B1(n_755), .B2(n_1239), .Y(n_1261) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_18), .A2(n_114), .B1(n_451), .B2(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_19), .B(n_405), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_20), .A2(n_197), .B1(n_474), .B2(n_477), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_21), .A2(n_264), .B1(n_954), .B2(n_955), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_22), .A2(n_245), .B1(n_520), .B2(n_521), .Y(n_727) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_23), .A2(n_207), .B1(n_504), .B2(n_527), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g1271 ( .A(n_24), .B(n_1272), .Y(n_1271) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_25), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_26), .A2(n_337), .B1(n_712), .B2(n_797), .Y(n_796) );
AOI22xp5_ASAP7_75t_L g995 ( .A1(n_27), .A2(n_269), .B1(n_996), .B2(n_998), .Y(n_995) );
AOI22xp5_ASAP7_75t_L g1270 ( .A1(n_28), .A2(n_78), .B1(n_934), .B2(n_1236), .Y(n_1270) );
AOI22xp5_ASAP7_75t_L g836 ( .A1(n_29), .A2(n_151), .B1(n_699), .B2(n_837), .Y(n_836) );
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_30), .A2(n_688), .B(n_689), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_31), .A2(n_46), .B1(n_749), .B2(n_751), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g1013 ( .A1(n_33), .A2(n_204), .B1(n_996), .B2(n_998), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_34), .A2(n_147), .B1(n_398), .B2(n_423), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_35), .A2(n_353), .B1(n_1000), .B2(n_1006), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_36), .A2(n_212), .B1(n_505), .B2(n_510), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_37), .A2(n_211), .B1(n_983), .B2(n_987), .Y(n_982) );
INVxp33_ASAP7_75t_SL g1039 ( .A(n_38), .Y(n_1039) );
AOI21xp5_ASAP7_75t_L g921 ( .A1(n_39), .A2(n_922), .B(n_924), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_40), .A2(n_55), .B1(n_990), .B2(n_993), .Y(n_989) );
INVx1_ASAP7_75t_L g925 ( .A(n_41), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_42), .A2(n_104), .B1(n_526), .B2(n_527), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_43), .A2(n_372), .B1(n_504), .B2(n_527), .Y(n_826) );
XOR2x2_ASAP7_75t_L g603 ( .A(n_44), .B(n_604), .Y(n_603) );
AOI22xp33_ASAP7_75t_SL g869 ( .A1(n_45), .A2(n_360), .B1(n_505), .B2(n_712), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_47), .A2(n_54), .B1(n_754), .B2(n_755), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_48), .A2(n_150), .B1(n_445), .B2(n_553), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_49), .A2(n_113), .B1(n_474), .B2(n_477), .Y(n_473) );
INVx1_ASAP7_75t_L g710 ( .A(n_50), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_51), .A2(n_138), .B1(n_474), .B2(n_477), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_52), .A2(n_160), .B1(n_627), .B2(n_800), .Y(n_799) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_53), .A2(n_98), .B1(n_428), .B2(n_677), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_56), .A2(n_167), .B1(n_704), .B2(n_750), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_57), .A2(n_179), .B1(n_555), .B2(n_706), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_58), .A2(n_109), .B1(n_520), .B2(n_521), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_59), .A2(n_235), .B1(n_518), .B2(n_524), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_60), .A2(n_253), .B1(n_523), .B2(n_567), .Y(n_566) );
OA22x2_ASAP7_75t_L g411 ( .A1(n_61), .A2(n_164), .B1(n_405), .B2(n_409), .Y(n_411) );
INVx1_ASAP7_75t_L g440 ( .A(n_61), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_62), .A2(n_310), .B1(n_699), .B2(n_700), .Y(n_698) );
XNOR2x1_ASAP7_75t_L g673 ( .A(n_63), .B(n_674), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g999 ( .A1(n_63), .A2(n_287), .B1(n_1000), .B2(n_1001), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_64), .A2(n_70), .B1(n_782), .B2(n_783), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_65), .A2(n_67), .B1(n_520), .B2(n_521), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_66), .A2(n_299), .B1(n_551), .B2(n_590), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_68), .A2(n_356), .B1(n_685), .B2(n_841), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_69), .A2(n_257), .B1(n_553), .B2(n_704), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_71), .A2(n_249), .B1(n_507), .B2(n_508), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_72), .A2(n_303), .B1(n_520), .B2(n_521), .Y(n_663) );
INVx1_ASAP7_75t_L g1117 ( .A(n_73), .Y(n_1117) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_74), .A2(n_260), .B1(n_549), .B2(n_702), .Y(n_792) );
INVx1_ASAP7_75t_L g885 ( .A(n_75), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_76), .A2(n_108), .B1(n_549), .B2(n_551), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_77), .A2(n_262), .B1(n_504), .B2(n_527), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g605 ( .A1(n_79), .A2(n_187), .B1(n_606), .B2(n_607), .C(n_608), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_80), .B(n_181), .Y(n_384) );
INVx1_ASAP7_75t_L g408 ( .A(n_80), .Y(n_408) );
OAI21xp33_ASAP7_75t_L g441 ( .A1(n_80), .A2(n_164), .B(n_442), .Y(n_441) );
AOI21xp33_ASAP7_75t_L g1267 ( .A1(n_81), .A2(n_541), .B(n_1268), .Y(n_1267) );
AOI221xp5_ASAP7_75t_L g598 ( .A1(n_82), .A2(n_314), .B1(n_541), .B2(n_599), .C(n_600), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_83), .A2(n_351), .B1(n_520), .B2(n_521), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_84), .A2(n_300), .B1(n_505), .B2(n_507), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g1262 ( .A1(n_85), .A2(n_278), .B1(n_760), .B2(n_761), .Y(n_1262) );
INVx1_ASAP7_75t_L g659 ( .A(n_87), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_88), .A2(n_185), .B1(n_428), .B2(n_547), .Y(n_546) );
AOI22xp33_ASAP7_75t_SL g1263 ( .A1(n_89), .A2(n_215), .B1(n_428), .B2(n_837), .Y(n_1263) );
INVx1_ASAP7_75t_L g803 ( .A(n_90), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_91), .A2(n_131), .B1(n_754), .B2(n_755), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_92), .B(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_93), .B(n_841), .Y(n_891) );
INVxp33_ASAP7_75t_L g1032 ( .A(n_94), .Y(n_1032) );
AND2x4_ASAP7_75t_L g986 ( .A(n_95), .B(n_273), .Y(n_986) );
INVx1_ASAP7_75t_L g992 ( .A(n_95), .Y(n_992) );
HB1xp67_ASAP7_75t_L g1282 ( .A(n_95), .Y(n_1282) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_96), .A2(n_316), .B1(n_504), .B2(n_527), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_97), .A2(n_239), .B1(n_450), .B2(n_837), .Y(n_898) );
INVx1_ASAP7_75t_L g845 ( .A(n_99), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_100), .A2(n_220), .B1(n_445), .B2(n_681), .Y(n_680) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_101), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g1257 ( .A1(n_102), .A2(n_103), .B1(n_897), .B2(n_1258), .Y(n_1257) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_105), .A2(n_195), .B1(n_508), .B2(n_625), .Y(n_822) );
INVx1_ASAP7_75t_L g970 ( .A(n_106), .Y(n_970) );
AOI221xp5_ASAP7_75t_L g842 ( .A1(n_107), .A2(n_111), .B1(n_773), .B2(n_817), .C(n_843), .Y(n_842) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_110), .A2(n_523), .B(n_709), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g1234 ( .A1(n_112), .A2(n_128), .B1(n_461), .B2(n_782), .Y(n_1234) );
XNOR2x1_ASAP7_75t_L g880 ( .A(n_115), .B(n_881), .Y(n_880) );
AOI21xp5_ASAP7_75t_L g816 ( .A1(n_116), .A2(n_817), .B(n_819), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_117), .A2(n_322), .B1(n_523), .B2(n_524), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_118), .B(n_537), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_119), .A2(n_154), .B1(n_555), .B2(n_948), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_120), .A2(n_202), .B1(n_474), .B2(n_477), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_121), .A2(n_155), .B1(n_454), .B2(n_456), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_122), .A2(n_180), .B1(n_505), .B2(n_508), .Y(n_656) );
INVx1_ASAP7_75t_L g844 ( .A(n_123), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_124), .A2(n_142), .B1(n_699), .B2(n_700), .Y(n_789) );
INVx1_ASAP7_75t_L g985 ( .A(n_125), .Y(n_985) );
AND2x4_ASAP7_75t_L g988 ( .A(n_125), .B(n_380), .Y(n_988) );
INVx1_ASAP7_75t_SL g997 ( .A(n_125), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_126), .A2(n_258), .B1(n_477), .B2(n_625), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g1230 ( .A1(n_127), .A2(n_352), .B1(n_677), .B2(n_750), .Y(n_1230) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_129), .A2(n_294), .B1(n_914), .B2(n_915), .Y(n_913) );
XNOR2x2_ASAP7_75t_SL g720 ( .A(n_130), .B(n_721), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g1017 ( .A1(n_130), .A2(n_233), .B1(n_1000), .B2(n_1001), .Y(n_1017) );
INVx1_ASAP7_75t_L g636 ( .A(n_132), .Y(n_636) );
INVx1_ASAP7_75t_L g490 ( .A(n_133), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_134), .B(n_599), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_135), .A2(n_266), .B1(n_454), .B2(n_553), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_136), .A2(n_343), .B1(n_706), .B2(n_757), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_137), .A2(n_355), .B1(n_507), .B2(n_523), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g738 ( .A1(n_139), .A2(n_362), .B1(n_607), .B2(n_739), .C(n_740), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_140), .A2(n_276), .B1(n_983), .B2(n_987), .Y(n_1021) );
XNOR2x1_ASAP7_75t_L g807 ( .A(n_141), .B(n_808), .Y(n_807) );
AO22x1_ASAP7_75t_L g1231 ( .A1(n_143), .A2(n_318), .B1(n_681), .B2(n_760), .Y(n_1231) );
INVx1_ASAP7_75t_L g814 ( .A(n_144), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_145), .A2(n_178), .B1(n_517), .B2(n_526), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_146), .A2(n_361), .B1(n_520), .B2(n_521), .Y(n_630) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_148), .A2(n_541), .B(n_542), .Y(n_540) );
INVx1_ASAP7_75t_L g730 ( .A(n_149), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_156), .B(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g601 ( .A(n_157), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_158), .A2(n_229), .B1(n_535), .B2(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g1020 ( .A1(n_159), .A2(n_371), .B1(n_990), .B2(n_993), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_161), .A2(n_302), .B1(n_398), .B2(n_423), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_162), .A2(n_346), .B1(n_504), .B2(n_527), .Y(n_631) );
INVx1_ASAP7_75t_L g422 ( .A(n_163), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_163), .B(n_218), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_163), .B(n_438), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_164), .B(n_285), .Y(n_383) );
AOI22xp5_ASAP7_75t_L g1016 ( .A1(n_165), .A2(n_173), .B1(n_996), .B2(n_998), .Y(n_1016) );
INVx1_ASAP7_75t_L g1269 ( .A(n_168), .Y(n_1269) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_169), .A2(n_280), .B1(n_461), .B2(n_716), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_170), .A2(n_176), .B1(n_461), .B2(n_463), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_171), .A2(n_240), .B1(n_423), .B2(n_555), .Y(n_835) );
AOI221xp5_ASAP7_75t_L g899 ( .A1(n_172), .A2(n_182), .B1(n_481), .B2(n_773), .C(n_900), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_174), .A2(n_313), .B1(n_749), .B2(n_957), .Y(n_956) );
INVx1_ASAP7_75t_L g543 ( .A(n_175), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g862 ( .A1(n_177), .A2(n_502), .B(n_863), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_181), .B(n_415), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_183), .A2(n_213), .B1(n_553), .B2(n_704), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_184), .A2(n_255), .B1(n_517), .B2(n_526), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_186), .A2(n_373), .B1(n_423), .B2(n_555), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g896 ( .A1(n_188), .A2(n_374), .B1(n_423), .B2(n_897), .Y(n_896) );
AO22x2_ASAP7_75t_L g856 ( .A1(n_189), .A2(n_857), .B1(n_875), .B2(n_876), .Y(n_856) );
INVxp67_ASAP7_75t_SL g875 ( .A(n_189), .Y(n_875) );
INVx1_ASAP7_75t_L g820 ( .A(n_190), .Y(n_820) );
INVx1_ASAP7_75t_L g690 ( .A(n_191), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_192), .A2(n_301), .B1(n_454), .B2(n_833), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_194), .B(n_692), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_196), .B(n_694), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_198), .A2(n_348), .B1(n_461), .B2(n_535), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_199), .A2(n_205), .B1(n_547), .B2(n_587), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_201), .A2(n_394), .B1(n_395), .B2(n_497), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_201), .Y(n_394) );
AOI21xp33_ASAP7_75t_L g801 ( .A1(n_203), .A2(n_625), .B(n_802), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g1119 ( .A1(n_206), .A2(n_263), .B1(n_1006), .B2(n_1037), .Y(n_1119) );
XNOR2x1_ASAP7_75t_L g695 ( .A(n_208), .B(n_696), .Y(n_695) );
AOI22xp33_ASAP7_75t_SL g1014 ( .A1(n_208), .A2(n_275), .B1(n_1000), .B2(n_1001), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_209), .A2(n_363), .B1(n_963), .B2(n_964), .Y(n_962) );
BUFx2_ASAP7_75t_L g865 ( .A(n_210), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g1238 ( .A1(n_214), .A2(n_317), .B1(n_592), .B2(n_1239), .Y(n_1238) );
INVx1_ASAP7_75t_L g901 ( .A(n_216), .Y(n_901) );
AOI22xp5_ASAP7_75t_L g811 ( .A1(n_217), .A2(n_345), .B1(n_704), .B2(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g406 ( .A(n_218), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g1007 ( .A1(n_219), .A2(n_222), .B1(n_996), .B2(n_998), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_221), .A2(n_334), .B1(n_706), .B2(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g1221 ( .A(n_222), .Y(n_1221) );
OAI222xp33_ASAP7_75t_L g1232 ( .A1(n_222), .A2(n_1233), .B1(n_1237), .B2(n_1238), .C1(n_1285), .C2(n_1286), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1243 ( .A(n_222), .B(n_1238), .Y(n_1243) );
AOI22xp33_ASAP7_75t_L g1251 ( .A1(n_222), .A2(n_1252), .B1(n_1278), .B2(n_1280), .Y(n_1251) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_223), .A2(n_368), .B1(n_585), .B2(n_757), .Y(n_756) );
XNOR2x1_ASAP7_75t_L g498 ( .A(n_224), .B(n_499), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g1273 ( .A1(n_225), .A2(n_341), .B1(n_1274), .B2(n_1275), .Y(n_1273) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_226), .A2(n_339), .B1(n_461), .B2(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_227), .A2(n_315), .B1(n_454), .B2(n_592), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_228), .A2(n_282), .B1(n_628), .B2(n_929), .Y(n_928) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_230), .A2(n_238), .B1(n_627), .B2(n_628), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_231), .B(n_502), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g1253 ( .A1(n_232), .A2(n_1254), .B1(n_1276), .B2(n_1277), .Y(n_1253) );
CKINVDCx5p33_ASAP7_75t_R g1276 ( .A(n_232), .Y(n_1276) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_234), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_236), .A2(n_326), .B1(n_549), .B2(n_702), .Y(n_701) );
OR2x2_ASAP7_75t_L g794 ( .A(n_237), .B(n_795), .Y(n_794) );
INVxp67_ASAP7_75t_L g806 ( .A(n_237), .Y(n_806) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_241), .A2(n_261), .B1(n_517), .B2(n_526), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_242), .A2(n_312), .B1(n_428), .B2(n_433), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_243), .A2(n_296), .B1(n_518), .B2(n_524), .Y(n_726) );
INVx1_ASAP7_75t_L g1118 ( .A(n_244), .Y(n_1118) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_246), .B(n_565), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_247), .A2(n_248), .B1(n_555), .B2(n_585), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_250), .A2(n_292), .B1(n_507), .B2(n_508), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_251), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_252), .A2(n_293), .B1(n_553), .B2(n_704), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_254), .A2(n_354), .B1(n_433), .B2(n_587), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_265), .A2(n_279), .B1(n_507), .B2(n_508), .Y(n_562) );
AOI221xp5_ASAP7_75t_L g965 ( .A1(n_267), .A2(n_268), .B1(n_628), .B2(n_966), .C(n_969), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_270), .A2(n_305), .B1(n_517), .B2(n_518), .Y(n_516) );
INVx1_ASAP7_75t_L g737 ( .A(n_271), .Y(n_737) );
AOI22x1_ASAP7_75t_L g580 ( .A1(n_272), .A2(n_581), .B1(n_582), .B2(n_602), .Y(n_580) );
INVx1_ASAP7_75t_L g602 ( .A(n_272), .Y(n_602) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_273), .Y(n_385) );
AND2x4_ASAP7_75t_L g991 ( .A(n_273), .B(n_992), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_274), .B(n_481), .Y(n_480) );
XNOR2x2_ASAP7_75t_L g944 ( .A(n_276), .B(n_945), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_277), .A2(n_309), .B1(n_517), .B2(n_526), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g933 ( .A1(n_281), .A2(n_369), .B1(n_776), .B2(n_934), .Y(n_933) );
INVx1_ASAP7_75t_L g887 ( .A(n_283), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_284), .A2(n_327), .B1(n_505), .B2(n_523), .Y(n_615) );
INVx1_ASAP7_75t_L g420 ( .A(n_285), .Y(n_420) );
INVxp67_ASAP7_75t_L g472 ( .A(n_285), .Y(n_472) );
AOI21xp33_ASAP7_75t_SL g859 ( .A1(n_288), .A2(n_625), .B(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g609 ( .A(n_289), .Y(n_609) );
INVx1_ASAP7_75t_L g642 ( .A(n_290), .Y(n_642) );
INVx1_ASAP7_75t_L g559 ( .A(n_291), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_295), .A2(n_311), .B1(n_518), .B2(n_524), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g1237 ( .A1(n_297), .A2(n_329), .B1(n_585), .B2(n_897), .Y(n_1237) );
INVx2_ASAP7_75t_L g380 ( .A(n_298), .Y(n_380) );
INVx1_ASAP7_75t_L g1034 ( .A(n_306), .Y(n_1034) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_307), .A2(n_308), .B1(n_504), .B2(n_505), .Y(n_503) );
INVx1_ASAP7_75t_L g741 ( .A(n_319), .Y(n_741) );
INVx1_ASAP7_75t_L g861 ( .A(n_320), .Y(n_861) );
AOI21xp33_ASAP7_75t_L g509 ( .A1(n_323), .A2(n_510), .B(n_511), .Y(n_509) );
INVx1_ASAP7_75t_L g512 ( .A(n_324), .Y(n_512) );
INVx1_ASAP7_75t_L g889 ( .A(n_325), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_328), .A2(n_344), .B1(n_477), .B2(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g531 ( .A(n_330), .Y(n_531) );
OAI21xp5_ASAP7_75t_L g910 ( .A1(n_331), .A2(n_911), .B(n_936), .Y(n_910) );
INVx1_ASAP7_75t_L g938 ( .A(n_331), .Y(n_938) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_332), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_333), .A2(n_366), .B1(n_504), .B2(n_527), .Y(n_569) );
INVx1_ASAP7_75t_L g651 ( .A(n_336), .Y(n_651) );
XNOR2x2_ASAP7_75t_L g746 ( .A(n_338), .B(n_747), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_340), .A2(n_359), .B1(n_760), .B2(n_761), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_342), .A2(n_365), .B1(n_960), .B2(n_961), .Y(n_959) );
INVx1_ASAP7_75t_L g644 ( .A(n_347), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_349), .B(n_565), .Y(n_654) );
BUFx2_ASAP7_75t_L g867 ( .A(n_350), .Y(n_867) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_358), .A2(n_640), .B(n_641), .Y(n_639) );
AOI21xp33_ASAP7_75t_L g657 ( .A1(n_364), .A2(n_510), .B(n_658), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_367), .Y(n_764) );
AOI21xp33_ASAP7_75t_SL g485 ( .A1(n_370), .A2(n_486), .B(n_489), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_386), .B(n_975), .Y(n_375) );
INVx2_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
NAND3xp33_ASAP7_75t_L g377 ( .A(n_378), .B(n_381), .C(n_385), .Y(n_377) );
AND2x2_ASAP7_75t_L g1248 ( .A(n_378), .B(n_1249), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_378), .B(n_1250), .Y(n_1279) );
AOI21xp5_ASAP7_75t_L g1283 ( .A1(n_378), .A2(n_385), .B(n_997), .Y(n_1283) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AO21x1_ASAP7_75t_L g1281 ( .A1(n_379), .A2(n_1282), .B(n_1283), .Y(n_1281) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g984 ( .A(n_380), .B(n_985), .Y(n_984) );
AND3x4_ASAP7_75t_L g996 ( .A(n_380), .B(n_991), .C(n_997), .Y(n_996) );
NOR2xp33_ASAP7_75t_L g1249 ( .A(n_381), .B(n_1250), .Y(n_1249) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AO21x2_ASAP7_75t_L g493 ( .A1(n_382), .A2(n_494), .B(n_495), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
INVx1_ASAP7_75t_L g1250 ( .A(n_385), .Y(n_1250) );
XNOR2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_667), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
XNOR2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_575), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B1(n_528), .B2(n_574), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
XOR2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_498), .Y(n_392) );
INVx1_ASAP7_75t_L g497 ( .A(n_395), .Y(n_497) );
NAND4xp75_ASAP7_75t_L g395 ( .A(n_396), .B(n_443), .C(n_459), .D(n_479), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_427), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g758 ( .A(n_399), .Y(n_758) );
INVx1_ASAP7_75t_L g791 ( .A(n_399), .Y(n_791) );
INVx3_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
BUFx12f_ASAP7_75t_L g555 ( .A(n_400), .Y(n_555) );
BUFx6f_ASAP7_75t_L g897 ( .A(n_400), .Y(n_897) );
AND2x4_ASAP7_75t_L g400 ( .A(n_401), .B(n_412), .Y(n_400) );
AND2x2_ASAP7_75t_L g424 ( .A(n_401), .B(n_425), .Y(n_424) );
AND2x4_ASAP7_75t_L g429 ( .A(n_401), .B(n_430), .Y(n_429) );
AND2x4_ASAP7_75t_L g455 ( .A(n_401), .B(n_448), .Y(n_455) );
AND2x4_ASAP7_75t_L g504 ( .A(n_401), .B(n_452), .Y(n_504) );
AND2x4_ASAP7_75t_L g517 ( .A(n_401), .B(n_448), .Y(n_517) );
AND2x4_ASAP7_75t_L g520 ( .A(n_401), .B(n_412), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_401), .B(n_425), .Y(n_521) );
AND2x4_ASAP7_75t_L g401 ( .A(n_402), .B(n_410), .Y(n_401) );
AND2x2_ASAP7_75t_L g476 ( .A(n_402), .B(n_411), .Y(n_476) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g447 ( .A(n_403), .B(n_411), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_407), .Y(n_403) );
NAND2xp33_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
INVx2_ASAP7_75t_L g409 ( .A(n_405), .Y(n_409) );
INVx3_ASAP7_75t_L g415 ( .A(n_405), .Y(n_415) );
NAND2xp33_ASAP7_75t_L g421 ( .A(n_405), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g442 ( .A(n_405), .Y(n_442) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_405), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_406), .B(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
OAI21xp5_ASAP7_75t_L g471 ( .A1(n_408), .A2(n_442), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g470 ( .A(n_411), .B(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g462 ( .A(n_412), .B(n_447), .Y(n_462) );
AND2x4_ASAP7_75t_L g488 ( .A(n_412), .B(n_476), .Y(n_488) );
AND2x4_ASAP7_75t_L g507 ( .A(n_412), .B(n_447), .Y(n_507) );
AND2x4_ASAP7_75t_L g523 ( .A(n_412), .B(n_476), .Y(n_523) );
AND2x4_ASAP7_75t_L g412 ( .A(n_413), .B(n_417), .Y(n_412) );
INVx2_ASAP7_75t_L g426 ( .A(n_413), .Y(n_426) );
OR2x2_ASAP7_75t_L g431 ( .A(n_413), .B(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_L g448 ( .A(n_413), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g466 ( .A(n_413), .B(n_467), .Y(n_466) );
AND2x4_ASAP7_75t_L g413 ( .A(n_414), .B(n_416), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_415), .B(n_420), .Y(n_419) );
INVxp67_ASAP7_75t_L g438 ( .A(n_415), .Y(n_438) );
NAND3xp33_ASAP7_75t_L g495 ( .A(n_416), .B(n_437), .C(n_496), .Y(n_495) );
AND2x4_ASAP7_75t_L g425 ( .A(n_417), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g432 ( .A(n_418), .Y(n_432) );
AND2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_421), .Y(n_418) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
BUFx5_ASAP7_75t_L g585 ( .A(n_424), .Y(n_585) );
BUFx3_ASAP7_75t_L g706 ( .A(n_424), .Y(n_706) );
INVx1_ASAP7_75t_L g1260 ( .A(n_424), .Y(n_1260) );
AND2x4_ASAP7_75t_L g475 ( .A(n_425), .B(n_476), .Y(n_475) );
AND2x4_ASAP7_75t_L g478 ( .A(n_425), .B(n_436), .Y(n_478) );
AND2x2_ASAP7_75t_L g484 ( .A(n_425), .B(n_447), .Y(n_484) );
AND2x4_ASAP7_75t_L g505 ( .A(n_425), .B(n_436), .Y(n_505) );
AND2x2_ASAP7_75t_L g510 ( .A(n_425), .B(n_476), .Y(n_510) );
AND2x2_ASAP7_75t_L g640 ( .A(n_425), .B(n_447), .Y(n_640) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_429), .Y(n_587) );
BUFx6f_ASAP7_75t_L g699 ( .A(n_429), .Y(n_699) );
BUFx6f_ASAP7_75t_L g750 ( .A(n_429), .Y(n_750) );
AND2x4_ASAP7_75t_L g435 ( .A(n_430), .B(n_436), .Y(n_435) );
AND2x4_ASAP7_75t_L g518 ( .A(n_430), .B(n_447), .Y(n_518) );
AND2x4_ASAP7_75t_L g527 ( .A(n_430), .B(n_436), .Y(n_527) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g452 ( .A(n_431), .Y(n_452) );
INVx1_ASAP7_75t_L g449 ( .A(n_432), .Y(n_449) );
INVx3_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g547 ( .A(n_434), .Y(n_547) );
INVx1_ASAP7_75t_L g677 ( .A(n_434), .Y(n_677) );
INVx5_ASAP7_75t_L g700 ( .A(n_434), .Y(n_700) );
INVx1_ASAP7_75t_L g915 ( .A(n_434), .Y(n_915) );
INVx6_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx12f_ASAP7_75t_L g837 ( .A(n_435), .Y(n_837) );
AND2x4_ASAP7_75t_L g458 ( .A(n_436), .B(n_448), .Y(n_458) );
AND2x4_ASAP7_75t_L g526 ( .A(n_436), .B(n_448), .Y(n_526) );
AND2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_441), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_453), .Y(n_443) );
BUFx3_ASAP7_75t_L g954 ( .A(n_445), .Y(n_954) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx8_ASAP7_75t_L g760 ( .A(n_446), .Y(n_760) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
AND2x4_ASAP7_75t_L g451 ( .A(n_447), .B(n_452), .Y(n_451) );
AND2x4_ASAP7_75t_L g524 ( .A(n_447), .B(n_448), .Y(n_524) );
AND2x2_ASAP7_75t_L g550 ( .A(n_447), .B(n_448), .Y(n_550) );
BUFx3_ASAP7_75t_L g917 ( .A(n_450), .Y(n_917) );
BUFx12f_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_451), .Y(n_551) );
BUFx6f_ASAP7_75t_L g681 ( .A(n_451), .Y(n_681) );
BUFx6f_ASAP7_75t_L g702 ( .A(n_451), .Y(n_702) );
BUFx3_ASAP7_75t_L g761 ( .A(n_451), .Y(n_761) );
BUFx2_ASAP7_75t_SL g950 ( .A(n_454), .Y(n_950) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx12f_ASAP7_75t_L g704 ( .A(n_455), .Y(n_704) );
BUFx6f_ASAP7_75t_L g1239 ( .A(n_455), .Y(n_1239) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g553 ( .A(n_457), .Y(n_553) );
INVx4_ASAP7_75t_L g592 ( .A(n_457), .Y(n_592) );
INVx4_ASAP7_75t_L g755 ( .A(n_457), .Y(n_755) );
INVx1_ASAP7_75t_L g812 ( .A(n_457), .Y(n_812) );
INVx4_ASAP7_75t_L g833 ( .A(n_457), .Y(n_833) );
INVx8_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_473), .Y(n_459) );
BUFx2_ASAP7_75t_L g961 ( .A(n_461), .Y(n_961) );
BUFx3_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g597 ( .A(n_462), .Y(n_597) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_462), .Y(n_627) );
INVx4_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g535 ( .A(n_464), .Y(n_535) );
INVx3_ASAP7_75t_L g628 ( .A(n_464), .Y(n_628) );
INVx2_ASAP7_75t_L g782 ( .A(n_464), .Y(n_782) );
INVx2_ASAP7_75t_L g1274 ( .A(n_464), .Y(n_1274) );
INVx5_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx2_ASAP7_75t_L g716 ( .A(n_465), .Y(n_716) );
BUFx2_ASAP7_75t_L g800 ( .A(n_465), .Y(n_800) );
BUFx4f_ASAP7_75t_L g841 ( .A(n_465), .Y(n_841) );
AND2x4_ASAP7_75t_L g465 ( .A(n_466), .B(n_470), .Y(n_465) );
AND2x2_ASAP7_75t_L g508 ( .A(n_466), .B(n_470), .Y(n_508) );
AND2x4_ASAP7_75t_L g692 ( .A(n_466), .B(n_470), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
INVx1_ASAP7_75t_L g494 ( .A(n_468), .Y(n_494) );
BUFx3_ASAP7_75t_L g963 ( .A(n_474), .Y(n_963) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx8_ASAP7_75t_SL g638 ( .A(n_475), .Y(n_638) );
BUFx6f_ASAP7_75t_L g712 ( .A(n_475), .Y(n_712) );
BUFx3_ASAP7_75t_L g773 ( .A(n_475), .Y(n_773) );
INVx2_ASAP7_75t_L g935 ( .A(n_475), .Y(n_935) );
BUFx3_ASAP7_75t_L g776 ( .A(n_477), .Y(n_776) );
INVx3_ASAP7_75t_L g886 ( .A(n_477), .Y(n_886) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx3_ASAP7_75t_L g798 ( .A(n_478), .Y(n_798) );
BUFx6f_ASAP7_75t_L g1236 ( .A(n_478), .Y(n_1236) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_485), .Y(n_479) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g688 ( .A(n_482), .Y(n_688) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g565 ( .A(n_483), .Y(n_565) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx3_ASAP7_75t_L g502 ( .A(n_484), .Y(n_502) );
INVx3_ASAP7_75t_L g538 ( .A(n_484), .Y(n_538) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g766 ( .A(n_487), .Y(n_766) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_488), .Y(n_541) );
BUFx3_ASAP7_75t_L g625 ( .A(n_488), .Y(n_625) );
BUFx3_ASAP7_75t_L g685 ( .A(n_488), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
INVx1_ASAP7_75t_L g694 ( .A(n_491), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_491), .B(n_710), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_491), .B(n_741), .Y(n_740) );
NOR2xp33_ASAP7_75t_L g802 ( .A(n_491), .B(n_803), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_491), .B(n_820), .Y(n_819) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_492), .Y(n_544) );
INVx2_ASAP7_75t_L g927 ( .A(n_492), .Y(n_927) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx3_ASAP7_75t_L g514 ( .A(n_493), .Y(n_514) );
OA22x2_ASAP7_75t_L g556 ( .A1(n_498), .A2(n_557), .B1(n_558), .B2(n_573), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_498), .Y(n_557) );
OR2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_515), .Y(n_499) );
NAND4xp25_ASAP7_75t_L g500 ( .A(n_501), .B(n_503), .C(n_506), .D(n_509), .Y(n_500) );
BUFx3_ASAP7_75t_L g932 ( .A(n_502), .Y(n_932) );
INVx2_ASAP7_75t_L g1225 ( .A(n_502), .Y(n_1225) );
INVx2_ASAP7_75t_L g736 ( .A(n_505), .Y(n_736) );
INVx1_ASAP7_75t_L g734 ( .A(n_507), .Y(n_734) );
INVx2_ASAP7_75t_L g868 ( .A(n_507), .Y(n_868) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_510), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .Y(n_511) );
INVx1_ASAP7_75t_L g567 ( .A(n_513), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_513), .B(n_601), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_513), .B(n_609), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_513), .B(n_659), .Y(n_658) );
INVx4_ASAP7_75t_L g903 ( .A(n_513), .Y(n_903) );
NOR2xp33_ASAP7_75t_L g1226 ( .A(n_513), .B(n_1227), .Y(n_1226) );
INVx4_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx3_ASAP7_75t_L g643 ( .A(n_514), .Y(n_643) );
NAND4xp25_ASAP7_75t_L g515 ( .A(n_516), .B(n_519), .C(n_522), .D(n_525), .Y(n_515) );
INVx2_ASAP7_75t_L g731 ( .A(n_523), .Y(n_731) );
INVx1_ASAP7_75t_L g574 ( .A(n_528), .Y(n_574) );
XOR2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_556), .Y(n_528) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
XNOR2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
NOR2xp67_ASAP7_75t_L g532 ( .A(n_533), .B(n_545), .Y(n_532) );
NAND4xp25_ASAP7_75t_L g533 ( .A(n_534), .B(n_536), .C(n_539), .D(n_540), .Y(n_533) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g599 ( .A(n_538), .Y(n_599) );
INVx2_ASAP7_75t_L g606 ( .A(n_538), .Y(n_606) );
INVx2_ASAP7_75t_L g714 ( .A(n_538), .Y(n_714) );
INVx3_ASAP7_75t_SL g780 ( .A(n_538), .Y(n_780) );
INVx2_ASAP7_75t_L g968 ( .A(n_538), .Y(n_968) );
INVx4_ASAP7_75t_L g890 ( .A(n_541), .Y(n_890) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
NAND4xp25_ASAP7_75t_SL g545 ( .A(n_546), .B(n_548), .C(n_552), .D(n_554), .Y(n_545) );
BUFx4f_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
BUFx6f_ASAP7_75t_L g590 ( .A(n_550), .Y(n_590) );
BUFx2_ASAP7_75t_SL g951 ( .A(n_553), .Y(n_951) );
XNOR2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
XOR2xp5_ASAP7_75t_L g573 ( .A(n_559), .B(n_560), .Y(n_573) );
OR2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_568), .Y(n_560) );
NAND4xp25_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .C(n_564), .D(n_566), .Y(n_561) );
NAND4xp25_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .C(n_571), .D(n_572), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_648), .B1(n_649), .B2(n_665), .Y(n_575) );
OAI21xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_619), .B(n_645), .Y(n_576) );
AOI22x1_ASAP7_75t_SL g665 ( .A1(n_577), .A2(n_620), .B1(n_646), .B2(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g647 ( .A(n_578), .Y(n_647) );
AO22x2_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_580), .B1(n_603), .B2(n_618), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND4xp75_ASAP7_75t_L g582 ( .A(n_583), .B(n_588), .C(n_593), .D(n_598), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_586), .Y(n_583) );
BUFx3_ASAP7_75t_L g948 ( .A(n_585), .Y(n_948) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .Y(n_588) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
BUFx3_ASAP7_75t_L g769 ( .A(n_596), .Y(n_769) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
BUFx6f_ASAP7_75t_L g930 ( .A(n_597), .Y(n_930) );
INVx1_ASAP7_75t_L g618 ( .A(n_603), .Y(n_618) );
NAND3x1_ASAP7_75t_L g604 ( .A(n_605), .B(n_610), .C(n_613), .Y(n_604) );
HB1xp67_ASAP7_75t_L g1272 ( .A(n_606), .Y(n_1272) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
AND4x1_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .C(n_616), .D(n_617), .Y(n_613) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_621), .Y(n_646) );
XOR2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_644), .Y(n_621) );
NOR4xp75_ASAP7_75t_L g622 ( .A(n_623), .B(n_629), .C(n_632), .D(n_635), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
INVx2_ASAP7_75t_L g923 ( .A(n_625), .Y(n_923) );
INVx3_ASAP7_75t_L g884 ( .A(n_627), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_633), .B(n_634), .Y(n_632) );
OAI21x1_ASAP7_75t_SL g635 ( .A1(n_636), .A2(n_637), .B(n_639), .Y(n_635) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_640), .Y(n_739) );
INVx2_ASAP7_75t_L g818 ( .A(n_640), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
INVx4_ASAP7_75t_L g783 ( .A(n_643), .Y(n_783) );
NOR2xp33_ASAP7_75t_L g843 ( .A(n_643), .B(n_844), .Y(n_843) );
NOR2xp33_ASAP7_75t_L g860 ( .A(n_643), .B(n_861), .Y(n_860) );
NOR2xp33_ASAP7_75t_L g969 ( .A(n_643), .B(n_970), .Y(n_969) );
NOR2xp33_ASAP7_75t_L g1268 ( .A(n_643), .B(n_1269), .Y(n_1268) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
INVx2_ASAP7_75t_L g666 ( .A(n_647), .Y(n_666) );
INVx3_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
BUFx3_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
XNOR2x1_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
OR2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_660), .Y(n_652) );
NAND4xp25_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .C(n_656), .D(n_657), .Y(n_653) );
NAND4xp25_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .C(n_663), .D(n_664), .Y(n_660) );
XNOR2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_850), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_744), .B1(n_848), .B2(n_849), .Y(n_668) );
BUFx3_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g848 ( .A(n_670), .Y(n_848) );
OAI22x1_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_718), .B1(n_742), .B2(n_743), .Y(n_670) );
INVx2_ASAP7_75t_L g742 ( .A(n_671), .Y(n_742) );
OA22x2_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .B1(n_695), .B2(n_717), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NAND4xp75_ASAP7_75t_L g674 ( .A(n_675), .B(n_679), .C(n_683), .D(n_687), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .Y(n_675) );
AND2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_682), .Y(n_679) );
HB1xp67_ASAP7_75t_L g955 ( .A(n_681), .Y(n_955) );
AND2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_686), .Y(n_683) );
BUFx2_ASAP7_75t_L g960 ( .A(n_685), .Y(n_960) );
OAI21xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_691), .B(n_693), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g863 ( .A1(n_691), .A2(n_864), .B1(n_866), .B2(n_868), .Y(n_863) );
INVx4_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx2_ASAP7_75t_L g717 ( .A(n_695), .Y(n_717) );
INVx1_ASAP7_75t_SL g941 ( .A(n_695), .Y(n_941) );
NOR2x1_ASAP7_75t_L g696 ( .A(n_697), .B(n_707), .Y(n_696) );
NAND4xp25_ASAP7_75t_L g697 ( .A(n_698), .B(n_701), .C(n_703), .D(n_705), .Y(n_697) );
BUFx3_ASAP7_75t_L g914 ( .A(n_699), .Y(n_914) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_700), .Y(n_751) );
BUFx12f_ASAP7_75t_L g754 ( .A(n_704), .Y(n_754) );
NAND4xp25_ASAP7_75t_SL g707 ( .A(n_708), .B(n_711), .C(n_713), .D(n_715), .Y(n_707) );
INVx2_ASAP7_75t_L g815 ( .A(n_712), .Y(n_815) );
INVx1_ASAP7_75t_L g940 ( .A(n_717), .Y(n_940) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g743 ( .A(n_720), .Y(n_743) );
NAND4xp75_ASAP7_75t_L g721 ( .A(n_722), .B(n_725), .C(n_728), .D(n_738), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
AND2x2_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_729), .B(n_733), .Y(n_728) );
OAI21xp33_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_731), .B(n_732), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_735), .B1(n_736), .B2(n_737), .Y(n_733) );
INVx1_ASAP7_75t_L g849 ( .A(n_744), .Y(n_849) );
XNOR2x1_ASAP7_75t_SL g744 ( .A(n_745), .B(n_784), .Y(n_744) );
BUFx3_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NAND3xp33_ASAP7_75t_SL g747 ( .A(n_748), .B(n_752), .C(n_762), .Y(n_747) );
BUFx3_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
AND3x1_ASAP7_75t_L g752 ( .A(n_753), .B(n_756), .C(n_759), .Y(n_752) );
BUFx4f_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
NOR3xp33_ASAP7_75t_L g762 ( .A(n_763), .B(n_770), .C(n_777), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_765), .B1(n_767), .B2(n_768), .Y(n_763) );
INVx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVxp67_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_772), .B1(n_774), .B2(n_775), .Y(n_770) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
OAI21xp33_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_779), .B(n_781), .Y(n_777) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
AO22x2_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_827), .B1(n_846), .B2(n_847), .Y(n_784) );
INVx2_ASAP7_75t_L g847 ( .A(n_785), .Y(n_847) );
XNOR2x1_ASAP7_75t_L g785 ( .A(n_786), .B(n_807), .Y(n_785) );
OAI22x1_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_794), .B1(n_805), .B2(n_806), .Y(n_786) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_788), .B(n_795), .Y(n_805) );
NAND4xp25_ASAP7_75t_L g788 ( .A(n_789), .B(n_790), .C(n_792), .D(n_793), .Y(n_788) );
NAND4xp25_ASAP7_75t_L g795 ( .A(n_796), .B(n_799), .C(n_801), .D(n_804), .Y(n_795) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g964 ( .A(n_798), .Y(n_964) );
NAND4xp75_ASAP7_75t_L g808 ( .A(n_809), .B(n_813), .C(n_821), .D(n_824), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .Y(n_809) );
OA21x2_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_815), .B(n_816), .Y(n_813) );
INVx2_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
AND2x2_ASAP7_75t_L g821 ( .A(n_822), .B(n_823), .Y(n_821) );
AND2x2_ASAP7_75t_L g824 ( .A(n_825), .B(n_826), .Y(n_824) );
BUFx3_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g846 ( .A(n_828), .Y(n_846) );
XNOR2x1_ASAP7_75t_L g828 ( .A(n_829), .B(n_845), .Y(n_828) );
NAND4xp75_ASAP7_75t_L g829 ( .A(n_830), .B(n_834), .C(n_838), .D(n_842), .Y(n_829) );
AND2x2_ASAP7_75t_L g830 ( .A(n_831), .B(n_832), .Y(n_830) );
AND2x2_ASAP7_75t_L g834 ( .A(n_835), .B(n_836), .Y(n_834) );
BUFx3_ASAP7_75t_L g957 ( .A(n_837), .Y(n_957) );
AND2x2_ASAP7_75t_L g838 ( .A(n_839), .B(n_840), .Y(n_838) );
XNOR2xp5_ASAP7_75t_L g850 ( .A(n_851), .B(n_904), .Y(n_850) );
AO22x1_ASAP7_75t_L g851 ( .A1(n_852), .A2(n_853), .B1(n_877), .B2(n_878), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g876 ( .A(n_857), .Y(n_876) );
NOR2x1_ASAP7_75t_L g857 ( .A(n_858), .B(n_870), .Y(n_857) );
NAND3xp33_ASAP7_75t_L g858 ( .A(n_859), .B(n_862), .C(n_869), .Y(n_858) );
CKINVDCx16_ASAP7_75t_R g864 ( .A(n_865), .Y(n_864) );
CKINVDCx9p33_ASAP7_75t_R g866 ( .A(n_867), .Y(n_866) );
NAND4xp25_ASAP7_75t_L g870 ( .A(n_871), .B(n_872), .C(n_873), .D(n_874), .Y(n_870) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx2_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
NAND4xp75_ASAP7_75t_L g881 ( .A(n_882), .B(n_892), .C(n_895), .D(n_899), .Y(n_881) );
NOR2xp67_ASAP7_75t_L g882 ( .A(n_883), .B(n_888), .Y(n_882) );
OAI22xp5_ASAP7_75t_L g883 ( .A1(n_884), .A2(n_885), .B1(n_886), .B2(n_887), .Y(n_883) );
OAI21xp5_ASAP7_75t_L g888 ( .A1(n_889), .A2(n_890), .B(n_891), .Y(n_888) );
AND2x2_ASAP7_75t_L g892 ( .A(n_893), .B(n_894), .Y(n_892) );
AND2x2_ASAP7_75t_L g895 ( .A(n_896), .B(n_898), .Y(n_895) );
NOR2xp33_ASAP7_75t_L g900 ( .A(n_901), .B(n_902), .Y(n_900) );
INVx2_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
AOI22x1_ASAP7_75t_L g904 ( .A1(n_905), .A2(n_942), .B1(n_971), .B2(n_973), .Y(n_904) );
INVx2_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
INVx2_ASAP7_75t_SL g907 ( .A(n_908), .Y(n_907) );
INVx1_ASAP7_75t_L g972 ( .A(n_908), .Y(n_972) );
OA22x2_ASAP7_75t_L g908 ( .A1(n_909), .A2(n_910), .B1(n_940), .B2(n_941), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
NOR2xp33_ASAP7_75t_L g911 ( .A(n_912), .B(n_920), .Y(n_911) );
INVxp67_ASAP7_75t_L g939 ( .A(n_912), .Y(n_939) );
NAND4xp25_ASAP7_75t_L g912 ( .A(n_913), .B(n_916), .C(n_918), .D(n_919), .Y(n_912) );
NOR2xp33_ASAP7_75t_L g937 ( .A(n_920), .B(n_938), .Y(n_937) );
NAND4xp25_ASAP7_75t_L g920 ( .A(n_921), .B(n_928), .C(n_931), .D(n_933), .Y(n_920) );
INVx2_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
NOR2xp33_ASAP7_75t_L g924 ( .A(n_925), .B(n_926), .Y(n_924) );
INVx3_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
INVx2_ASAP7_75t_L g1275 ( .A(n_930), .Y(n_1275) );
INVx3_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_937), .B(n_939), .Y(n_936) );
OAI22xp5_ASAP7_75t_L g1035 ( .A1(n_938), .A2(n_1036), .B1(n_1038), .B2(n_1039), .Y(n_1035) );
INVx1_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
BUFx3_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
INVx2_ASAP7_75t_SL g974 ( .A(n_944), .Y(n_974) );
NAND4xp75_ASAP7_75t_L g945 ( .A(n_946), .B(n_952), .C(n_958), .D(n_965), .Y(n_945) );
AND2x2_ASAP7_75t_L g946 ( .A(n_947), .B(n_949), .Y(n_946) );
AND2x2_ASAP7_75t_L g952 ( .A(n_953), .B(n_956), .Y(n_952) );
AND2x2_ASAP7_75t_L g958 ( .A(n_959), .B(n_962), .Y(n_958) );
INVx1_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
INVx2_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
INVx1_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
OAI221xp5_ASAP7_75t_L g975 ( .A1(n_976), .A2(n_1216), .B1(n_1219), .B2(n_1247), .C(n_1251), .Y(n_975) );
AOI211xp5_ASAP7_75t_L g976 ( .A1(n_977), .A2(n_1115), .B(n_1120), .C(n_1188), .Y(n_976) );
NAND4xp25_ASAP7_75t_L g977 ( .A(n_978), .B(n_1060), .C(n_1083), .D(n_1104), .Y(n_977) );
AOI211xp5_ASAP7_75t_L g978 ( .A1(n_979), .A2(n_1002), .B(n_1022), .C(n_1047), .Y(n_978) );
AOI21xp33_ASAP7_75t_L g1157 ( .A1(n_979), .A2(n_1158), .B(n_1159), .Y(n_1157) );
INVx1_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
NOR2xp33_ASAP7_75t_L g1079 ( .A(n_980), .B(n_1059), .Y(n_1079) );
OR2x2_ASAP7_75t_L g980 ( .A(n_981), .B(n_994), .Y(n_980) );
INVx1_ASAP7_75t_L g1042 ( .A(n_981), .Y(n_1042) );
INVx1_ASAP7_75t_L g1050 ( .A(n_981), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_982), .B(n_989), .Y(n_981) );
AND2x2_ASAP7_75t_L g983 ( .A(n_984), .B(n_986), .Y(n_983) );
AND2x4_ASAP7_75t_L g990 ( .A(n_984), .B(n_991), .Y(n_990) );
AND2x2_ASAP7_75t_L g1000 ( .A(n_984), .B(n_986), .Y(n_1000) );
AND2x4_ASAP7_75t_L g1037 ( .A(n_984), .B(n_986), .Y(n_1037) );
AND2x2_ASAP7_75t_L g987 ( .A(n_986), .B(n_988), .Y(n_987) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_986), .B(n_988), .Y(n_1001) );
AND2x4_ASAP7_75t_L g1006 ( .A(n_986), .B(n_988), .Y(n_1006) );
AND2x4_ASAP7_75t_L g993 ( .A(n_988), .B(n_991), .Y(n_993) );
AND2x4_ASAP7_75t_L g998 ( .A(n_988), .B(n_991), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g1033 ( .A(n_988), .B(n_991), .Y(n_1033) );
INVx3_ASAP7_75t_L g1031 ( .A(n_990), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_994), .B(n_1041), .Y(n_1040) );
OR2x2_ASAP7_75t_L g1043 ( .A(n_994), .B(n_1029), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_994), .B(n_1059), .Y(n_1058) );
INVx2_ASAP7_75t_L g1075 ( .A(n_994), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_994), .B(n_1042), .Y(n_1082) );
OR2x2_ASAP7_75t_L g1087 ( .A(n_994), .B(n_1059), .Y(n_1087) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_994), .B(n_1029), .Y(n_1100) );
OR2x2_ASAP7_75t_L g1113 ( .A(n_994), .B(n_1042), .Y(n_1113) );
HB1xp67_ASAP7_75t_L g1135 ( .A(n_994), .Y(n_1135) );
AND2x2_ASAP7_75t_L g994 ( .A(n_995), .B(n_999), .Y(n_994) );
NOR2x1_ASAP7_75t_R g1002 ( .A(n_1003), .B(n_1008), .Y(n_1002) );
NAND2xp5_ASAP7_75t_L g1025 ( .A(n_1003), .B(n_1012), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_1003), .B(n_1046), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_1003), .B(n_1053), .Y(n_1077) );
NOR2xp33_ASAP7_75t_L g1092 ( .A(n_1003), .B(n_1093), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g1132 ( .A(n_1003), .B(n_1015), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1003), .B(n_1091), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1003), .B(n_1011), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1003), .B(n_1158), .Y(n_1193) );
INVx1_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
INVx1_ASAP7_75t_SL g1056 ( .A(n_1004), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1090 ( .A(n_1004), .B(n_1091), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g1125 ( .A(n_1004), .B(n_1126), .Y(n_1125) );
OR2x2_ASAP7_75t_L g1140 ( .A(n_1004), .B(n_1065), .Y(n_1140) );
NAND2xp5_ASAP7_75t_L g1172 ( .A(n_1004), .B(n_1012), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1004), .B(n_1158), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1007), .Y(n_1004) );
INVx2_ASAP7_75t_L g1038 ( .A(n_1006), .Y(n_1038) );
NAND2xp5_ASAP7_75t_SL g1008 ( .A(n_1009), .B(n_1018), .Y(n_1008) );
INVx3_ASAP7_75t_SL g1009 ( .A(n_1010), .Y(n_1009) );
NOR2x1_ASAP7_75t_L g1158 ( .A(n_1010), .B(n_1018), .Y(n_1158) );
OR2x2_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1015), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1053 ( .A(n_1011), .B(n_1015), .Y(n_1053) );
INVx1_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_1012), .B(n_1015), .Y(n_1046) );
OR2x2_ASAP7_75t_L g1065 ( .A(n_1012), .B(n_1015), .Y(n_1065) );
AOI221xp5_ASAP7_75t_L g1178 ( .A1(n_1012), .A2(n_1027), .B1(n_1108), .B2(n_1179), .C(n_1181), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_1013), .B(n_1014), .Y(n_1012) );
O2A1O1Ixp33_ASAP7_75t_L g1047 ( .A1(n_1015), .A2(n_1048), .B(n_1051), .C(n_1057), .Y(n_1047) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1015), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1015), .B(n_1055), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1015 ( .A(n_1016), .B(n_1017), .Y(n_1015) );
NAND2xp5_ASAP7_75t_SL g1023 ( .A(n_1018), .B(n_1024), .Y(n_1023) );
NOR2xp33_ASAP7_75t_L g1049 ( .A(n_1018), .B(n_1050), .Y(n_1049) );
INVx2_ASAP7_75t_L g1062 ( .A(n_1018), .Y(n_1062) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1018), .Y(n_1096) );
INVx2_ASAP7_75t_L g1099 ( .A(n_1018), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1018), .B(n_1053), .Y(n_1126) );
BUFx6f_ASAP7_75t_L g1138 ( .A(n_1018), .Y(n_1138) );
NAND2xp5_ASAP7_75t_L g1161 ( .A(n_1018), .B(n_1162), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1018), .B(n_1028), .Y(n_1173) );
INVx4_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
OR2x2_ASAP7_75t_L g1054 ( .A(n_1019), .B(n_1055), .Y(n_1054) );
NAND2xp5_ASAP7_75t_L g1130 ( .A(n_1019), .B(n_1059), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1019), .B(n_1029), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_1020), .B(n_1021), .Y(n_1019) );
OAI22xp5_ASAP7_75t_L g1022 ( .A1(n_1023), .A2(n_1026), .B1(n_1043), .B2(n_1044), .Y(n_1022) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
NAND2xp5_ASAP7_75t_L g1026 ( .A(n_1027), .B(n_1040), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_1027), .B(n_1071), .Y(n_1070) );
INVx2_ASAP7_75t_L g1027 ( .A(n_1028), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g1101 ( .A(n_1028), .B(n_1085), .Y(n_1101) );
NAND2xp5_ASAP7_75t_L g1201 ( .A(n_1028), .B(n_1061), .Y(n_1201) );
INVx1_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
INVx2_ASAP7_75t_L g1059 ( .A(n_1029), .Y(n_1059) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_1029), .B(n_1082), .Y(n_1081) );
OR2x2_ASAP7_75t_L g1029 ( .A(n_1030), .B(n_1035), .Y(n_1029) );
OAI22xp5_ASAP7_75t_L g1030 ( .A1(n_1031), .A2(n_1032), .B1(n_1033), .B2(n_1034), .Y(n_1030) );
OAI221xp5_ASAP7_75t_L g1116 ( .A1(n_1031), .A2(n_1033), .B1(n_1117), .B2(n_1118), .C(n_1119), .Y(n_1116) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1031), .Y(n_1218) );
INVx3_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
AOI221xp5_ASAP7_75t_L g1143 ( .A1(n_1040), .A2(n_1144), .B1(n_1146), .B2(n_1149), .C(n_1156), .Y(n_1143) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1041), .Y(n_1071) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
NOR2xp33_ASAP7_75t_L g1095 ( .A(n_1043), .B(n_1096), .Y(n_1095) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1043), .Y(n_1148) );
NOR2xp33_ASAP7_75t_L g1164 ( .A(n_1043), .B(n_1050), .Y(n_1164) );
OAI22xp5_ASAP7_75t_L g1206 ( .A1(n_1043), .A2(n_1207), .B1(n_1208), .B2(n_1210), .Y(n_1206) );
OAI221xp5_ASAP7_75t_L g1156 ( .A1(n_1044), .A2(n_1115), .B1(n_1157), .B2(n_1163), .C(n_1165), .Y(n_1156) );
INVx1_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1045), .B(n_1058), .Y(n_1142) );
NAND2xp5_ASAP7_75t_L g1067 ( .A(n_1046), .B(n_1068), .Y(n_1067) );
NAND2xp5_ASAP7_75t_L g1080 ( .A(n_1046), .B(n_1081), .Y(n_1080) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1046), .Y(n_1094) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_1046), .B(n_1055), .Y(n_1103) );
INVx1_ASAP7_75t_L g1048 ( .A(n_1049), .Y(n_1048) );
INVx2_ASAP7_75t_L g1085 ( .A(n_1050), .Y(n_1085) );
BUFx3_ASAP7_75t_L g1147 ( .A(n_1050), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1050), .B(n_1059), .Y(n_1176) );
OR2x2_ASAP7_75t_L g1051 ( .A(n_1052), .B(n_1054), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1053), .B(n_1055), .Y(n_1108) );
INVx1_ASAP7_75t_L g1068 ( .A(n_1054), .Y(n_1068) );
AND2x4_ASAP7_75t_L g1063 ( .A(n_1055), .B(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
INVx2_ASAP7_75t_L g1106 ( .A(n_1059), .Y(n_1106) );
AOI21xp33_ASAP7_75t_SL g1192 ( .A1(n_1059), .A2(n_1193), .B(n_1194), .Y(n_1192) );
O2A1O1Ixp33_ASAP7_75t_L g1060 ( .A1(n_1061), .A2(n_1066), .B(n_1069), .C(n_1072), .Y(n_1060) );
AND2x2_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1063), .Y(n_1061) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1062), .Y(n_1074) );
NAND2xp5_ASAP7_75t_L g1089 ( .A(n_1062), .B(n_1090), .Y(n_1089) );
NAND2xp5_ASAP7_75t_L g1111 ( .A(n_1062), .B(n_1077), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_1062), .B(n_1155), .Y(n_1154) );
NOR2xp33_ASAP7_75t_L g1214 ( .A(n_1062), .B(n_1065), .Y(n_1214) );
NAND2xp5_ASAP7_75t_L g1073 ( .A(n_1063), .B(n_1074), .Y(n_1073) );
INVx2_ASAP7_75t_SL g1152 ( .A(n_1063), .Y(n_1152) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_1065), .B(n_1094), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g1186 ( .A1(n_1066), .A2(n_1082), .B1(n_1169), .B2(n_1187), .Y(n_1186) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
INVx1_ASAP7_75t_L g1069 ( .A(n_1070), .Y(n_1069) );
NOR2xp33_ASAP7_75t_L g1184 ( .A(n_1071), .B(n_1132), .Y(n_1184) );
OAI221xp5_ASAP7_75t_L g1072 ( .A1(n_1073), .A2(n_1075), .B1(n_1076), .B2(n_1078), .C(n_1080), .Y(n_1072) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_1074), .B(n_1103), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1075), .B(n_1180), .Y(n_1179) );
CKINVDCx14_ASAP7_75t_R g1205 ( .A(n_1075), .Y(n_1205) );
NAND2xp5_ASAP7_75t_L g1208 ( .A(n_1075), .B(n_1209), .Y(n_1208) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1077), .Y(n_1076) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1081), .Y(n_1215) );
AOI211xp5_ASAP7_75t_L g1104 ( .A1(n_1082), .A2(n_1105), .B(n_1109), .C(n_1112), .Y(n_1104) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1082), .Y(n_1160) );
AOI221xp5_ASAP7_75t_L g1083 ( .A1(n_1084), .A2(n_1088), .B1(n_1092), .B2(n_1095), .C(n_1097), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_1085), .B(n_1086), .Y(n_1084) );
NOR2xp33_ASAP7_75t_L g1174 ( .A(n_1085), .B(n_1115), .Y(n_1174) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1085), .Y(n_1194) );
NAND2xp5_ASAP7_75t_L g1195 ( .A(n_1085), .B(n_1116), .Y(n_1195) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
NOR2xp33_ASAP7_75t_L g1199 ( .A(n_1087), .B(n_1096), .Y(n_1199) );
INVxp67_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_1091), .B(n_1138), .Y(n_1145) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1095), .Y(n_1185) );
AOI21xp5_ASAP7_75t_L g1097 ( .A1(n_1098), .A2(n_1101), .B(n_1102), .Y(n_1097) );
NAND2xp5_ASAP7_75t_L g1098 ( .A(n_1099), .B(n_1100), .Y(n_1098) );
NAND2xp67_ASAP7_75t_L g1107 ( .A(n_1099), .B(n_1108), .Y(n_1107) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1100), .Y(n_1139) );
AOI221xp5_ASAP7_75t_SL g1175 ( .A1(n_1100), .A2(n_1124), .B1(n_1154), .B2(n_1176), .C(n_1177), .Y(n_1175) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1101), .Y(n_1187) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1103), .Y(n_1102) );
NOR2xp33_ASAP7_75t_L g1207 ( .A(n_1103), .B(n_1155), .Y(n_1207) );
NOR2xp67_ASAP7_75t_SL g1105 ( .A(n_1106), .B(n_1107), .Y(n_1105) );
INVx2_ASAP7_75t_L g1110 ( .A(n_1106), .Y(n_1110) );
NOR2xp33_ASAP7_75t_L g1151 ( .A(n_1106), .B(n_1152), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g1153 ( .A(n_1106), .B(n_1154), .Y(n_1153) );
AOI221xp5_ASAP7_75t_L g1196 ( .A1(n_1106), .A2(n_1172), .B1(n_1197), .B2(n_1199), .C(n_1200), .Y(n_1196) );
NOR2xp33_ASAP7_75t_L g1203 ( .A(n_1107), .B(n_1110), .Y(n_1203) );
NOR2xp33_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1111), .Y(n_1109) );
NAND2xp5_ASAP7_75t_L g1190 ( .A(n_1110), .B(n_1191), .Y(n_1190) );
AOI21xp33_ASAP7_75t_L g1212 ( .A1(n_1111), .A2(n_1213), .B(n_1215), .Y(n_1212) );
NOR2xp33_ASAP7_75t_L g1112 ( .A(n_1113), .B(n_1114), .Y(n_1112) );
OAI211xp5_ASAP7_75t_L g1144 ( .A1(n_1115), .A2(n_1125), .B(n_1140), .C(n_1145), .Y(n_1144) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1115), .Y(n_1209) );
INVx2_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
HB1xp67_ASAP7_75t_L g1122 ( .A(n_1116), .Y(n_1122) );
OAI211xp5_ASAP7_75t_L g1120 ( .A1(n_1121), .A2(n_1123), .B(n_1143), .C(n_1175), .Y(n_1120) );
INVx2_ASAP7_75t_L g1121 ( .A(n_1122), .Y(n_1121) );
O2A1O1Ixp33_ASAP7_75t_L g1123 ( .A1(n_1124), .A2(n_1127), .B(n_1133), .C(n_1136), .Y(n_1123) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
NAND3xp33_ASAP7_75t_L g1149 ( .A(n_1125), .B(n_1150), .C(n_1153), .Y(n_1149) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1126), .Y(n_1198) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_1129), .B(n_1131), .Y(n_1128) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1130), .Y(n_1129) );
NOR2xp33_ASAP7_75t_L g1166 ( .A(n_1130), .B(n_1167), .Y(n_1166) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1134), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
A2O1A1Ixp33_ASAP7_75t_L g1136 ( .A1(n_1137), .A2(n_1139), .B(n_1140), .C(n_1141), .Y(n_1136) );
AOI221xp5_ASAP7_75t_L g1202 ( .A1(n_1137), .A2(n_1203), .B1(n_1204), .B2(n_1206), .C(n_1212), .Y(n_1202) );
INVx2_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1140), .Y(n_1155) );
NAND2xp5_ASAP7_75t_L g1197 ( .A(n_1140), .B(n_1198), .Y(n_1197) );
CKINVDCx5p33_ASAP7_75t_R g1141 ( .A(n_1142), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_1147), .B(n_1148), .Y(n_1146) );
OAI321xp33_ASAP7_75t_L g1188 ( .A1(n_1148), .A2(n_1189), .A3(n_1192), .B1(n_1195), .B2(n_1196), .C(n_1202), .Y(n_1188) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
NOR2xp33_ASAP7_75t_L g1159 ( .A(n_1160), .B(n_1161), .Y(n_1159) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
OAI21xp33_ASAP7_75t_L g1165 ( .A1(n_1166), .A2(n_1169), .B(n_1174), .Y(n_1165) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1171), .B(n_1173), .Y(n_1170) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1172), .Y(n_1171) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1174), .Y(n_1182) );
OAI221xp5_ASAP7_75t_L g1177 ( .A1(n_1178), .A2(n_1182), .B1(n_1183), .B2(n_1185), .C(n_1186), .Y(n_1177) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1181), .Y(n_1191) );
INVxp67_ASAP7_75t_L g1183 ( .A(n_1184), .Y(n_1183) );
INVxp67_ASAP7_75t_SL g1189 ( .A(n_1190), .Y(n_1189) );
INVxp67_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
CKINVDCx14_ASAP7_75t_R g1204 ( .A(n_1205), .Y(n_1204) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
CKINVDCx5p33_ASAP7_75t_R g1216 ( .A(n_1217), .Y(n_1216) );
HB1xp67_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
AND2x4_ASAP7_75t_L g1219 ( .A(n_1220), .B(n_1240), .Y(n_1219) );
AOI21x1_ASAP7_75t_L g1220 ( .A1(n_1221), .A2(n_1222), .B(n_1232), .Y(n_1220) );
NAND2xp5_ASAP7_75t_L g1222 ( .A(n_1223), .B(n_1228), .Y(n_1222) );
BUFx2_ASAP7_75t_L g1241 ( .A(n_1223), .Y(n_1241) );
INVx2_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
NOR2xp33_ASAP7_75t_L g1228 ( .A(n_1229), .B(n_1231), .Y(n_1228) );
INVxp67_ASAP7_75t_SL g1229 ( .A(n_1230), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_1230), .B(n_1237), .Y(n_1245) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1231), .Y(n_1246) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1233), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1234), .B(n_1235), .Y(n_1233) );
NAND4xp75_ASAP7_75t_L g1240 ( .A(n_1241), .B(n_1242), .C(n_1245), .D(n_1246), .Y(n_1240) );
NOR2x1_ASAP7_75t_L g1242 ( .A(n_1243), .B(n_1244), .Y(n_1242) );
CKINVDCx16_ASAP7_75t_R g1247 ( .A(n_1248), .Y(n_1247) );
INVxp33_ASAP7_75t_L g1252 ( .A(n_1253), .Y(n_1252) );
INVx1_ASAP7_75t_SL g1277 ( .A(n_1254), .Y(n_1277) );
HB1xp67_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
NOR2x1_ASAP7_75t_L g1255 ( .A(n_1256), .B(n_1264), .Y(n_1255) );
NAND4xp25_ASAP7_75t_L g1256 ( .A(n_1257), .B(n_1261), .C(n_1262), .D(n_1263), .Y(n_1256) );
BUFx6f_ASAP7_75t_L g1258 ( .A(n_1259), .Y(n_1258) );
INVx2_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
NAND3xp33_ASAP7_75t_L g1264 ( .A(n_1265), .B(n_1271), .C(n_1273), .Y(n_1264) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_1267), .B(n_1270), .Y(n_1266) );
BUFx2_ASAP7_75t_SL g1278 ( .A(n_1279), .Y(n_1278) );
HB1xp67_ASAP7_75t_L g1280 ( .A(n_1281), .Y(n_1280) );
endmodule