module fake_ibex_295_n_1871 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_193, n_108, n_350, n_165, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_371, n_357, n_88, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_244, n_73, n_343, n_310, n_323, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_370, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_22, n_136, n_261, n_30, n_367, n_221, n_355, n_102, n_52, n_99, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_141, n_222, n_186, n_349, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_335, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_75, n_137, n_338, n_173, n_363, n_180, n_369, n_201, n_14, n_351, n_368, n_257, n_77, n_44, n_66, n_305, n_307, n_192, n_140, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_26, n_188, n_200, n_199, n_308, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_381, n_382, n_95, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_342, n_233, n_385, n_118, n_378, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_345, n_119, n_361, n_72, n_319, n_195, n_212, n_311, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_344, n_393, n_297, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_399, n_254, n_213, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_1871);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_350;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_371;
input n_357;
input n_88;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_244;
input n_73;
input n_343;
input n_310;
input n_323;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_370;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_367;
input n_221;
input n_355;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_349;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_335;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_338;
input n_173;
input n_363;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_257;
input n_77;
input n_44;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_26;
input n_188;
input n_200;
input n_199;
input n_308;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_381;
input n_382;
input n_95;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_118;
input n_378;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_345;
input n_119;
input n_361;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_344;
input n_393;
input n_297;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_399;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;

output n_1871;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_1582;
wire n_766;
wire n_1110;
wire n_1382;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_1594;
wire n_1802;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_1125;
wire n_733;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_1766;
wire n_550;
wire n_557;
wire n_641;
wire n_893;
wire n_527;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_1081;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_1778;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_420;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_666;
wire n_1638;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_793;
wire n_937;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1863;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_553;
wire n_554;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_745;
wire n_447;
wire n_1753;
wire n_564;
wire n_562;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_579;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_422;
wire n_1717;
wire n_1609;
wire n_1613;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_1742;
wire n_1818;
wire n_870;
wire n_1709;
wire n_1610;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_455;
wire n_1701;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_737;
wire n_606;
wire n_1571;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_435;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_1786;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1031;
wire n_981;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_974;
wire n_1036;
wire n_1831;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_846;
wire n_471;
wire n_1793;
wire n_1237;
wire n_859;
wire n_1109;
wire n_965;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_1032;
wire n_936;
wire n_469;
wire n_1825;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_1792;
wire n_1712;
wire n_590;
wire n_1568;
wire n_1184;
wire n_1477;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_1751;
wire n_669;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_1776;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_488;
wire n_705;
wire n_1548;
wire n_429;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_1704;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_1545;
wire n_456;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_1470;
wire n_444;
wire n_1761;
wire n_1836;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_411;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1615;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_650;
wire n_409;
wire n_1575;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_951;
wire n_468;
wire n_1580;
wire n_1574;
wire n_780;
wire n_502;
wire n_1705;
wire n_633;
wire n_1746;
wire n_726;
wire n_532;
wire n_1439;
wire n_863;
wire n_597;
wire n_1832;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_1785;
wire n_486;
wire n_1870;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_1683;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1845;
wire n_1104;
wire n_1667;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1679;
wire n_1497;
wire n_1578;
wire n_1143;
wire n_1783;
wire n_418;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_1857;
wire n_545;
wire n_887;
wire n_1162;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_1323;
wire n_578;
wire n_1739;
wire n_432;
wire n_1777;
wire n_403;
wire n_1353;
wire n_423;
wire n_1429;
wire n_1546;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1834;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_1830;
wire n_1629;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_1340;
wire n_1626;
wire n_674;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_400;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_404;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1517;
wire n_690;
wire n_1225;
wire n_982;
wire n_1624;
wire n_785;
wire n_604;
wire n_1598;
wire n_977;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_1625;
wire n_933;
wire n_1774;
wire n_1797;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_1538;
wire n_487;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_1725;
wire n_1135;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_1066;
wire n_1169;
wire n_648;
wire n_571;
wire n_1726;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1337;
wire n_1647;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_480;
wire n_1057;
wire n_1473;
wire n_516;
wire n_1403;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_1718;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1740;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_1788;
wire n_786;
wire n_505;
wire n_1621;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1570;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1769;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_1632;
wire n_688;
wire n_1542;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1547;
wire n_1097;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1199;
wire n_1767;
wire n_1768;
wire n_1443;
wire n_478;
wire n_1585;
wire n_1861;
wire n_1564;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_828;
wire n_1438;
wire n_753;
wire n_747;
wire n_645;
wire n_1147;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1518;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_1693;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_1686;
wire n_1302;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_854;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1734;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_1720;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1866;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_1692;
wire n_438;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_1868;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1757;
wire n_699;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1414;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_405;
wire n_1807;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1611;
wire n_955;
wire n_440;
wire n_1333;
wire n_414;
wire n_952;
wire n_1675;
wire n_1640;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1732;
wire n_1354;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_1843;
wire n_408;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_227),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_327),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_148),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_164),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_351),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_305),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_325),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g407 ( 
.A(n_127),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_60),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_64),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_320),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_103),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_4),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_380),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_304),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_319),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_93),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_76),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_357),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_338),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_349),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_260),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_375),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_388),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_359),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_376),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_326),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_124),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_381),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_268),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_364),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_225),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_24),
.Y(n_432)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_121),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_35),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_132),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_154),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_293),
.Y(n_437)
);

INVxp67_ASAP7_75t_SL g438 ( 
.A(n_130),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_204),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_39),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_362),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_322),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_255),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_384),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_78),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_29),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_218),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_342),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_149),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_339),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_311),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_296),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_54),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_222),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_12),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_192),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_262),
.Y(n_457)
);

BUFx10_ASAP7_75t_L g458 ( 
.A(n_298),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_63),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_53),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_280),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g462 ( 
.A(n_119),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_117),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_101),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_22),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_323),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_286),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_167),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_119),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_52),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_336),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_354),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_316),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_229),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_122),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_66),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_294),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_13),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_301),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_265),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_281),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_105),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_217),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_383),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_254),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_313),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_374),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_162),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_348),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_247),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_300),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_299),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_355),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_175),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_208),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_122),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_248),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_360),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_83),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_346),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_372),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_2),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_363),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_219),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_23),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_22),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_66),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_312),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_114),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_353),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_302),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_37),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_205),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_373),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_214),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_361),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_161),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_15),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_345),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_91),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_366),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_76),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_26),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_173),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_287),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_259),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_234),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_99),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_272),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_379),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_308),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_297),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_393),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_170),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_65),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_110),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_133),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_250),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_91),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_371),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_87),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_182),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_288),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_256),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_88),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_159),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_352),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_340),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_310),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_228),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_231),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_278),
.Y(n_552)
);

BUFx5_ASAP7_75t_L g553 ( 
.A(n_165),
.Y(n_553)
);

INVx1_ASAP7_75t_SL g554 ( 
.A(n_94),
.Y(n_554)
);

BUFx8_ASAP7_75t_SL g555 ( 
.A(n_290),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_377),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_292),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_369),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_230),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_382),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_321),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_270),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_395),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_39),
.Y(n_564)
);

CKINVDCx16_ASAP7_75t_R g565 ( 
.A(n_368),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_120),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_68),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_176),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_64),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_151),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_221),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_387),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_391),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_25),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_291),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_385),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_238),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_334),
.Y(n_578)
);

INVx1_ASAP7_75t_SL g579 ( 
.A(n_118),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_126),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_51),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_370),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_58),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_275),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_244),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_146),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_125),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_67),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_187),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_18),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_137),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_390),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_224),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_174),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_367),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_179),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_335),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_95),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_156),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_226),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_246),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_50),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_309),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_32),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_32),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_27),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_77),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_45),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_48),
.Y(n_609)
);

CKINVDCx16_ASAP7_75t_R g610 ( 
.A(n_141),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_274),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_3),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_166),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_249),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_48),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_317),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_33),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_181),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_303),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_329),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_108),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_328),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_350),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_5),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_33),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_223),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_13),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_356),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_20),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_314),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_344),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_386),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_365),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_79),
.Y(n_634)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_389),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_178),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_258),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_53),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_341),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_81),
.Y(n_640)
);

INVx1_ASAP7_75t_SL g641 ( 
.A(n_315),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_54),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_93),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_307),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_82),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_347),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_295),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_100),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_18),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_343),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_136),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_215),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_318),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_306),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_97),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_139),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_358),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_378),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_324),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_269),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g661 ( 
.A(n_459),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_555),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_557),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_553),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_598),
.B(n_0),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_407),
.B(n_0),
.Y(n_666)
);

INVx1_ASAP7_75t_SL g667 ( 
.A(n_555),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_589),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g669 ( 
.A(n_408),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g670 ( 
.A(n_460),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_414),
.Y(n_671)
);

INVxp33_ASAP7_75t_L g672 ( 
.A(n_605),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_408),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_496),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_578),
.B(n_1),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_605),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_609),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_520),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_449),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_609),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_456),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_638),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_638),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_457),
.Y(n_684)
);

CKINVDCx20_ASAP7_75t_R g685 ( 
.A(n_574),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_440),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_468),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_474),
.Y(n_688)
);

INVxp67_ASAP7_75t_L g689 ( 
.A(n_409),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_463),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_465),
.Y(n_691)
);

NOR2xp67_ASAP7_75t_L g692 ( 
.A(n_416),
.B(n_1),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_480),
.Y(n_693)
);

CKINVDCx20_ASAP7_75t_R g694 ( 
.A(n_583),
.Y(n_694)
);

HB1xp67_ASAP7_75t_L g695 ( 
.A(n_412),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_481),
.Y(n_696)
);

INVxp67_ASAP7_75t_SL g697 ( 
.A(n_470),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_475),
.Y(n_698)
);

CKINVDCx20_ASAP7_75t_R g699 ( 
.A(n_627),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_482),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_458),
.B(n_2),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_405),
.B(n_3),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_525),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_497),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_506),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_518),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_600),
.Y(n_707)
);

HB1xp67_ASAP7_75t_L g708 ( 
.A(n_417),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_410),
.B(n_4),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_523),
.Y(n_710)
);

BUFx2_ASAP7_75t_L g711 ( 
.A(n_432),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_603),
.Y(n_712)
);

CKINVDCx14_ASAP7_75t_R g713 ( 
.A(n_458),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_626),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_528),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_628),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_539),
.B(n_5),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_565),
.Y(n_718)
);

INVxp67_ASAP7_75t_SL g719 ( 
.A(n_545),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_564),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_610),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_413),
.B(n_6),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_424),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_571),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_567),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_612),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_571),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_621),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_572),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_624),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_648),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_572),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_649),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_655),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_458),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_423),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_657),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_427),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_553),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_430),
.Y(n_740)
);

INVxp33_ASAP7_75t_L g741 ( 
.A(n_615),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_436),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_439),
.Y(n_743)
);

INVxp67_ASAP7_75t_L g744 ( 
.A(n_433),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_686),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_662),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_671),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_703),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_713),
.B(n_434),
.Y(n_749)
);

BUFx10_ASAP7_75t_L g750 ( 
.A(n_735),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_669),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_713),
.B(n_445),
.Y(n_752)
);

AND2x4_ASAP7_75t_L g753 ( 
.A(n_663),
.B(n_615),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_668),
.B(n_615),
.Y(n_754)
);

INVx3_ASAP7_75t_L g755 ( 
.A(n_723),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_736),
.B(n_401),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_679),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_703),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_673),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_690),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_691),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_723),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_718),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_698),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_700),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_705),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_664),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_706),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_703),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_744),
.B(n_615),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_710),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_715),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_664),
.B(n_401),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_720),
.Y(n_774)
);

BUFx2_ASAP7_75t_L g775 ( 
.A(n_711),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_739),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_681),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_725),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_684),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_728),
.Y(n_780)
);

OA21x2_ASAP7_75t_L g781 ( 
.A1(n_739),
.A2(n_524),
.B(n_415),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_730),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_731),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_672),
.B(n_428),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_676),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_677),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_733),
.Y(n_787)
);

OA21x2_ASAP7_75t_L g788 ( 
.A1(n_738),
.A2(n_524),
.B(n_415),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_672),
.B(n_446),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_680),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_682),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_734),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_683),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_717),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_695),
.B(n_708),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_697),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_719),
.Y(n_797)
);

BUFx2_ASAP7_75t_L g798 ( 
.A(n_721),
.Y(n_798)
);

INVx1_ASAP7_75t_SL g799 ( 
.A(n_667),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_703),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_740),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_687),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_688),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_742),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_693),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_696),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_743),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_704),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_707),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_665),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_689),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_712),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_702),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_741),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_741),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_666),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_701),
.B(n_643),
.Y(n_817)
);

OA21x2_ASAP7_75t_L g818 ( 
.A1(n_675),
.A2(n_547),
.B(n_542),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_726),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_692),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_714),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_716),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_709),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_724),
.Y(n_824)
);

CKINVDCx16_ASAP7_75t_R g825 ( 
.A(n_661),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_722),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_729),
.Y(n_827)
);

AND2x2_ASAP7_75t_SL g828 ( 
.A(n_727),
.B(n_643),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_661),
.Y(n_829)
);

OAI21x1_ASAP7_75t_L g830 ( 
.A1(n_732),
.A2(n_547),
.B(n_542),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_737),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_670),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_727),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_670),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_674),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_674),
.B(n_611),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_678),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_678),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_699),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_685),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_685),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_694),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_694),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_699),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_723),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_662),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_R g847 ( 
.A(n_713),
.B(n_657),
.Y(n_847)
);

CKINVDCx20_ASAP7_75t_R g848 ( 
.A(n_727),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_723),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_723),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_686),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_713),
.B(n_453),
.Y(n_852)
);

BUFx2_ASAP7_75t_L g853 ( 
.A(n_711),
.Y(n_853)
);

CKINVDCx20_ASAP7_75t_R g854 ( 
.A(n_727),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_703),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_723),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_723),
.Y(n_857)
);

CKINVDCx20_ASAP7_75t_R g858 ( 
.A(n_727),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_686),
.Y(n_859)
);

CKINVDCx20_ASAP7_75t_R g860 ( 
.A(n_727),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_723),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_723),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_686),
.Y(n_863)
);

OA21x2_ASAP7_75t_L g864 ( 
.A1(n_664),
.A2(n_650),
.B(n_611),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_686),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_723),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_736),
.B(n_650),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_662),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_723),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_686),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_723),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_686),
.Y(n_872)
);

CKINVDCx20_ASAP7_75t_R g873 ( 
.A(n_727),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_703),
.Y(n_874)
);

CKINVDCx16_ASAP7_75t_R g875 ( 
.A(n_713),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_703),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_713),
.B(n_455),
.Y(n_877)
);

BUFx2_ASAP7_75t_L g878 ( 
.A(n_711),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_723),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_686),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_662),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_723),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_662),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_664),
.B(n_656),
.Y(n_884)
);

CKINVDCx14_ASAP7_75t_R g885 ( 
.A(n_713),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_703),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_703),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_686),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_686),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_686),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_662),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_686),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_662),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_794),
.B(n_411),
.Y(n_894)
);

BUFx4f_ASAP7_75t_L g895 ( 
.A(n_798),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_810),
.B(n_447),
.Y(n_896)
);

INVx4_ASAP7_75t_SL g897 ( 
.A(n_817),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_755),
.Y(n_898)
);

INVx4_ASAP7_75t_L g899 ( 
.A(n_755),
.Y(n_899)
);

CKINVDCx11_ASAP7_75t_R g900 ( 
.A(n_848),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_784),
.B(n_400),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_784),
.B(n_402),
.Y(n_902)
);

INVx4_ASAP7_75t_L g903 ( 
.A(n_845),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_796),
.A2(n_643),
.B1(n_442),
.B2(n_448),
.Y(n_904)
);

BUFx6f_ASAP7_75t_SL g905 ( 
.A(n_837),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_814),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_815),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_811),
.B(n_403),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_789),
.B(n_775),
.Y(n_909)
);

INVxp33_ASAP7_75t_L g910 ( 
.A(n_853),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_816),
.B(n_635),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_751),
.A2(n_476),
.B1(n_478),
.B2(n_464),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_750),
.B(n_404),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_878),
.B(n_499),
.Y(n_914)
);

INVx2_ASAP7_75t_SL g915 ( 
.A(n_750),
.Y(n_915)
);

NAND2xp33_ASAP7_75t_L g916 ( 
.A(n_813),
.B(n_553),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_753),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_797),
.A2(n_643),
.B1(n_443),
.B2(n_461),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_SL g919 ( 
.A(n_875),
.B(n_502),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_845),
.Y(n_920)
);

BUFx4f_ASAP7_75t_L g921 ( 
.A(n_837),
.Y(n_921)
);

INVxp67_ASAP7_75t_SL g922 ( 
.A(n_819),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_753),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_885),
.B(n_505),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_754),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_754),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_813),
.B(n_406),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_885),
.B(n_507),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_861),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_823),
.B(n_826),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_L g931 ( 
.A1(n_813),
.A2(n_452),
.B1(n_467),
.B2(n_466),
.Y(n_931)
);

INVxp67_ASAP7_75t_SL g932 ( 
.A(n_861),
.Y(n_932)
);

XNOR2xp5_ASAP7_75t_L g933 ( 
.A(n_848),
.B(n_509),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_749),
.B(n_641),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_762),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_752),
.B(n_644),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_849),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_847),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_770),
.Y(n_939)
);

INVx5_ASAP7_75t_L g940 ( 
.A(n_801),
.Y(n_940)
);

AND2x6_ASAP7_75t_L g941 ( 
.A(n_852),
.B(n_424),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_817),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_L g943 ( 
.A1(n_813),
.A2(n_486),
.B1(n_487),
.B2(n_485),
.Y(n_943)
);

INVx4_ASAP7_75t_SL g944 ( 
.A(n_877),
.Y(n_944)
);

AND2x6_ASAP7_75t_L g945 ( 
.A(n_795),
.B(n_472),
.Y(n_945)
);

INVx5_ASAP7_75t_L g946 ( 
.A(n_801),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_820),
.B(n_647),
.Y(n_947)
);

OAI22xp33_ASAP7_75t_L g948 ( 
.A1(n_799),
.A2(n_522),
.B1(n_535),
.B2(n_512),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_850),
.Y(n_949)
);

INVx5_ASAP7_75t_L g950 ( 
.A(n_801),
.Y(n_950)
);

NOR3xp33_ASAP7_75t_L g951 ( 
.A(n_825),
.B(n_469),
.C(n_462),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_856),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_804),
.B(n_418),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_857),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_862),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_866),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_786),
.Y(n_957)
);

INVxp67_ASAP7_75t_SL g958 ( 
.A(n_788),
.Y(n_958)
);

INVx4_ASAP7_75t_SL g959 ( 
.A(n_770),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_807),
.B(n_760),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_745),
.Y(n_961)
);

AND2x6_ASAP7_75t_L g962 ( 
.A(n_799),
.B(n_472),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_851),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_761),
.B(n_419),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_764),
.B(n_420),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_859),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_801),
.Y(n_967)
);

NAND2xp33_ASAP7_75t_L g968 ( 
.A(n_765),
.B(n_553),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_863),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_766),
.B(n_421),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_865),
.B(n_422),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_781),
.Y(n_972)
);

INVx4_ASAP7_75t_SL g973 ( 
.A(n_831),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_768),
.B(n_425),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_870),
.Y(n_975)
);

INVx4_ASAP7_75t_L g976 ( 
.A(n_786),
.Y(n_976)
);

NAND3xp33_ASAP7_75t_SL g977 ( 
.A(n_847),
.B(n_541),
.C(n_536),
.Y(n_977)
);

AOI22xp33_ASAP7_75t_L g978 ( 
.A1(n_771),
.A2(n_490),
.B1(n_493),
.B2(n_491),
.Y(n_978)
);

OR2x6_ASAP7_75t_L g979 ( 
.A(n_829),
.B(n_494),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_785),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_836),
.B(n_566),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_772),
.B(n_426),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_L g983 ( 
.A1(n_774),
.A2(n_495),
.B1(n_504),
.B2(n_498),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_836),
.B(n_569),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_872),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_880),
.Y(n_986)
);

NAND2xp33_ASAP7_75t_L g987 ( 
.A(n_778),
.B(n_553),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_869),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_888),
.B(n_429),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_780),
.B(n_431),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_782),
.B(n_435),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_783),
.B(n_437),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_889),
.Y(n_993)
);

OR2x2_ASAP7_75t_L g994 ( 
.A(n_834),
.B(n_554),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_787),
.B(n_581),
.Y(n_995)
);

INVx4_ASAP7_75t_L g996 ( 
.A(n_776),
.Y(n_996)
);

INVx4_ASAP7_75t_L g997 ( 
.A(n_776),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_890),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_790),
.Y(n_999)
);

AND2x6_ASAP7_75t_L g1000 ( 
.A(n_792),
.B(n_514),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_871),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_892),
.B(n_441),
.Y(n_1002)
);

INVx4_ASAP7_75t_L g1003 ( 
.A(n_788),
.Y(n_1003)
);

NOR2x1p5_ASAP7_75t_L g1004 ( 
.A(n_763),
.B(n_588),
.Y(n_1004)
);

INVxp67_ASAP7_75t_L g1005 ( 
.A(n_832),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_746),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_818),
.A2(n_508),
.B1(n_517),
.B2(n_510),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_759),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_791),
.Y(n_1009)
);

INVx4_ASAP7_75t_L g1010 ( 
.A(n_879),
.Y(n_1010)
);

BUFx10_ASAP7_75t_L g1011 ( 
.A(n_881),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_793),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_828),
.A2(n_602),
.B1(n_604),
.B2(n_590),
.Y(n_1013)
);

NOR2x1p5_ASAP7_75t_L g1014 ( 
.A(n_763),
.B(n_606),
.Y(n_1014)
);

AOI22xp33_ASAP7_75t_L g1015 ( 
.A1(n_818),
.A2(n_521),
.B1(n_526),
.B2(n_519),
.Y(n_1015)
);

AND2x6_ASAP7_75t_L g1016 ( 
.A(n_756),
.B(n_514),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_SL g1017 ( 
.A1(n_854),
.A2(n_608),
.B1(n_625),
.B2(n_607),
.Y(n_1017)
);

AOI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_828),
.A2(n_634),
.B1(n_640),
.B2(n_629),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_882),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_756),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_867),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_867),
.B(n_833),
.Y(n_1022)
);

BUFx10_ASAP7_75t_L g1023 ( 
.A(n_883),
.Y(n_1023)
);

BUFx10_ASAP7_75t_L g1024 ( 
.A(n_893),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_830),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_781),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_838),
.B(n_444),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_864),
.Y(n_1028)
);

BUFx10_ASAP7_75t_L g1029 ( 
.A(n_846),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_773),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_864),
.B(n_450),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_767),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_773),
.Y(n_1033)
);

INVxp67_ASAP7_75t_SL g1034 ( 
.A(n_884),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_884),
.B(n_451),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_837),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_748),
.Y(n_1037)
);

INVx4_ASAP7_75t_SL g1038 ( 
.A(n_837),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_800),
.Y(n_1039)
);

NAND2xp33_ASAP7_75t_L g1040 ( 
.A(n_846),
.B(n_553),
.Y(n_1040)
);

AOI22xp33_ASAP7_75t_L g1041 ( 
.A1(n_868),
.A2(n_532),
.B1(n_549),
.B2(n_534),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_748),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_824),
.B(n_454),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_748),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_748),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_758),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_758),
.Y(n_1047)
);

INVx4_ASAP7_75t_L g1048 ( 
.A(n_868),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_758),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_827),
.B(n_471),
.Y(n_1050)
);

AND2x6_ASAP7_75t_L g1051 ( 
.A(n_840),
.B(n_552),
.Y(n_1051)
);

INVx4_ASAP7_75t_L g1052 ( 
.A(n_891),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_758),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_769),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_747),
.Y(n_1055)
);

INVx1_ASAP7_75t_SL g1056 ( 
.A(n_757),
.Y(n_1056)
);

INVx2_ASAP7_75t_SL g1057 ( 
.A(n_777),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_769),
.Y(n_1058)
);

INVx5_ASAP7_75t_L g1059 ( 
.A(n_769),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_779),
.B(n_473),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_802),
.B(n_477),
.Y(n_1061)
);

INVx2_ASAP7_75t_SL g1062 ( 
.A(n_803),
.Y(n_1062)
);

INVx2_ASAP7_75t_SL g1063 ( 
.A(n_805),
.Y(n_1063)
);

INVxp67_ASAP7_75t_L g1064 ( 
.A(n_832),
.Y(n_1064)
);

INVx4_ASAP7_75t_L g1065 ( 
.A(n_891),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_769),
.Y(n_1066)
);

NOR3xp33_ASAP7_75t_L g1067 ( 
.A(n_841),
.B(n_843),
.C(n_842),
.Y(n_1067)
);

OR2x6_ASAP7_75t_L g1068 ( 
.A(n_844),
.B(n_556),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_806),
.Y(n_1069)
);

OR2x2_ASAP7_75t_L g1070 ( 
.A(n_808),
.B(n_579),
.Y(n_1070)
);

INVx6_ASAP7_75t_L g1071 ( 
.A(n_855),
.Y(n_1071)
);

BUFx10_ASAP7_75t_L g1072 ( 
.A(n_809),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_855),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_812),
.B(n_479),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_855),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_821),
.A2(n_561),
.B1(n_568),
.B2(n_558),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_822),
.B(n_483),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_887),
.A2(n_584),
.B1(n_597),
.B2(n_577),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_855),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_839),
.B(n_484),
.Y(n_1080)
);

INVx4_ASAP7_75t_L g1081 ( 
.A(n_874),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_874),
.B(n_488),
.Y(n_1082)
);

INVx5_ASAP7_75t_L g1083 ( 
.A(n_874),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_839),
.B(n_642),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_874),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_835),
.B(n_489),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_887),
.A2(n_613),
.B1(n_622),
.B2(n_599),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_876),
.Y(n_1088)
);

NAND2xp33_ASAP7_75t_L g1089 ( 
.A(n_876),
.B(n_553),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_854),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_858),
.B(n_492),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_876),
.B(n_500),
.Y(n_1092)
);

CKINVDCx16_ASAP7_75t_R g1093 ( 
.A(n_858),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_876),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_860),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_886),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_886),
.B(n_501),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_886),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_886),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_860),
.B(n_645),
.Y(n_1100)
);

BUFx4f_ASAP7_75t_L g1101 ( 
.A(n_887),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_887),
.B(n_503),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_873),
.Y(n_1103)
);

HB1xp67_ASAP7_75t_L g1104 ( 
.A(n_873),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_814),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_810),
.A2(n_632),
.B1(n_636),
.B2(n_633),
.Y(n_1106)
);

NAND3xp33_ASAP7_75t_L g1107 ( 
.A(n_784),
.B(n_658),
.C(n_654),
.Y(n_1107)
);

NAND2xp33_ASAP7_75t_L g1108 ( 
.A(n_794),
.B(n_511),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_753),
.Y(n_1109)
);

AND2x4_ASAP7_75t_L g1110 ( 
.A(n_794),
.B(n_617),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_810),
.B(n_513),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_794),
.B(n_515),
.Y(n_1112)
);

BUFx3_ASAP7_75t_L g1113 ( 
.A(n_775),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_847),
.Y(n_1114)
);

NAND2xp33_ASAP7_75t_L g1115 ( 
.A(n_794),
.B(n_516),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_789),
.B(n_438),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_915),
.B(n_527),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_1020),
.B(n_660),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1021),
.B(n_529),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_972),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_976),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_922),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_961),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_963),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_976),
.Y(n_1125)
);

NAND3xp33_ASAP7_75t_L g1126 ( 
.A(n_1007),
.B(n_1015),
.C(n_1107),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_L g1127 ( 
.A1(n_981),
.A2(n_659),
.B1(n_582),
.B2(n_552),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_966),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_969),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_894),
.B(n_1110),
.Y(n_1130)
);

AOI221xp5_ASAP7_75t_L g1131 ( 
.A1(n_930),
.A2(n_531),
.B1(n_537),
.B2(n_533),
.C(n_530),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_996),
.Y(n_1132)
);

NOR3xp33_ASAP7_75t_L g1133 ( 
.A(n_1017),
.B(n_540),
.C(n_538),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_975),
.Y(n_1134)
);

NAND2xp33_ASAP7_75t_L g1135 ( 
.A(n_1000),
.B(n_543),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_894),
.B(n_544),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1110),
.B(n_6),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_984),
.B(n_546),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_948),
.B(n_548),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_1113),
.B(n_895),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_996),
.Y(n_1141)
);

BUFx3_ASAP7_75t_L g1142 ( 
.A(n_1006),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_958),
.A2(n_960),
.B1(n_986),
.B2(n_985),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_909),
.B(n_7),
.Y(n_1144)
);

NOR3x1_ASAP7_75t_L g1145 ( 
.A(n_1069),
.B(n_7),
.C(n_8),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_972),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_1112),
.B(n_550),
.Y(n_1147)
);

NAND2xp33_ASAP7_75t_L g1148 ( 
.A(n_1000),
.B(n_551),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_993),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_998),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_L g1151 ( 
.A1(n_1116),
.A2(n_582),
.B1(n_656),
.B2(n_559),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_972),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_997),
.B(n_562),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1022),
.B(n_570),
.Y(n_1154)
);

AND2x6_ASAP7_75t_SL g1155 ( 
.A(n_1091),
.B(n_8),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_939),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_896),
.B(n_573),
.Y(n_1157)
);

HB1xp67_ASAP7_75t_L g1158 ( 
.A(n_910),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_995),
.B(n_575),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_1005),
.B(n_576),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_957),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1064),
.B(n_580),
.Y(n_1162)
);

NAND2xp33_ASAP7_75t_L g1163 ( 
.A(n_1000),
.B(n_585),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_906),
.B(n_586),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1109),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_925),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_945),
.A2(n_591),
.B1(n_592),
.B2(n_587),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_914),
.B(n_9),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_935),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_1048),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1056),
.B(n_9),
.Y(n_1171)
);

INVxp67_ASAP7_75t_L g1172 ( 
.A(n_919),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_907),
.B(n_593),
.Y(n_1173)
);

INVx4_ASAP7_75t_L g1174 ( 
.A(n_1048),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_997),
.B(n_594),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1105),
.B(n_595),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_917),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_945),
.B(n_596),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_1101),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_945),
.A2(n_942),
.B1(n_1067),
.B2(n_911),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1052),
.B(n_653),
.Y(n_1181)
);

NOR2x1p5_ASAP7_75t_L g1182 ( 
.A(n_1052),
.B(n_601),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_937),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_945),
.B(n_616),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_949),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1008),
.B(n_618),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_923),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_952),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_980),
.B(n_619),
.Y(n_1189)
);

NOR3xp33_ASAP7_75t_L g1190 ( 
.A(n_1093),
.B(n_623),
.C(n_620),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1065),
.B(n_630),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_926),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_921),
.Y(n_1193)
);

AOI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1009),
.A2(n_652),
.B1(n_637),
.B2(n_639),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_954),
.Y(n_1195)
);

OR2x6_ASAP7_75t_L g1196 ( 
.A(n_1065),
.B(n_525),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_999),
.B(n_631),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1106),
.B(n_646),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_899),
.B(n_651),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1080),
.B(n_10),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1012),
.B(n_10),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_899),
.Y(n_1202)
);

INVxp67_ASAP7_75t_L g1203 ( 
.A(n_1070),
.Y(n_1203)
);

INVx5_ASAP7_75t_L g1204 ( 
.A(n_1000),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_1072),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_959),
.Y(n_1206)
);

INVx2_ASAP7_75t_SL g1207 ( 
.A(n_1072),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_903),
.B(n_525),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1115),
.B(n_11),
.Y(n_1209)
);

NAND2xp33_ASAP7_75t_L g1210 ( 
.A(n_962),
.B(n_525),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_SL g1211 ( 
.A(n_1003),
.B(n_560),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_959),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_897),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_SL g1214 ( 
.A(n_1003),
.B(n_560),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1108),
.B(n_11),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_941),
.B(n_901),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_941),
.B(n_12),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1029),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_941),
.B(n_14),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_941),
.B(n_14),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_903),
.B(n_560),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_955),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_953),
.B(n_560),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_902),
.B(n_15),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_964),
.B(n_16),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_965),
.B(n_16),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_956),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_974),
.B(n_17),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_982),
.B(n_17),
.Y(n_1229)
);

OAI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1026),
.A2(n_614),
.B(n_563),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1055),
.B(n_19),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_990),
.B(n_19),
.Y(n_1232)
);

AND2x6_ASAP7_75t_SL g1233 ( 
.A(n_1100),
.B(n_20),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_991),
.B(n_563),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_992),
.B(n_934),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_900),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1011),
.Y(n_1237)
);

INVx5_ASAP7_75t_L g1238 ( 
.A(n_962),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_988),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1001),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_897),
.Y(n_1241)
);

NAND3xp33_ASAP7_75t_L g1242 ( 
.A(n_931),
.B(n_614),
.C(n_563),
.Y(n_1242)
);

AND2x6_ASAP7_75t_L g1243 ( 
.A(n_1025),
.B(n_563),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_1002),
.B(n_614),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_943),
.A2(n_1028),
.B1(n_979),
.B2(n_1018),
.Y(n_1245)
);

INVx8_ASAP7_75t_L g1246 ( 
.A(n_905),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_898),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_936),
.B(n_971),
.Y(n_1248)
);

NOR2x1_ASAP7_75t_L g1249 ( 
.A(n_977),
.B(n_614),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_924),
.B(n_21),
.Y(n_1250)
);

INVxp67_ASAP7_75t_L g1251 ( 
.A(n_962),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_929),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_989),
.B(n_21),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_908),
.B(n_23),
.Y(n_1254)
);

NOR3xp33_ASAP7_75t_L g1255 ( 
.A(n_1095),
.B(n_24),
.C(n_25),
.Y(n_1255)
);

AOI22x1_ASAP7_75t_L g1256 ( 
.A1(n_967),
.A2(n_128),
.B1(n_129),
.B2(n_123),
.Y(n_1256)
);

INVxp67_ASAP7_75t_L g1257 ( 
.A(n_962),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_912),
.B(n_26),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_978),
.B(n_27),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1032),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1016),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_983),
.B(n_28),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1016),
.A2(n_1051),
.B1(n_1010),
.B2(n_979),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1010),
.Y(n_1264)
);

AND2x6_ASAP7_75t_SL g1265 ( 
.A(n_1068),
.B(n_30),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_967),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_913),
.B(n_31),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_932),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1019),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1016),
.B(n_1111),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_928),
.B(n_31),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_967),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_940),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_994),
.B(n_34),
.Y(n_1274)
);

INVxp67_ASAP7_75t_L g1275 ( 
.A(n_1084),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1057),
.B(n_34),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1027),
.B(n_35),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_940),
.Y(n_1278)
);

OAI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1062),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_1279)
);

OAI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1031),
.A2(n_134),
.B(n_131),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_SL g1281 ( 
.A(n_1011),
.Y(n_1281)
);

O2A1O1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_951),
.A2(n_40),
.B(n_36),
.C(n_38),
.Y(n_1282)
);

AND2x6_ASAP7_75t_SL g1283 ( 
.A(n_1068),
.B(n_40),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1016),
.B(n_41),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_920),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_SL g1286 ( 
.A(n_944),
.B(n_41),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_1043),
.B(n_1050),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1051),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1036),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1013),
.B(n_947),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1076),
.B(n_42),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1086),
.B(n_43),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_940),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1041),
.B(n_44),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1051),
.B(n_45),
.Y(n_1295)
);

INVxp67_ASAP7_75t_L g1296 ( 
.A(n_1104),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1060),
.B(n_46),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_946),
.Y(n_1298)
);

NOR2xp67_ASAP7_75t_L g1299 ( 
.A(n_1063),
.B(n_46),
.Y(n_1299)
);

A2O1A1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1030),
.A2(n_1033),
.B(n_1034),
.C(n_918),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_946),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_946),
.Y(n_1302)
);

NOR3xp33_ASAP7_75t_L g1303 ( 
.A(n_1103),
.B(n_47),
.C(n_49),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_904),
.B(n_47),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_950),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1023),
.Y(n_1306)
);

O2A1O1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1130),
.A2(n_1040),
.B(n_927),
.C(n_1061),
.Y(n_1307)
);

OAI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1300),
.A2(n_916),
.B(n_968),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1123),
.B(n_944),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1124),
.B(n_1128),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1211),
.A2(n_1035),
.B(n_987),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1129),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1134),
.B(n_973),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1149),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1211),
.A2(n_970),
.B(n_1082),
.Y(n_1315)
);

BUFx6f_ASAP7_75t_L g1316 ( 
.A(n_1120),
.Y(n_1316)
);

HB1xp67_ASAP7_75t_L g1317 ( 
.A(n_1158),
.Y(n_1317)
);

AOI33xp33_ASAP7_75t_L g1318 ( 
.A1(n_1144),
.A2(n_1078),
.A3(n_1087),
.B1(n_1004),
.B2(n_1014),
.B3(n_933),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1170),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1203),
.B(n_1090),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1150),
.B(n_973),
.Y(n_1321)
);

BUFx8_ASAP7_75t_L g1322 ( 
.A(n_1281),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_R g1323 ( 
.A(n_1236),
.B(n_1237),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_SL g1324 ( 
.A(n_1174),
.B(n_1029),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1122),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1275),
.A2(n_1074),
.B1(n_1077),
.B2(n_938),
.Y(n_1326)
);

O2A1O1Ixp33_ASAP7_75t_L g1327 ( 
.A1(n_1248),
.A2(n_1092),
.B(n_1097),
.C(n_1102),
.Y(n_1327)
);

OAI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1230),
.A2(n_1039),
.B(n_1089),
.Y(n_1328)
);

AOI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1230),
.A2(n_1044),
.B(n_1042),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_SL g1330 ( 
.A(n_1174),
.B(n_1023),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1260),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1177),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1187),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1214),
.A2(n_1046),
.B(n_1045),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1290),
.B(n_1038),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1296),
.B(n_1114),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1192),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1214),
.A2(n_1054),
.B(n_1047),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1268),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_L g1340 ( 
.A(n_1287),
.B(n_1024),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_R g1341 ( 
.A(n_1306),
.B(n_1024),
.Y(n_1341)
);

A2O1A1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1277),
.A2(n_950),
.B(n_1066),
.C(n_1058),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1169),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1235),
.B(n_1038),
.Y(n_1344)
);

O2A1O1Ixp5_ASAP7_75t_L g1345 ( 
.A1(n_1223),
.A2(n_1081),
.B(n_1073),
.C(n_1075),
.Y(n_1345)
);

NOR2x1_ASAP7_75t_L g1346 ( 
.A(n_1205),
.B(n_1081),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1143),
.A2(n_950),
.B1(n_1083),
.B2(n_1059),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_1120),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1168),
.B(n_49),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1137),
.B(n_50),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1156),
.B(n_51),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1201),
.Y(n_1352)
);

A2O1A1Ixp33_ASAP7_75t_L g1353 ( 
.A1(n_1297),
.A2(n_1274),
.B(n_1126),
.C(n_1224),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1142),
.B(n_52),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1218),
.B(n_1059),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1171),
.B(n_55),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1180),
.B(n_55),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1294),
.B(n_56),
.Y(n_1358)
);

BUFx12f_ASAP7_75t_L g1359 ( 
.A(n_1265),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1291),
.B(n_56),
.Y(n_1360)
);

AOI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1250),
.A2(n_1094),
.B1(n_1088),
.B2(n_1071),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_SL g1362 ( 
.A(n_1172),
.B(n_1059),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_SL g1363 ( 
.A(n_1281),
.B(n_1083),
.Y(n_1363)
);

AOI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1271),
.A2(n_1071),
.B1(n_1085),
.B2(n_1079),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1160),
.B(n_57),
.Y(n_1365)
);

NAND2x1p5_ASAP7_75t_L g1366 ( 
.A(n_1207),
.B(n_1083),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1216),
.A2(n_1098),
.B(n_1096),
.Y(n_1367)
);

NOR3xp33_ASAP7_75t_L g1368 ( 
.A(n_1282),
.B(n_1099),
.C(n_57),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1136),
.B(n_58),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1119),
.A2(n_1049),
.B(n_1037),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1186),
.A2(n_1049),
.B(n_1037),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1245),
.B(n_59),
.Y(n_1372)
);

O2A1O1Ixp5_ASAP7_75t_L g1373 ( 
.A1(n_1234),
.A2(n_1049),
.B(n_1053),
.C(n_1037),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1183),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1259),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1258),
.B(n_59),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1138),
.B(n_60),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1120),
.Y(n_1378)
);

A2O1A1Ixp33_ASAP7_75t_L g1379 ( 
.A1(n_1126),
.A2(n_1053),
.B(n_63),
.C(n_61),
.Y(n_1379)
);

NOR3xp33_ASAP7_75t_L g1380 ( 
.A(n_1303),
.B(n_61),
.C(n_62),
.Y(n_1380)
);

A2O1A1Ixp33_ASAP7_75t_L g1381 ( 
.A1(n_1292),
.A2(n_1053),
.B(n_67),
.C(n_62),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1280),
.A2(n_138),
.B(n_135),
.Y(n_1382)
);

AO21x2_ASAP7_75t_L g1383 ( 
.A1(n_1280),
.A2(n_142),
.B(n_140),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1262),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1151),
.B(n_65),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1164),
.A2(n_144),
.B(n_143),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1173),
.A2(n_147),
.B(n_145),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1176),
.A2(n_152),
.B(n_150),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1146),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1270),
.A2(n_155),
.B(n_153),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1185),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1140),
.B(n_1162),
.Y(n_1392)
);

NAND2x1p5_ASAP7_75t_L g1393 ( 
.A(n_1179),
.B(n_68),
.Y(n_1393)
);

BUFx6f_ASAP7_75t_L g1394 ( 
.A(n_1146),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1231),
.B(n_69),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1276),
.B(n_69),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1133),
.B(n_1182),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1154),
.A2(n_158),
.B(n_157),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1159),
.B(n_70),
.Y(n_1399)
);

INVx3_ASAP7_75t_L g1400 ( 
.A(n_1302),
.Y(n_1400)
);

NAND3xp33_ASAP7_75t_L g1401 ( 
.A(n_1255),
.B(n_70),
.C(n_71),
.Y(n_1401)
);

INVx2_ASAP7_75t_SL g1402 ( 
.A(n_1246),
.Y(n_1402)
);

NAND3xp33_ASAP7_75t_L g1403 ( 
.A(n_1249),
.B(n_1210),
.C(n_1288),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1266),
.A2(n_163),
.B(n_160),
.Y(n_1404)
);

A2O1A1Ixp33_ASAP7_75t_L g1405 ( 
.A1(n_1225),
.A2(n_1226),
.B(n_1229),
.C(n_1228),
.Y(n_1405)
);

OAI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1232),
.A2(n_169),
.B(n_168),
.Y(n_1406)
);

BUFx2_ASAP7_75t_L g1407 ( 
.A(n_1196),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1127),
.B(n_71),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1194),
.B(n_1200),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_1246),
.Y(n_1410)
);

AOI22x1_ASAP7_75t_L g1411 ( 
.A1(n_1272),
.A2(n_172),
.B1(n_177),
.B2(n_171),
.Y(n_1411)
);

INVx11_ASAP7_75t_L g1412 ( 
.A(n_1246),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1118),
.A2(n_183),
.B(n_180),
.Y(n_1413)
);

A2O1A1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1253),
.A2(n_74),
.B(n_72),
.C(n_73),
.Y(n_1414)
);

O2A1O1Ixp33_ASAP7_75t_L g1415 ( 
.A1(n_1254),
.A2(n_74),
.B(n_72),
.C(n_73),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1147),
.A2(n_185),
.B(n_184),
.Y(n_1416)
);

INVx3_ASAP7_75t_L g1417 ( 
.A(n_1302),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1285),
.B(n_75),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1213),
.B(n_75),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1188),
.A2(n_188),
.B(n_186),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1194),
.B(n_1165),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1161),
.B(n_77),
.Y(n_1422)
);

OAI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1195),
.A2(n_190),
.B(n_189),
.Y(n_1423)
);

AOI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1190),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1222),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1227),
.A2(n_193),
.B(n_191),
.Y(n_1426)
);

OAI321xp33_ASAP7_75t_L g1427 ( 
.A1(n_1279),
.A2(n_80),
.A3(n_81),
.B1(n_82),
.B2(n_83),
.C(n_84),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_SL g1428 ( 
.A(n_1179),
.B(n_84),
.Y(n_1428)
);

OAI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1239),
.A2(n_195),
.B(n_194),
.Y(n_1429)
);

OR2x6_ASAP7_75t_SL g1430 ( 
.A(n_1265),
.B(n_85),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1240),
.A2(n_197),
.B(n_196),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_1146),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1152),
.A2(n_199),
.B(n_198),
.Y(n_1433)
);

NAND3xp33_ASAP7_75t_SL g1434 ( 
.A(n_1263),
.B(n_85),
.C(n_86),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1256),
.A2(n_201),
.B(n_200),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1166),
.B(n_86),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1132),
.B(n_87),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_L g1438 ( 
.A(n_1198),
.B(n_88),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1131),
.A2(n_89),
.B1(n_90),
.B2(n_92),
.Y(n_1439)
);

BUFx3_ASAP7_75t_L g1440 ( 
.A(n_1302),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1132),
.B(n_89),
.Y(n_1441)
);

INVx2_ASAP7_75t_SL g1442 ( 
.A(n_1179),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_1152),
.Y(n_1443)
);

BUFx4f_ASAP7_75t_L g1444 ( 
.A(n_1196),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1193),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1141),
.B(n_90),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1152),
.A2(n_203),
.B(n_202),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1264),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1157),
.B(n_96),
.Y(n_1449)
);

O2A1O1Ixp33_ASAP7_75t_L g1450 ( 
.A1(n_1209),
.A2(n_96),
.B(n_97),
.C(n_98),
.Y(n_1450)
);

NAND3xp33_ASAP7_75t_L g1451 ( 
.A(n_1261),
.B(n_98),
.C(n_99),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1208),
.A2(n_207),
.B(n_206),
.Y(n_1452)
);

INVx2_ASAP7_75t_SL g1453 ( 
.A(n_1241),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1141),
.B(n_100),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1312),
.B(n_1267),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1329),
.A2(n_1371),
.B(n_1370),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1314),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1353),
.A2(n_1304),
.B(n_1215),
.Y(n_1458)
);

AOI21xp33_ASAP7_75t_L g1459 ( 
.A1(n_1344),
.A2(n_1196),
.B(n_1217),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1334),
.A2(n_1221),
.B(n_1244),
.Y(n_1460)
);

AOI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1405),
.A2(n_1148),
.B(n_1135),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1311),
.A2(n_1163),
.B(n_1219),
.Y(n_1462)
);

NAND2x1_ASAP7_75t_L g1463 ( 
.A(n_1400),
.B(n_1243),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1338),
.A2(n_1284),
.B(n_1202),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1308),
.A2(n_1220),
.B(n_1251),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1315),
.A2(n_1257),
.B(n_1289),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1444),
.A2(n_1204),
.B1(n_1167),
.B2(n_1238),
.Y(n_1467)
);

AOI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1367),
.A2(n_1328),
.B(n_1335),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1373),
.A2(n_1202),
.B(n_1247),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1332),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1337),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1382),
.A2(n_1252),
.B(n_1295),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1325),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1310),
.B(n_1145),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1333),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1339),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1340),
.B(n_1299),
.Y(n_1477)
);

OAI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1349),
.A2(n_1204),
.B1(n_1238),
.B2(n_1178),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1342),
.A2(n_1199),
.B(n_1175),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1318),
.B(n_1269),
.Y(n_1480)
);

OAI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1409),
.A2(n_1139),
.B(n_1184),
.Y(n_1481)
);

OAI22x1_ASAP7_75t_L g1482 ( 
.A1(n_1419),
.A2(n_1283),
.B1(n_1233),
.B2(n_1155),
.Y(n_1482)
);

INVx6_ASAP7_75t_SL g1483 ( 
.A(n_1419),
.Y(n_1483)
);

AOI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1372),
.A2(n_1286),
.B(n_1242),
.Y(n_1484)
);

BUFx4f_ASAP7_75t_L g1485 ( 
.A(n_1359),
.Y(n_1485)
);

NAND2xp33_ASAP7_75t_L g1486 ( 
.A(n_1341),
.B(n_1204),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1421),
.B(n_1369),
.Y(n_1487)
);

AOI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1368),
.A2(n_1212),
.B1(n_1206),
.B2(n_1181),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1319),
.B(n_1189),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1375),
.B(n_1384),
.Y(n_1490)
);

AOI21xp5_ASAP7_75t_SL g1491 ( 
.A1(n_1316),
.A2(n_1243),
.B(n_1242),
.Y(n_1491)
);

O2A1O1Ixp5_ASAP7_75t_L g1492 ( 
.A1(n_1362),
.A2(n_1191),
.B(n_1153),
.C(n_1117),
.Y(n_1492)
);

AOI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1403),
.A2(n_1197),
.B(n_1273),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1435),
.A2(n_1125),
.B(n_1121),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1352),
.A2(n_1238),
.B(n_1278),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1407),
.A2(n_1305),
.B1(n_1301),
.B2(n_1298),
.Y(n_1496)
);

AOI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1307),
.A2(n_1293),
.B(n_1243),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1392),
.B(n_1397),
.Y(n_1498)
);

OA21x2_ASAP7_75t_L g1499 ( 
.A1(n_1406),
.A2(n_1243),
.B(n_210),
.Y(n_1499)
);

AOI21x1_ASAP7_75t_L g1500 ( 
.A1(n_1347),
.A2(n_1155),
.B(n_1233),
.Y(n_1500)
);

OAI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1438),
.A2(n_1283),
.B(n_101),
.Y(n_1501)
);

BUFx6f_ASAP7_75t_L g1502 ( 
.A(n_1316),
.Y(n_1502)
);

OA21x2_ASAP7_75t_L g1503 ( 
.A1(n_1423),
.A2(n_211),
.B(n_209),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1351),
.Y(n_1504)
);

INVx3_ASAP7_75t_L g1505 ( 
.A(n_1440),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1365),
.B(n_102),
.Y(n_1506)
);

AOI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1327),
.A2(n_213),
.B(n_212),
.Y(n_1507)
);

AOI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1380),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1345),
.A2(n_1447),
.B(n_1433),
.Y(n_1509)
);

AOI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1377),
.A2(n_220),
.B(n_216),
.Y(n_1510)
);

INVxp67_ASAP7_75t_SL g1511 ( 
.A(n_1317),
.Y(n_1511)
);

OAI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1376),
.A2(n_104),
.B(n_105),
.Y(n_1512)
);

AOI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1358),
.A2(n_233),
.B(n_232),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1356),
.B(n_106),
.Y(n_1514)
);

BUFx2_ASAP7_75t_SL g1515 ( 
.A(n_1402),
.Y(n_1515)
);

CKINVDCx16_ASAP7_75t_R g1516 ( 
.A(n_1323),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1331),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1320),
.B(n_106),
.Y(n_1518)
);

AOI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1439),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1411),
.A2(n_236),
.B(n_235),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1399),
.A2(n_1360),
.B(n_1383),
.Y(n_1521)
);

INVxp67_ASAP7_75t_L g1522 ( 
.A(n_1354),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1449),
.B(n_107),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1343),
.Y(n_1524)
);

A2O1A1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1415),
.A2(n_109),
.B(n_110),
.C(n_111),
.Y(n_1525)
);

O2A1O1Ixp5_ASAP7_75t_L g1526 ( 
.A1(n_1357),
.A2(n_330),
.B(n_399),
.C(n_398),
.Y(n_1526)
);

AO21x2_ASAP7_75t_L g1527 ( 
.A1(n_1379),
.A2(n_239),
.B(n_237),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1350),
.B(n_111),
.Y(n_1528)
);

OAI21x1_ASAP7_75t_L g1529 ( 
.A1(n_1390),
.A2(n_241),
.B(n_240),
.Y(n_1529)
);

OAI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1385),
.A2(n_112),
.B(n_113),
.Y(n_1530)
);

OAI21x1_ASAP7_75t_L g1531 ( 
.A1(n_1429),
.A2(n_243),
.B(n_242),
.Y(n_1531)
);

OAI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1408),
.A2(n_112),
.B(n_113),
.Y(n_1532)
);

OAI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1395),
.A2(n_114),
.B(n_115),
.Y(n_1533)
);

OAI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1398),
.A2(n_332),
.B(n_397),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1418),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1374),
.Y(n_1536)
);

AOI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1316),
.A2(n_333),
.B(n_396),
.Y(n_1537)
);

AOI21xp5_ASAP7_75t_L g1538 ( 
.A1(n_1348),
.A2(n_331),
.B(n_394),
.Y(n_1538)
);

BUFx6f_ASAP7_75t_L g1539 ( 
.A(n_1348),
.Y(n_1539)
);

INVxp67_ASAP7_75t_SL g1540 ( 
.A(n_1348),
.Y(n_1540)
);

INVx1_ASAP7_75t_SL g1541 ( 
.A(n_1410),
.Y(n_1541)
);

OAI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1396),
.A2(n_116),
.B(n_118),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1378),
.A2(n_337),
.B(n_392),
.Y(n_1543)
);

NAND3xp33_ASAP7_75t_L g1544 ( 
.A(n_1401),
.B(n_1381),
.C(n_1414),
.Y(n_1544)
);

O2A1O1Ixp33_ASAP7_75t_L g1545 ( 
.A1(n_1501),
.A2(n_1434),
.B(n_1450),
.C(n_1336),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1511),
.Y(n_1546)
);

AOI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1521),
.A2(n_1389),
.B(n_1378),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1482),
.A2(n_1451),
.B1(n_1422),
.B2(n_1424),
.Y(n_1548)
);

AOI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1461),
.A2(n_1389),
.B(n_1378),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1490),
.B(n_1391),
.Y(n_1550)
);

BUFx10_ASAP7_75t_L g1551 ( 
.A(n_1516),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1457),
.B(n_1425),
.Y(n_1552)
);

INVx4_ASAP7_75t_L g1553 ( 
.A(n_1485),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1483),
.A2(n_1430),
.B1(n_1393),
.B2(n_1448),
.Y(n_1554)
);

BUFx4f_ASAP7_75t_SL g1555 ( 
.A(n_1483),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1473),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1475),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1470),
.B(n_1326),
.Y(n_1558)
);

BUFx12f_ASAP7_75t_L g1559 ( 
.A(n_1485),
.Y(n_1559)
);

NOR2x1_ASAP7_75t_SL g1560 ( 
.A(n_1467),
.B(n_1389),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1498),
.A2(n_1428),
.B1(n_1436),
.B2(n_1454),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1476),
.B(n_1400),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1502),
.Y(n_1563)
);

AOI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1462),
.A2(n_1432),
.B(n_1394),
.Y(n_1564)
);

AOI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1458),
.A2(n_1432),
.B(n_1394),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1474),
.A2(n_1446),
.B1(n_1437),
.B2(n_1441),
.Y(n_1566)
);

CKINVDCx20_ASAP7_75t_R g1567 ( 
.A(n_1541),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1505),
.Y(n_1568)
);

BUFx4f_ASAP7_75t_SL g1569 ( 
.A(n_1505),
.Y(n_1569)
);

INVx6_ASAP7_75t_L g1570 ( 
.A(n_1489),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1471),
.B(n_1417),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1487),
.B(n_1445),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1480),
.B(n_1442),
.Y(n_1573)
);

CKINVDCx20_ASAP7_75t_R g1574 ( 
.A(n_1515),
.Y(n_1574)
);

AOI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1499),
.A2(n_1432),
.B(n_1394),
.Y(n_1575)
);

OR2x6_ASAP7_75t_L g1576 ( 
.A(n_1463),
.B(n_1500),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1524),
.Y(n_1577)
);

AOI21xp5_ASAP7_75t_SL g1578 ( 
.A1(n_1499),
.A2(n_1443),
.B(n_1321),
.Y(n_1578)
);

INVx2_ASAP7_75t_R g1579 ( 
.A(n_1504),
.Y(n_1579)
);

INVx3_ASAP7_75t_L g1580 ( 
.A(n_1502),
.Y(n_1580)
);

NOR2x1_ASAP7_75t_SL g1581 ( 
.A(n_1496),
.B(n_1443),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1517),
.Y(n_1582)
);

AOI222xp33_ASAP7_75t_L g1583 ( 
.A1(n_1522),
.A2(n_1427),
.B1(n_1322),
.B2(n_1324),
.C1(n_1330),
.C2(n_1309),
.Y(n_1583)
);

NAND2x1p5_ASAP7_75t_L g1584 ( 
.A(n_1502),
.B(n_1417),
.Y(n_1584)
);

OAI21xp33_ASAP7_75t_L g1585 ( 
.A1(n_1508),
.A2(n_1363),
.B(n_1313),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1536),
.Y(n_1586)
);

AOI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1519),
.A2(n_1355),
.B1(n_1322),
.B2(n_1453),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1455),
.B(n_1355),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1514),
.Y(n_1589)
);

INVx4_ASAP7_75t_L g1590 ( 
.A(n_1539),
.Y(n_1590)
);

BUFx3_ASAP7_75t_L g1591 ( 
.A(n_1539),
.Y(n_1591)
);

INVx3_ASAP7_75t_L g1592 ( 
.A(n_1576),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1577),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1552),
.Y(n_1594)
);

CKINVDCx16_ASAP7_75t_R g1595 ( 
.A(n_1574),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1552),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1554),
.A2(n_1508),
.B1(n_1542),
.B2(n_1533),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1554),
.A2(n_1544),
.B1(n_1519),
.B2(n_1523),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1556),
.Y(n_1599)
);

INVx8_ASAP7_75t_L g1600 ( 
.A(n_1576),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1590),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1586),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1557),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1582),
.B(n_1512),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1546),
.B(n_1530),
.Y(n_1605)
);

BUFx4f_ASAP7_75t_SL g1606 ( 
.A(n_1559),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1571),
.Y(n_1607)
);

BUFx6f_ASAP7_75t_L g1608 ( 
.A(n_1576),
.Y(n_1608)
);

BUFx6f_ASAP7_75t_SL g1609 ( 
.A(n_1553),
.Y(n_1609)
);

OR2x6_ASAP7_75t_L g1610 ( 
.A(n_1578),
.B(n_1491),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1571),
.Y(n_1611)
);

INVx3_ASAP7_75t_L g1612 ( 
.A(n_1590),
.Y(n_1612)
);

AND2x4_ASAP7_75t_L g1613 ( 
.A(n_1560),
.B(n_1456),
.Y(n_1613)
);

INVx3_ASAP7_75t_L g1614 ( 
.A(n_1580),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1580),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1563),
.Y(n_1616)
);

BUFx8_ASAP7_75t_L g1617 ( 
.A(n_1568),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1563),
.Y(n_1618)
);

CKINVDCx20_ASAP7_75t_R g1619 ( 
.A(n_1567),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1550),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_SL g1621 ( 
.A1(n_1570),
.A2(n_1532),
.B1(n_1544),
.B2(n_1486),
.Y(n_1621)
);

BUFx12f_ASAP7_75t_L g1622 ( 
.A(n_1553),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1570),
.A2(n_1477),
.B1(n_1488),
.B2(n_1518),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1620),
.B(n_1579),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1593),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1616),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1593),
.Y(n_1627)
);

BUFx3_ASAP7_75t_L g1628 ( 
.A(n_1617),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1599),
.Y(n_1629)
);

INVx2_ASAP7_75t_SL g1630 ( 
.A(n_1600),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1617),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1620),
.B(n_1464),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1616),
.Y(n_1633)
);

INVx3_ASAP7_75t_L g1634 ( 
.A(n_1613),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1599),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1594),
.B(n_1589),
.Y(n_1636)
);

OA21x2_ASAP7_75t_L g1637 ( 
.A1(n_1598),
.A2(n_1575),
.B(n_1494),
.Y(n_1637)
);

INVx3_ASAP7_75t_L g1638 ( 
.A(n_1613),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1618),
.Y(n_1639)
);

INVx1_ASAP7_75t_SL g1640 ( 
.A(n_1601),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1602),
.Y(n_1641)
);

INVx3_ASAP7_75t_L g1642 ( 
.A(n_1613),
.Y(n_1642)
);

BUFx3_ASAP7_75t_L g1643 ( 
.A(n_1617),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1602),
.Y(n_1644)
);

INVx3_ASAP7_75t_L g1645 ( 
.A(n_1613),
.Y(n_1645)
);

OR2x6_ASAP7_75t_L g1646 ( 
.A(n_1600),
.B(n_1547),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1603),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1603),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1607),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1607),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1611),
.Y(n_1651)
);

BUFx3_ASAP7_75t_L g1652 ( 
.A(n_1617),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1651),
.B(n_1592),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1647),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1647),
.Y(n_1655)
);

BUFx3_ASAP7_75t_L g1656 ( 
.A(n_1628),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1644),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1644),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1651),
.B(n_1592),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1648),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1648),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1649),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1651),
.B(n_1592),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1641),
.Y(n_1664)
);

INVx2_ASAP7_75t_SL g1665 ( 
.A(n_1628),
.Y(n_1665)
);

AND2x4_ASAP7_75t_L g1666 ( 
.A(n_1634),
.B(n_1638),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1644),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1627),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1649),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1650),
.Y(n_1670)
);

BUFx6f_ASAP7_75t_L g1671 ( 
.A(n_1646),
.Y(n_1671)
);

OAI221xp5_ASAP7_75t_L g1672 ( 
.A1(n_1636),
.A2(n_1597),
.B1(n_1587),
.B2(n_1623),
.C(n_1621),
.Y(n_1672)
);

AOI22xp33_ASAP7_75t_SL g1673 ( 
.A1(n_1628),
.A2(n_1604),
.B1(n_1600),
.B2(n_1605),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1640),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1641),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1672),
.A2(n_1604),
.B1(n_1605),
.B2(n_1643),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1662),
.B(n_1650),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1653),
.B(n_1634),
.Y(n_1678)
);

OAI221xp5_ASAP7_75t_SL g1679 ( 
.A1(n_1673),
.A2(n_1548),
.B1(n_1631),
.B2(n_1545),
.C(n_1643),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1665),
.B(n_1640),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1656),
.A2(n_1643),
.B1(n_1652),
.B2(n_1583),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1669),
.B(n_1636),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1670),
.B(n_1624),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1665),
.B(n_1624),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1660),
.B(n_1624),
.Y(n_1685)
);

AOI221x1_ASAP7_75t_SL g1686 ( 
.A1(n_1660),
.A2(n_1558),
.B1(n_1572),
.B2(n_1596),
.C(n_1594),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1661),
.B(n_1596),
.Y(n_1687)
);

NAND4xp25_ASAP7_75t_L g1688 ( 
.A(n_1656),
.B(n_1583),
.C(n_1652),
.D(n_1566),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1661),
.B(n_1632),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1674),
.B(n_1634),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1654),
.B(n_1655),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1653),
.B(n_1634),
.Y(n_1692)
);

AND2x4_ASAP7_75t_SL g1693 ( 
.A(n_1681),
.B(n_1551),
.Y(n_1693)
);

INVx5_ASAP7_75t_L g1694 ( 
.A(n_1680),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1678),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1691),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1684),
.B(n_1666),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1692),
.B(n_1666),
.Y(n_1698)
);

INVxp67_ASAP7_75t_L g1699 ( 
.A(n_1688),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1689),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1685),
.B(n_1659),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1683),
.B(n_1682),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1677),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1686),
.B(n_1659),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1678),
.B(n_1663),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1690),
.B(n_1663),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1687),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1681),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1676),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1676),
.B(n_1666),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1679),
.B(n_1657),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1685),
.B(n_1657),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1703),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_SL g1714 ( 
.A(n_1694),
.B(n_1595),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1697),
.B(n_1671),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1708),
.B(n_1664),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1702),
.B(n_1658),
.Y(n_1717)
);

AND3x2_ASAP7_75t_L g1718 ( 
.A(n_1699),
.B(n_1609),
.C(n_1606),
.Y(n_1718)
);

AOI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1708),
.A2(n_1709),
.B1(n_1711),
.B2(n_1704),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1697),
.B(n_1710),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1703),
.B(n_1664),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1696),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1721),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1720),
.B(n_1694),
.Y(n_1724)
);

OAI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1719),
.A2(n_1694),
.B(n_1619),
.Y(n_1725)
);

INVx1_ASAP7_75t_SL g1726 ( 
.A(n_1718),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1722),
.Y(n_1727)
);

OAI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1714),
.A2(n_1652),
.B1(n_1595),
.B2(n_1630),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1727),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1726),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1723),
.B(n_1719),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1728),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1730),
.B(n_1725),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1732),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1729),
.B(n_1731),
.Y(n_1735)
);

INVx2_ASAP7_75t_SL g1736 ( 
.A(n_1730),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1736),
.B(n_1724),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1733),
.B(n_1718),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1734),
.B(n_1716),
.Y(n_1739)
);

INVxp67_ASAP7_75t_SL g1740 ( 
.A(n_1735),
.Y(n_1740)
);

NAND2x1p5_ASAP7_75t_L g1741 ( 
.A(n_1735),
.B(n_1551),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1736),
.B(n_1728),
.Y(n_1742)
);

O2A1O1Ixp33_ASAP7_75t_L g1743 ( 
.A1(n_1740),
.A2(n_1525),
.B(n_1506),
.C(n_1366),
.Y(n_1743)
);

OAI32xp33_ASAP7_75t_L g1744 ( 
.A1(n_1742),
.A2(n_1713),
.A3(n_1717),
.B1(n_1715),
.B2(n_1695),
.Y(n_1744)
);

AOI322xp5_ASAP7_75t_L g1745 ( 
.A1(n_1738),
.A2(n_1737),
.A3(n_1739),
.B1(n_1741),
.B2(n_1622),
.C1(n_1700),
.C2(n_1707),
.Y(n_1745)
);

AOI221xp5_ASAP7_75t_L g1746 ( 
.A1(n_1742),
.A2(n_1693),
.B1(n_1609),
.B2(n_1700),
.C(n_1585),
.Y(n_1746)
);

AOI21xp33_ASAP7_75t_SL g1747 ( 
.A1(n_1741),
.A2(n_120),
.B(n_121),
.Y(n_1747)
);

OAI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1742),
.A2(n_1535),
.B(n_1492),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1742),
.B(n_1712),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1742),
.B(n_1701),
.Y(n_1750)
);

OAI211xp5_ASAP7_75t_L g1751 ( 
.A1(n_1740),
.A2(n_1412),
.B(n_1555),
.C(n_1622),
.Y(n_1751)
);

OAI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1742),
.A2(n_1609),
.B1(n_1705),
.B2(n_1706),
.Y(n_1752)
);

NOR4xp25_ASAP7_75t_L g1753 ( 
.A(n_1751),
.B(n_1528),
.C(n_1561),
.D(n_1481),
.Y(n_1753)
);

NAND3xp33_ASAP7_75t_L g1754 ( 
.A(n_1745),
.B(n_1346),
.C(n_1479),
.Y(n_1754)
);

INVxp33_ASAP7_75t_L g1755 ( 
.A(n_1747),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1749),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1750),
.B(n_1698),
.Y(n_1757)
);

BUFx2_ASAP7_75t_L g1758 ( 
.A(n_1746),
.Y(n_1758)
);

NOR3xp33_ASAP7_75t_SL g1759 ( 
.A(n_1744),
.B(n_1413),
.C(n_1416),
.Y(n_1759)
);

NOR3xp33_ASAP7_75t_L g1760 ( 
.A(n_1748),
.B(n_1459),
.C(n_1526),
.Y(n_1760)
);

NAND3xp33_ASAP7_75t_L g1761 ( 
.A(n_1752),
.B(n_1488),
.C(n_1510),
.Y(n_1761)
);

AO22x2_ASAP7_75t_L g1762 ( 
.A1(n_1743),
.A2(n_1588),
.B1(n_1601),
.B2(n_1612),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1747),
.B(n_1675),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1749),
.Y(n_1764)
);

OAI211xp5_ASAP7_75t_L g1765 ( 
.A1(n_1751),
.A2(n_1569),
.B(n_1573),
.C(n_1671),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1749),
.Y(n_1766)
);

NAND3xp33_ASAP7_75t_L g1767 ( 
.A(n_1745),
.B(n_1513),
.C(n_1507),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1749),
.Y(n_1768)
);

NAND3xp33_ASAP7_75t_L g1769 ( 
.A(n_1745),
.B(n_1538),
.C(n_1537),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1755),
.B(n_1601),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_L g1771 ( 
.A(n_1758),
.B(n_1612),
.Y(n_1771)
);

NAND4xp75_ASAP7_75t_L g1772 ( 
.A(n_1756),
.B(n_1543),
.C(n_1503),
.D(n_1630),
.Y(n_1772)
);

AND4x1_ASAP7_75t_L g1773 ( 
.A(n_1753),
.B(n_1386),
.C(n_1387),
.D(n_1388),
.Y(n_1773)
);

NOR3xp33_ASAP7_75t_L g1774 ( 
.A(n_1765),
.B(n_1754),
.C(n_1769),
.Y(n_1774)
);

NAND4xp25_ASAP7_75t_L g1775 ( 
.A(n_1764),
.B(n_1591),
.C(n_1612),
.D(n_1592),
.Y(n_1775)
);

NAND4xp25_ASAP7_75t_L g1776 ( 
.A(n_1766),
.B(n_1612),
.C(n_1495),
.D(n_1550),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1757),
.B(n_1671),
.Y(n_1777)
);

NOR3xp33_ASAP7_75t_L g1778 ( 
.A(n_1768),
.B(n_1426),
.C(n_1420),
.Y(n_1778)
);

AOI221xp5_ASAP7_75t_L g1779 ( 
.A1(n_1762),
.A2(n_1562),
.B1(n_1671),
.B2(n_1614),
.C(n_1615),
.Y(n_1779)
);

NAND3xp33_ASAP7_75t_L g1780 ( 
.A(n_1759),
.B(n_1767),
.C(n_1760),
.Y(n_1780)
);

OAI221xp5_ASAP7_75t_L g1781 ( 
.A1(n_1763),
.A2(n_1761),
.B1(n_1762),
.B2(n_1671),
.C(n_1630),
.Y(n_1781)
);

AOI221xp5_ASAP7_75t_L g1782 ( 
.A1(n_1753),
.A2(n_1562),
.B1(n_1614),
.B2(n_1615),
.C(n_1675),
.Y(n_1782)
);

AOI33xp33_ASAP7_75t_L g1783 ( 
.A1(n_1756),
.A2(n_1611),
.A3(n_1618),
.B1(n_1632),
.B2(n_1629),
.B3(n_1625),
.Y(n_1783)
);

NOR3x1_ASAP7_75t_L g1784 ( 
.A(n_1758),
.B(n_1534),
.C(n_1478),
.Y(n_1784)
);

NOR2xp33_ASAP7_75t_L g1785 ( 
.A(n_1755),
.B(n_1614),
.Y(n_1785)
);

NOR3xp33_ASAP7_75t_L g1786 ( 
.A(n_1765),
.B(n_1431),
.C(n_1520),
.Y(n_1786)
);

NAND4xp25_ASAP7_75t_L g1787 ( 
.A(n_1756),
.B(n_1642),
.C(n_1638),
.D(n_1645),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1780),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1771),
.B(n_1774),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1777),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1770),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1776),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1784),
.B(n_1638),
.Y(n_1793)
);

NOR2xp33_ASAP7_75t_L g1794 ( 
.A(n_1781),
.B(n_1614),
.Y(n_1794)
);

NOR2x1_ASAP7_75t_L g1795 ( 
.A(n_1785),
.B(n_1404),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1772),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1783),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1773),
.Y(n_1798)
);

AOI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1775),
.A2(n_1527),
.B1(n_1610),
.B2(n_1608),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1782),
.Y(n_1800)
);

INVx1_ASAP7_75t_SL g1801 ( 
.A(n_1778),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1787),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1779),
.B(n_1638),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1786),
.B(n_1642),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1780),
.Y(n_1805)
);

INVxp67_ASAP7_75t_L g1806 ( 
.A(n_1780),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_L g1807 ( 
.A(n_1806),
.B(n_1608),
.Y(n_1807)
);

NAND3xp33_ASAP7_75t_SL g1808 ( 
.A(n_1788),
.B(n_1805),
.C(n_1801),
.Y(n_1808)
);

NOR2x1_ASAP7_75t_L g1809 ( 
.A(n_1789),
.B(n_1452),
.Y(n_1809)
);

BUFx3_ASAP7_75t_L g1810 ( 
.A(n_1790),
.Y(n_1810)
);

NOR3xp33_ASAP7_75t_L g1811 ( 
.A(n_1798),
.B(n_1531),
.C(n_1361),
.Y(n_1811)
);

NAND4xp25_ASAP7_75t_L g1812 ( 
.A(n_1791),
.B(n_1497),
.C(n_1645),
.D(n_1642),
.Y(n_1812)
);

NOR3x1_ASAP7_75t_L g1813 ( 
.A(n_1792),
.B(n_1529),
.C(n_1509),
.Y(n_1813)
);

NOR2xp33_ASAP7_75t_SL g1814 ( 
.A(n_1796),
.B(n_1608),
.Y(n_1814)
);

NOR3xp33_ASAP7_75t_L g1815 ( 
.A(n_1800),
.B(n_1364),
.C(n_1493),
.Y(n_1815)
);

NAND2xp33_ASAP7_75t_L g1816 ( 
.A(n_1802),
.B(n_1608),
.Y(n_1816)
);

AND2x2_ASAP7_75t_SL g1817 ( 
.A(n_1797),
.B(n_1503),
.Y(n_1817)
);

NAND4xp75_ASAP7_75t_L g1818 ( 
.A(n_1795),
.B(n_1565),
.C(n_1466),
.D(n_1549),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1804),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1803),
.B(n_1642),
.Y(n_1820)
);

NOR2x1_ASAP7_75t_L g1821 ( 
.A(n_1794),
.B(n_1527),
.Y(n_1821)
);

XOR2x1_ASAP7_75t_SL g1822 ( 
.A(n_1808),
.B(n_1793),
.Y(n_1822)
);

NOR3xp33_ASAP7_75t_L g1823 ( 
.A(n_1810),
.B(n_1799),
.C(n_1484),
.Y(n_1823)
);

AOI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1807),
.A2(n_1799),
.B1(n_1600),
.B2(n_1608),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1818),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_SL g1826 ( 
.A(n_1814),
.B(n_1539),
.Y(n_1826)
);

XNOR2xp5_ASAP7_75t_L g1827 ( 
.A(n_1819),
.B(n_1584),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1820),
.Y(n_1828)
);

AND2x4_ASAP7_75t_L g1829 ( 
.A(n_1809),
.B(n_1645),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1821),
.B(n_1645),
.Y(n_1830)
);

HB1xp67_ASAP7_75t_L g1831 ( 
.A(n_1817),
.Y(n_1831)
);

BUFx2_ASAP7_75t_L g1832 ( 
.A(n_1812),
.Y(n_1832)
);

NAND4xp75_ASAP7_75t_L g1833 ( 
.A(n_1813),
.B(n_1465),
.C(n_1637),
.D(n_1468),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1816),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1815),
.Y(n_1835)
);

OAI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1834),
.A2(n_1811),
.B1(n_1646),
.B2(n_1600),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1827),
.Y(n_1837)
);

AO22x2_ASAP7_75t_L g1838 ( 
.A1(n_1835),
.A2(n_1825),
.B1(n_1828),
.B2(n_1822),
.Y(n_1838)
);

XOR2xp5_ASAP7_75t_L g1839 ( 
.A(n_1827),
.B(n_245),
.Y(n_1839)
);

XNOR2x2_ASAP7_75t_L g1840 ( 
.A(n_1824),
.B(n_1460),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1829),
.Y(n_1841)
);

NOR4xp75_ASAP7_75t_L g1842 ( 
.A(n_1826),
.B(n_251),
.C(n_252),
.D(n_253),
.Y(n_1842)
);

XOR2xp5_ASAP7_75t_L g1843 ( 
.A(n_1832),
.B(n_257),
.Y(n_1843)
);

XOR2xp5_ASAP7_75t_L g1844 ( 
.A(n_1831),
.B(n_261),
.Y(n_1844)
);

OAI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1838),
.A2(n_1830),
.B1(n_1823),
.B2(n_1833),
.Y(n_1845)
);

NOR3xp33_ASAP7_75t_L g1846 ( 
.A(n_1837),
.B(n_263),
.C(n_264),
.Y(n_1846)
);

NAND5xp2_ASAP7_75t_L g1847 ( 
.A(n_1839),
.B(n_1584),
.C(n_1540),
.D(n_1564),
.E(n_273),
.Y(n_1847)
);

OAI221xp5_ASAP7_75t_L g1848 ( 
.A1(n_1843),
.A2(n_1610),
.B1(n_1646),
.B2(n_1626),
.C(n_1633),
.Y(n_1848)
);

NAND5xp2_ASAP7_75t_L g1849 ( 
.A(n_1838),
.B(n_266),
.C(n_267),
.D(n_271),
.E(n_276),
.Y(n_1849)
);

AOI221xp5_ASAP7_75t_L g1850 ( 
.A1(n_1844),
.A2(n_1626),
.B1(n_1639),
.B2(n_1633),
.C(n_1443),
.Y(n_1850)
);

OAI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1845),
.A2(n_1841),
.B1(n_1836),
.B2(n_1840),
.Y(n_1851)
);

OAI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1848),
.A2(n_1842),
.B1(n_1646),
.B2(n_1610),
.Y(n_1852)
);

OAI21xp33_ASAP7_75t_L g1853 ( 
.A1(n_1849),
.A2(n_1646),
.B(n_1610),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1847),
.Y(n_1854)
);

OAI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1846),
.A2(n_1646),
.B1(n_1610),
.B2(n_1639),
.Y(n_1855)
);

OAI22xp5_ASAP7_75t_SL g1856 ( 
.A1(n_1850),
.A2(n_1637),
.B1(n_1635),
.B2(n_1625),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1854),
.Y(n_1857)
);

AOI21xp5_ASAP7_75t_L g1858 ( 
.A1(n_1851),
.A2(n_1581),
.B(n_1469),
.Y(n_1858)
);

AOI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1852),
.A2(n_1632),
.B1(n_1637),
.B2(n_1658),
.Y(n_1859)
);

AO22x1_ASAP7_75t_L g1860 ( 
.A1(n_1855),
.A2(n_1853),
.B1(n_1856),
.B2(n_1667),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1857),
.A2(n_277),
.B(n_279),
.Y(n_1861)
);

AOI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1860),
.A2(n_282),
.B(n_283),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_SL g1863 ( 
.A(n_1859),
.B(n_1667),
.Y(n_1863)
);

OAI21xp5_ASAP7_75t_L g1864 ( 
.A1(n_1858),
.A2(n_1472),
.B(n_1668),
.Y(n_1864)
);

AOI22xp33_ASAP7_75t_L g1865 ( 
.A1(n_1862),
.A2(n_1863),
.B1(n_1861),
.B2(n_1864),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1862),
.B(n_284),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1862),
.B(n_285),
.Y(n_1867)
);

AOI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1866),
.A2(n_1668),
.B1(n_1637),
.B2(n_1635),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1867),
.Y(n_1869)
);

AOI221xp5_ASAP7_75t_L g1870 ( 
.A1(n_1869),
.A2(n_1865),
.B1(n_1629),
.B2(n_1627),
.C(n_1637),
.Y(n_1870)
);

AOI211xp5_ASAP7_75t_L g1871 ( 
.A1(n_1870),
.A2(n_1868),
.B(n_1627),
.C(n_289),
.Y(n_1871)
);


endmodule