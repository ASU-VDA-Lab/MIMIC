module fake_jpeg_26589_n_76 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_76);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_76;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_75;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_70;
wire n_15;
wire n_66;

INVx1_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx10_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_20),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_0),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_22),
.Y(n_24)
);

NOR2x1_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_17),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_13),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_14),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_30),
.B(n_33),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_8),
.B(n_10),
.C(n_13),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_16),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_15),
.B(n_14),
.C(n_10),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_15),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_36),
.B1(n_38),
.B2(n_9),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_16),
.B1(n_9),
.B2(n_8),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_18),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_39),
.Y(n_49)
);

OAI21xp33_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_21),
.B(n_16),
.Y(n_41)
);

XOR2x1_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_42),
.B(n_44),
.Y(n_52)
);

MAJx2_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_18),
.C(n_19),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_SL g57 ( 
.A(n_46),
.B(n_19),
.Y(n_57)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_49),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_54),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_55),
.Y(n_61)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_19),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_58),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_57),
.C(n_55),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_63),
.B(n_66),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_61),
.B(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_60),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_61),
.A2(n_52),
.B1(n_47),
.B2(n_46),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_68),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_40),
.B(n_45),
.Y(n_68)
);

AOI211xp5_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_63),
.B(n_45),
.C(n_3),
.Y(n_71)
);

BUFx24_ASAP7_75t_SL g73 ( 
.A(n_71),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_48),
.Y(n_72)
);

AOI322xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_73),
.A3(n_22),
.B1(n_4),
.B2(n_6),
.C1(n_2),
.C2(n_1),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_74),
.A2(n_1),
.B(n_21),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_1),
.Y(n_76)
);


endmodule