module fake_jpeg_17032_n_165 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_165);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_SL g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_41),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_13),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_33),
.A2(n_48),
.B1(n_22),
.B2(n_26),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_2),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_34),
.B(n_35),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_6),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_36),
.B(n_39),
.Y(n_61)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_6),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_6),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_20),
.B(n_9),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_47),
.Y(n_65)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_23),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_20),
.B(n_11),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_49),
.B(n_25),
.Y(n_54)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_51),
.Y(n_67)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_22),
.A2(n_12),
.B1(n_29),
.B2(n_21),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_52),
.A2(n_26),
.B1(n_18),
.B2(n_21),
.Y(n_58)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_54),
.B(n_66),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_58),
.A2(n_70),
.B1(n_56),
.B2(n_65),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_29),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_62),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_27),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_35),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_69),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_19),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_47),
.A2(n_31),
.B1(n_30),
.B2(n_12),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_34),
.B(n_31),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_45),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_39),
.B(n_30),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_73),
.B(n_77),
.Y(n_89)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_79),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_40),
.C(n_46),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_37),
.C(n_53),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_43),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_51),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_32),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_82),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_41),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_76),
.A2(n_45),
.B1(n_53),
.B2(n_41),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_88),
.Y(n_105)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_87),
.Y(n_110)
);

BUFx12_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_55),
.B(n_61),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_93),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_55),
.B(n_61),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_66),
.A2(n_60),
.B1(n_59),
.B2(n_71),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_95),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_102),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_77),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_103),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_78),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_58),
.B(n_63),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_SL g117 ( 
.A(n_104),
.B(n_56),
.C(n_64),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_98),
.A2(n_62),
.B(n_70),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_72),
.B(n_78),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_84),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_112),
.Y(n_133)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_92),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_113),
.B(n_116),
.Y(n_123)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_117),
.A2(n_102),
.B1(n_96),
.B2(n_95),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_120),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_64),
.C(n_72),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_119),
.B(n_89),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_86),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_111),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_SL g124 ( 
.A1(n_117),
.A2(n_104),
.B(n_83),
.C(n_98),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_128),
.B1(n_135),
.B2(n_109),
.Y(n_144)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_107),
.A2(n_98),
.B1(n_100),
.B2(n_99),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_127),
.A2(n_130),
.B1(n_131),
.B2(n_115),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_119),
.C(n_115),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_101),
.B1(n_97),
.B2(n_91),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_116),
.A2(n_97),
.B1(n_74),
.B2(n_80),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_134),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_110),
.A2(n_86),
.B(n_78),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_105),
.A2(n_80),
.B1(n_88),
.B2(n_108),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_122),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_137),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_130),
.B(n_114),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_138),
.A2(n_140),
.B(n_144),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_134),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_106),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_110),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_127),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_123),
.B(n_114),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_145),
.A2(n_113),
.B1(n_112),
.B2(n_141),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_147),
.C(n_151),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_148),
.A2(n_133),
.B1(n_144),
.B2(n_126),
.Y(n_154)
);

MAJx2_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_124),
.C(n_132),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_141),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_152),
.A2(n_128),
.B(n_143),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_150),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_153),
.A2(n_155),
.B(n_157),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_137),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_152),
.A2(n_143),
.B(n_124),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_156),
.A2(n_151),
.B(n_149),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_159),
.A2(n_160),
.B(n_124),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_162),
.C(n_120),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_158),
.Y(n_162)
);

OAI321xp33_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_139),
.A3(n_146),
.B1(n_156),
.B2(n_109),
.C(n_106),
.Y(n_163)
);

AOI221xp5_ASAP7_75t_L g165 ( 
.A1(n_163),
.A2(n_164),
.B1(n_121),
.B2(n_118),
.C(n_88),
.Y(n_165)
);


endmodule