module real_jpeg_6546_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_0),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_0),
.B(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_0),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_0),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_0),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_1),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_1),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_1),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_1),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_1),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_1),
.B(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_1),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_1),
.B(n_377),
.Y(n_376)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_3),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_3),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_4),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_4),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_4),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_4),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_4),
.B(n_210),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_4),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_4),
.B(n_269),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_5),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_5),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_SL g50 ( 
.A(n_5),
.B(n_51),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_5),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_5),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_5),
.B(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_5),
.Y(n_145)
);

AND2x2_ASAP7_75t_SL g174 ( 
.A(n_5),
.B(n_175),
.Y(n_174)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_7),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_8),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_8),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_8),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_8),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_8),
.B(n_239),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_9),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_9),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_9),
.B(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_9),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_9),
.B(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_9),
.B(n_372),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_9),
.B(n_402),
.Y(n_401)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_11),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_11),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g189 ( 
.A(n_11),
.Y(n_189)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_11),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_11),
.Y(n_251)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_12),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_12),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_12),
.Y(n_148)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_12),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_13),
.B(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_13),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_13),
.B(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_13),
.B(n_259),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_13),
.B(n_385),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_14),
.Y(n_102)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_14),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_14),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_15),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_15),
.B(n_127),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_15),
.B(n_272),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_15),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_15),
.B(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_15),
.B(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_196),
.B1(n_449),
.B2(n_450),
.Y(n_17)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_18),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_195),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_164),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_21),
.B(n_164),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_96),
.C(n_135),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_22),
.B(n_332),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_66),
.C(n_85),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_23),
.B(n_326),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_40),
.C(n_55),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_24),
.B(n_283),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_36),
.B2(n_39),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_31),
.B2(n_35),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_27),
.A2(n_28),
.B1(n_147),
.B2(n_149),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_27),
.A2(n_28),
.B1(n_341),
.B2(n_342),
.Y(n_378)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_28),
.B(n_31),
.C(n_36),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_28),
.B(n_144),
.C(n_147),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_28),
.B(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_30),
.Y(n_241)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_30),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_30),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_31),
.B(n_225),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_31),
.A2(n_35),
.B1(n_225),
.B2(n_226),
.Y(n_312)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_34),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_36),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_36),
.A2(n_39),
.B1(n_191),
.B2(n_193),
.Y(n_190)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_37),
.Y(n_260)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_38),
.Y(n_131)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_38),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_40),
.B(n_55),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_45),
.C(n_50),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_41),
.B(n_50),
.Y(n_277)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_43),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_44),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g305 ( 
.A(n_44),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_45),
.B(n_277),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_50),
.A2(n_129),
.B1(n_132),
.B2(n_133),
.Y(n_128)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_50),
.Y(n_133)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_53),
.Y(n_217)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_54),
.Y(n_354)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_54),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_56),
.Y(n_142)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_58),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_58),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_64),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_60),
.B(n_64),
.C(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_62),
.B(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_62),
.Y(n_348)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_63),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_66),
.B(n_85),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_79),
.C(n_82),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_68),
.B(n_289),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.C(n_77),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_69),
.A2(n_70),
.B1(n_77),
.B2(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_70),
.B(n_106),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_70),
.B(n_106),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_72),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_72),
.Y(n_231)
);

OR2x2_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OR2x2_ASAP7_75t_SL g99 ( 
.A(n_76),
.B(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_111),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_76),
.B(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_77),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_79),
.B(n_82),
.Y(n_289)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_80),
.Y(n_171)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_81),
.B(n_248),
.Y(n_306)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_95),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_92),
.B2(n_94),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_88),
.B(n_92),
.C(n_95),
.Y(n_154)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_92),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_92),
.A2(n_94),
.B1(n_160),
.B2(n_163),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_94),
.B(n_156),
.C(n_163),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_96),
.B(n_135),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_114),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_97),
.B(n_115),
.C(n_124),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_103),
.B2(n_104),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_98),
.A2(n_99),
.B1(n_174),
.B2(n_177),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_98),
.A2(n_99),
.B1(n_218),
.B2(n_299),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_99),
.B(n_106),
.C(n_110),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_99),
.B(n_216),
.C(n_218),
.Y(n_215)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_102),
.Y(n_246)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_110),
.B2(n_113),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_105),
.A2(n_106),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_116),
.C(n_120),
.Y(n_115)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_109),
.Y(n_374)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_110),
.Y(n_113)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_124),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_116),
.A2(n_117),
.B1(n_120),
.B2(n_121),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_128),
.B2(n_134),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_126),
.B(n_129),
.C(n_133),
.Y(n_181)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_128),
.Y(n_134)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_152),
.B2(n_153),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_154),
.C(n_155),
.Y(n_165)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.C(n_143),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_138),
.B(n_141),
.Y(n_324)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_143),
.B(n_324),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_146),
.B1(n_150),
.B2(n_151),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_144),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_144),
.A2(n_150),
.B1(n_258),
.B2(n_261),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_144),
.B(n_254),
.C(n_258),
.Y(n_275)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_146),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_147),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

AO22x1_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_160),
.Y(n_163)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx24_ASAP7_75t_SL g452 ( 
.A(n_164),
.Y(n_452)
);

FAx1_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_166),
.CI(n_182),
.CON(n_164),
.SN(n_164)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_178),
.B2(n_179),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_169),
.A2(n_170),
.B1(n_205),
.B2(n_208),
.Y(n_204)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_170),
.B(n_205),
.C(n_209),
.Y(n_278)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_174),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_175),
.Y(n_256)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_194),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_190),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_191),
.Y(n_193)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_196),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_333),
.Y(n_196)
);

O2A1O1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_319),
.B(n_328),
.C(n_329),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_290),
.B(n_318),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_199),
.B(n_447),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_279),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_200),
.B(n_279),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_252),
.C(n_273),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_201),
.B(n_317),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_229),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_202),
.B(n_230),
.C(n_235),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_215),
.C(n_223),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_203),
.B(n_314),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_209),
.Y(n_203)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_205),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx8_ASAP7_75t_L g345 ( 
.A(n_214),
.Y(n_345)
);

BUFx5_ASAP7_75t_L g408 ( 
.A(n_214),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_215),
.A2(n_223),
.B1(n_224),
.B2(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_215),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_216),
.B(n_298),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_218),
.Y(n_299)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_222),
.Y(n_311)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_235),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_242),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_236),
.A2(n_237),
.B(n_238),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_236),
.B(n_243),
.C(n_247),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_240),
.Y(n_269)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_247),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

INVx8_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_252),
.B(n_273),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_262),
.C(n_264),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_253),
.A2(n_262),
.B1(n_263),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_253),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_255),
.B(n_407),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_255),
.B(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_258),
.Y(n_261)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_264),
.B(n_294),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.C(n_270),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_265),
.A2(n_266),
.B1(n_436),
.B2(n_437),
.Y(n_435)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_267),
.A2(n_268),
.B1(n_270),
.B2(n_271),
.Y(n_437)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_278),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_276),
.C(n_278),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_280),
.B(n_282),
.C(n_284),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_285),
.B(n_287),
.C(n_288),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_316),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_291),
.B(n_316),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_296),
.C(n_313),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_292),
.A2(n_293),
.B1(n_441),
.B2(n_442),
.Y(n_440)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_296),
.B(n_313),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_300),
.C(n_312),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_297),
.B(n_431),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_300),
.B(n_312),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_306),
.C(n_307),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_301),
.A2(n_302),
.B1(n_307),
.B2(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx6_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_306),
.B(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_307),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_308),
.B(n_353),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_308),
.B(n_410),
.Y(n_409)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx8_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_320),
.B(n_330),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_322),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_331),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_322),
.B(n_331),
.Y(n_448)
);

FAx1_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_325),
.CI(n_327),
.CON(n_322),
.SN(n_322)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

OAI31xp33_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_445),
.A3(n_446),
.B(n_448),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_439),
.B(n_444),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_336),
.A2(n_426),
.B(n_438),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_379),
.B(n_425),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_338),
.B(n_365),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_338),
.B(n_365),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_350),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_339),
.B(n_351),
.C(n_362),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_346),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_340),
.B(n_347),
.C(n_349),
.Y(n_434)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx8_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_349),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_362),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_355),
.C(n_357),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_352),
.B(n_367),
.Y(n_366)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_355),
.A2(n_356),
.B1(n_357),
.B2(n_358),
.Y(n_367)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx8_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

BUFx5_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_368),
.C(n_378),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_366),
.B(n_422),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_368),
.A2(n_369),
.B1(n_378),
.B2(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_375),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_370),
.A2(n_371),
.B1(n_375),
.B2(n_376),
.Y(n_392)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx5_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_378),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_380),
.A2(n_419),
.B(n_424),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_404),
.B(n_418),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_382),
.B(n_393),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_382),
.B(n_393),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_392),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_390),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_384),
.B(n_390),
.C(n_392),
.Y(n_420)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx5_ASAP7_75t_SL g386 ( 
.A(n_387),
.Y(n_386)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_400),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_394),
.A2(n_395),
.B1(n_400),
.B2(n_401),
.Y(n_416)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx6_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx8_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_412),
.B(n_417),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_409),
.Y(n_405)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_416),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_413),
.B(n_416),
.Y(n_417)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_421),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_420),
.B(n_421),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_428),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_427),
.B(n_428),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_429),
.A2(n_430),
.B1(n_432),
.B2(n_433),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_434),
.C(n_435),
.Y(n_443)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_435),
.Y(n_433)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_440),
.B(n_443),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_440),
.B(n_443),
.Y(n_444)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_441),
.Y(n_442)
);


endmodule