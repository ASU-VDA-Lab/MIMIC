module fake_jpeg_1876_n_275 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_275);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_275;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g113 ( 
.A(n_43),
.Y(n_113)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx4f_ASAP7_75t_SL g97 ( 
.A(n_45),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_46),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_33),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_48),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_23),
.B(n_11),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_52),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_33),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_32),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_53),
.B(n_62),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_29),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_30),
.B(n_1),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_69),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_29),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_25),
.B(n_1),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_70),
.B(n_16),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_37),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_74),
.B(n_91),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_26),
.B1(n_35),
.B2(n_28),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_79),
.A2(n_9),
.B1(n_15),
.B2(n_110),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_48),
.B(n_37),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_82),
.B(n_87),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_31),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_84),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_53),
.B(n_35),
.Y(n_87)
);

BUFx12_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_90),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_41),
.B(n_28),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_47),
.B(n_39),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_93),
.B(n_78),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_65),
.A2(n_27),
.B1(n_39),
.B2(n_17),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_95),
.Y(n_124)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_27),
.C(n_17),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_101),
.C(n_111),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_64),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_101),
.B(n_117),
.Y(n_148)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_45),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_111),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_L g118 ( 
.A1(n_45),
.A2(n_16),
.B(n_5),
.Y(n_118)
);

OR2x2_ASAP7_75t_SL g135 ( 
.A(n_118),
.B(n_3),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_117),
.B(n_112),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_119),
.B(n_125),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_79),
.A2(n_24),
.B1(n_5),
.B2(n_7),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_120),
.A2(n_130),
.B1(n_138),
.B2(n_146),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_99),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_106),
.A2(n_24),
.B1(n_5),
.B2(n_8),
.Y(n_130)
);

OR2x4_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_64),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_131),
.A2(n_127),
.B(n_136),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_133),
.Y(n_160)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_135),
.Y(n_175)
);

O2A1O1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_99),
.A2(n_50),
.B(n_8),
.C(n_10),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_82),
.A2(n_9),
.B1(n_10),
.B2(n_15),
.Y(n_138)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_92),
.Y(n_139)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_140),
.A2(n_147),
.B1(n_124),
.B2(n_142),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_103),
.Y(n_155)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_97),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_145),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_94),
.B(n_96),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_102),
.A2(n_77),
.B1(n_80),
.B2(n_113),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_109),
.A2(n_104),
.B1(n_85),
.B2(n_81),
.Y(n_147)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_88),
.B(n_113),
.C(n_94),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_75),
.C(n_86),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_162),
.C(n_168),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_156),
.B(n_174),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_97),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_170),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_90),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_108),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_178),
.Y(n_190)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_169),
.Y(n_193)
);

NOR2x1p5_ASAP7_75t_SL g170 ( 
.A(n_131),
.B(n_75),
.Y(n_170)
);

AND2x2_ASAP7_75t_SL g171 ( 
.A(n_141),
.B(n_108),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_180),
.Y(n_188)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_133),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_123),
.B(n_135),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_177),
.B(n_121),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_129),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_182),
.B(n_196),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_170),
.A2(n_139),
.B(n_126),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_184),
.A2(n_163),
.B(n_180),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_128),
.C(n_137),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_191),
.C(n_197),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_147),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_134),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_192),
.B(n_194),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_149),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_158),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_203),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_177),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_155),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_154),
.B(n_168),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_198),
.B(n_199),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_159),
.B(n_179),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_157),
.Y(n_201)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_164),
.Y(n_202)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_175),
.B(n_164),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_205),
.A2(n_193),
.B(n_200),
.Y(n_234)
);

AO22x1_ASAP7_75t_L g206 ( 
.A1(n_187),
.A2(n_163),
.B1(n_176),
.B2(n_171),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_210),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_181),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_204),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_172),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_185),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_161),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_161),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_219),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_188),
.A2(n_172),
.B1(n_160),
.B2(n_166),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_220),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_187),
.A2(n_191),
.B1(n_189),
.B2(n_190),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_221),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_212),
.A2(n_193),
.B1(n_201),
.B2(n_189),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_222),
.A2(n_232),
.B1(n_219),
.B2(n_220),
.Y(n_245)
);

INVxp33_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_205),
.A2(n_184),
.B(n_197),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_227),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_215),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_L g228 ( 
.A1(n_221),
.A2(n_211),
.B(n_199),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_228),
.B(n_234),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_214),
.C(n_186),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_215),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_216),
.Y(n_241)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_231),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_236),
.A2(n_239),
.B1(n_242),
.B2(n_245),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_208),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_214),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_223),
.A2(n_218),
.B1(n_210),
.B2(n_206),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_225),
.C(n_226),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_241),
.Y(n_248)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_231),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_244),
.A2(n_232),
.B1(n_206),
.B2(n_235),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_247),
.B(n_253),
.Y(n_256)
);

NOR2xp67_ASAP7_75t_SL g257 ( 
.A(n_249),
.B(n_241),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_240),
.C(n_237),
.Y(n_255)
);

NAND2xp67_ASAP7_75t_SL g251 ( 
.A(n_243),
.B(n_226),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_251),
.A2(n_252),
.B(n_246),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_239),
.A2(n_238),
.B1(n_235),
.B2(n_234),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_183),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_254),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_257),
.C(n_248),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_250),
.C(n_229),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_258),
.B(n_259),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_229),
.C(n_227),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_233),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_242),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_256),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_251),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_213),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_266),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_236),
.C(n_217),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_267),
.A2(n_268),
.B(n_264),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_264),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_270),
.B(n_271),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_202),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_272),
.B(n_166),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_273),
.Y(n_275)
);


endmodule