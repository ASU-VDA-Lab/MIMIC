module fake_netlist_5_68_n_2195 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_2195);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_2195;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_2142;
wire n_320;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_223;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2140;
wire n_1819;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_944;
wire n_345;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_561;
wire n_1319;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_604;
wire n_368;
wire n_433;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2137;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_2176;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_2131;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_2153;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2080;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1834;
wire n_1659;
wire n_2097;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1912;
wire n_1771;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_2148;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_2136;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_994;
wire n_386;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1478;
wire n_1339;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2183;
wire n_328;
wire n_1250;
wire n_2173;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1495;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_2135;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

BUFx2_ASAP7_75t_L g222 ( 
.A(n_164),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_129),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_168),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_38),
.Y(n_225)
);

BUFx5_ASAP7_75t_L g226 ( 
.A(n_44),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_68),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_55),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_100),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_77),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_143),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_30),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_204),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_16),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_216),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_169),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_22),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_5),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_99),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_179),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_102),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_149),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_75),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_119),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_174),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_155),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_52),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_91),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_131),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_2),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_153),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_162),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_2),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_66),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_118),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_11),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_181),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_135),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_74),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_208),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_171),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_195),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_127),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_50),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_180),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_141),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_113),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_150),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_110),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_163),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_194),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_193),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_46),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_128),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_51),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_77),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_23),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_75),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_17),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_85),
.Y(n_281)
);

BUFx10_ASAP7_75t_L g282 ( 
.A(n_176),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_157),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_38),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_188),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_62),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_8),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_103),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_25),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_151),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_44),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_42),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_24),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_66),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_4),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_39),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_68),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_147),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_94),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_0),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_142),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_133),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_198),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_137),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_124),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_31),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_39),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_189),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_52),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_45),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_83),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_8),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_161),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_82),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_202),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_154),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_25),
.Y(n_317)
);

BUFx5_ASAP7_75t_L g318 ( 
.A(n_210),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_60),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_64),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_71),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_73),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_112),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_191),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_82),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_200),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_160),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_72),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_104),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_173),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_185),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_108),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_156),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_43),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_190),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_47),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_166),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_14),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_41),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_36),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_56),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_138),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_40),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_64),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_136),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_54),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_196),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_114),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_47),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_183),
.Y(n_350)
);

BUFx5_ASAP7_75t_L g351 ( 
.A(n_85),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_5),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_177),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_79),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_69),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_41),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_90),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_48),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_172),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_148),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_159),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_79),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_46),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_53),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_212),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_205),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_74),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_71),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_201),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_132),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_15),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_197),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_90),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_123),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_51),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_69),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_16),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_17),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_4),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_89),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_192),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_144),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_88),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_49),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_40),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_49),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_36),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_186),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_199),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_117),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_48),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_42),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_93),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_33),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_30),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_122),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_182),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_50),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_55),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_62),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_101),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_89),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_54),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_31),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_19),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_96),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_105),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_84),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_6),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_0),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_9),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_45),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_158),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_18),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_78),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_67),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_165),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_111),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_187),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_6),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_211),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_218),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_24),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_86),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_139),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_213),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_98),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_125),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_35),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_86),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_121),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_22),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_37),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_57),
.Y(n_434)
);

INVx2_ASAP7_75t_SL g435 ( 
.A(n_57),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_11),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_303),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_314),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_409),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_305),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_332),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g442 ( 
.A(n_227),
.B(n_233),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_226),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_314),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_409),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_319),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_319),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_396),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_422),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_434),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_226),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_268),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_226),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_226),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_226),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_434),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_268),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_225),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_228),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_L g460 ( 
.A(n_286),
.B(n_1),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_239),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_231),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_248),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_251),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_287),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_222),
.B(n_1),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_384),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_254),
.Y(n_468)
);

NOR2xp67_ASAP7_75t_L g469 ( 
.A(n_286),
.B(n_3),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_222),
.B(n_3),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_255),
.Y(n_471)
);

INVxp33_ASAP7_75t_SL g472 ( 
.A(n_257),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_260),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_226),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_279),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_226),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_308),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_226),
.B(n_7),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_308),
.Y(n_479)
);

NOR2xp67_ASAP7_75t_L g480 ( 
.A(n_286),
.B(n_7),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_390),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_226),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_224),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_351),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_351),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_351),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_281),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_235),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_291),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_390),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_267),
.B(n_9),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_351),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_351),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_417),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_223),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_229),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_292),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_351),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_293),
.Y(n_499)
);

NOR2xp67_ASAP7_75t_L g500 ( 
.A(n_286),
.B(n_10),
.Y(n_500)
);

NOR2xp67_ASAP7_75t_L g501 ( 
.A(n_238),
.B(n_10),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_R g502 ( 
.A(n_234),
.B(n_236),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_351),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_351),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_296),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_351),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_232),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_232),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_237),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_297),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_237),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_267),
.B(n_12),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_392),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_235),
.Y(n_514)
);

INVxp67_ASAP7_75t_SL g515 ( 
.A(n_298),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_300),
.Y(n_516)
);

CKINVDCx14_ASAP7_75t_R g517 ( 
.A(n_249),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_235),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_240),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_230),
.B(n_299),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_306),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_235),
.Y(n_522)
);

NOR2xp67_ASAP7_75t_L g523 ( 
.A(n_238),
.B(n_12),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_241),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_241),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_230),
.B(n_13),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_235),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_307),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_250),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_250),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_311),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_320),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_243),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_252),
.Y(n_534)
);

CKINVDCx16_ASAP7_75t_R g535 ( 
.A(n_249),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_252),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_253),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_245),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_246),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_253),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_256),
.Y(n_541)
);

INVxp33_ASAP7_75t_L g542 ( 
.A(n_227),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_235),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_417),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_430),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_256),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_322),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_325),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_392),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_247),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_328),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_258),
.Y(n_552)
);

CKINVDCx16_ASAP7_75t_R g553 ( 
.A(n_249),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_494),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_488),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_488),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_535),
.B(n_249),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_460),
.B(n_348),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_488),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_514),
.B(n_518),
.Y(n_560)
);

NOR2x1_ASAP7_75t_L g561 ( 
.A(n_520),
.B(n_230),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_456),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_514),
.Y(n_563)
);

OAI21x1_ASAP7_75t_L g564 ( 
.A1(n_451),
.A2(n_361),
.B(n_326),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_469),
.B(n_365),
.Y(n_565)
);

BUFx2_ASAP7_75t_L g566 ( 
.A(n_438),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_494),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_518),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_438),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_494),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_522),
.B(n_430),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_494),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_494),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_522),
.B(n_430),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_527),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_544),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_527),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_444),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_544),
.Y(n_579)
);

BUFx2_ASAP7_75t_L g580 ( 
.A(n_444),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_544),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_543),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_543),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_545),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_544),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_544),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_545),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_453),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_480),
.B(n_361),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_453),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_454),
.Y(n_591)
);

CKINVDCx6p67_ASAP7_75t_R g592 ( 
.A(n_479),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_513),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_454),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_455),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_443),
.B(n_430),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_487),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_455),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_451),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_485),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_474),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_476),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_446),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_482),
.B(n_430),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_484),
.B(n_430),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_513),
.B(n_392),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_486),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g608 ( 
.A(n_551),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_492),
.B(n_259),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_485),
.Y(n_610)
);

CKINVDCx8_ASAP7_75t_R g611 ( 
.A(n_553),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_502),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_493),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_SL g614 ( 
.A(n_466),
.B(n_265),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_549),
.B(n_284),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_498),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_503),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_504),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_472),
.B(n_282),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_506),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_442),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_442),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_483),
.B(n_242),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_478),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_507),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_508),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_509),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_511),
.Y(n_628)
);

OAI21x1_ASAP7_75t_L g629 ( 
.A1(n_526),
.A2(n_326),
.B(n_299),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_524),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_525),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_529),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_446),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_549),
.B(n_284),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_530),
.Y(n_635)
);

INVxp67_ASAP7_75t_L g636 ( 
.A(n_462),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_515),
.B(n_264),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_534),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_536),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_537),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_540),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_541),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_546),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_500),
.Y(n_644)
);

BUFx10_ASAP7_75t_L g645 ( 
.A(n_612),
.Y(n_645)
);

AO22x2_ASAP7_75t_L g646 ( 
.A1(n_624),
.A2(n_512),
.B1(n_439),
.B2(n_445),
.Y(n_646)
);

BUFx6f_ASAP7_75t_SL g647 ( 
.A(n_558),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_554),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_554),
.Y(n_649)
);

INVx5_ASAP7_75t_L g650 ( 
.A(n_613),
.Y(n_650)
);

AOI21x1_ASAP7_75t_L g651 ( 
.A1(n_596),
.A2(n_326),
.B(n_299),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_601),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_588),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_623),
.B(n_458),
.Y(n_654)
);

INVx4_ASAP7_75t_L g655 ( 
.A(n_613),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_624),
.B(n_517),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_601),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_588),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_592),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_599),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_599),
.Y(n_661)
);

BUFx4f_ASAP7_75t_L g662 ( 
.A(n_613),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_590),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_624),
.A2(n_491),
.B1(n_470),
.B2(n_336),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_614),
.B(n_495),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_614),
.B(n_496),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_637),
.B(n_458),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_644),
.B(n_542),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_599),
.Y(n_669)
);

INVx4_ASAP7_75t_L g670 ( 
.A(n_613),
.Y(n_670)
);

NAND2xp33_ASAP7_75t_R g671 ( 
.A(n_566),
.B(n_447),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_554),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_597),
.B(n_459),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_600),
.Y(n_674)
);

INVx4_ASAP7_75t_L g675 ( 
.A(n_613),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_554),
.Y(n_676)
);

AO22x2_ASAP7_75t_L g677 ( 
.A1(n_557),
.A2(n_435),
.B1(n_349),
.B2(n_375),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_600),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_600),
.Y(n_679)
);

BUFx4f_ASAP7_75t_L g680 ( 
.A(n_613),
.Y(n_680)
);

NOR2x1p5_ASAP7_75t_L g681 ( 
.A(n_592),
.B(n_447),
.Y(n_681)
);

XNOR2xp5_ASAP7_75t_L g682 ( 
.A(n_619),
.B(n_437),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_610),
.Y(n_683)
);

INVx1_ASAP7_75t_SL g684 ( 
.A(n_593),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_606),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_597),
.B(n_519),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_610),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_610),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_590),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_591),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_563),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_563),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_608),
.B(n_533),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_608),
.B(n_459),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_591),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_568),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_568),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_602),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_594),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_621),
.B(n_538),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_594),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_595),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_595),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_575),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_598),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_575),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_621),
.A2(n_539),
.B1(n_552),
.B2(n_550),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_622),
.B(n_461),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_593),
.B(n_450),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_606),
.Y(n_710)
);

AND2x6_ASAP7_75t_L g711 ( 
.A(n_561),
.B(n_417),
.Y(n_711)
);

OAI22xp33_ASAP7_75t_L g712 ( 
.A1(n_562),
.A2(n_309),
.B1(n_312),
.B2(n_276),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_609),
.B(n_461),
.Y(n_713)
);

OAI22xp33_ASAP7_75t_L g714 ( 
.A1(n_562),
.A2(n_405),
.B1(n_467),
.B2(n_465),
.Y(n_714)
);

INVx5_ASAP7_75t_L g715 ( 
.A(n_613),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_577),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_577),
.Y(n_717)
);

BUFx6f_ASAP7_75t_SL g718 ( 
.A(n_558),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_582),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_609),
.B(n_463),
.Y(n_720)
);

INVxp67_ASAP7_75t_SL g721 ( 
.A(n_596),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_554),
.Y(n_722)
);

BUFx10_ASAP7_75t_L g723 ( 
.A(n_558),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_622),
.B(n_463),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_598),
.Y(n_725)
);

INVxp33_ASAP7_75t_L g726 ( 
.A(n_615),
.Y(n_726)
);

NAND2xp33_ASAP7_75t_L g727 ( 
.A(n_644),
.B(n_464),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_602),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_SL g729 ( 
.A(n_611),
.B(n_282),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_607),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_615),
.Y(n_731)
);

AND2x6_ASAP7_75t_L g732 ( 
.A(n_561),
.B(n_417),
.Y(n_732)
);

AOI22xp5_ASAP7_75t_L g733 ( 
.A1(n_634),
.A2(n_321),
.B1(n_340),
.B2(n_310),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_582),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_583),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_607),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_616),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_616),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_558),
.B(n_464),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_617),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_583),
.Y(n_741)
);

OAI22xp33_ASAP7_75t_L g742 ( 
.A1(n_636),
.A2(n_450),
.B1(n_523),
.B2(n_501),
.Y(n_742)
);

INVx5_ASAP7_75t_L g743 ( 
.A(n_618),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_617),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_584),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_584),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_565),
.B(n_468),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_634),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_620),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_565),
.B(n_468),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_620),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_587),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_628),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_554),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_628),
.Y(n_755)
);

INVxp33_ASAP7_75t_SL g756 ( 
.A(n_569),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_587),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_555),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_628),
.Y(n_759)
);

OR2x6_ASAP7_75t_L g760 ( 
.A(n_565),
.B(n_629),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_554),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_570),
.Y(n_762)
);

BUFx10_ASAP7_75t_L g763 ( 
.A(n_565),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_570),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_636),
.B(n_471),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_570),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_628),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_555),
.Y(n_768)
);

OR2x2_ASAP7_75t_L g769 ( 
.A(n_566),
.B(n_471),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_570),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_556),
.Y(n_771)
);

OR2x6_ASAP7_75t_L g772 ( 
.A(n_629),
.B(n_262),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_556),
.Y(n_773)
);

HB1xp67_ASAP7_75t_L g774 ( 
.A(n_633),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_SL g775 ( 
.A(n_611),
.B(n_282),
.Y(n_775)
);

AND3x2_ASAP7_75t_L g776 ( 
.A(n_578),
.B(n_370),
.C(n_349),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_589),
.A2(n_336),
.B1(n_375),
.B2(n_349),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_589),
.B(n_473),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_635),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_559),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_589),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_589),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_626),
.A2(n_336),
.B1(n_415),
.B2(n_375),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_559),
.Y(n_784)
);

INVx6_ASAP7_75t_L g785 ( 
.A(n_618),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_635),
.B(n_473),
.Y(n_786)
);

INVx4_ASAP7_75t_L g787 ( 
.A(n_618),
.Y(n_787)
);

INVx4_ASAP7_75t_L g788 ( 
.A(n_618),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_567),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_564),
.B(n_262),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_635),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_626),
.B(n_475),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_611),
.A2(n_489),
.B1(n_497),
.B2(n_475),
.Y(n_793)
);

BUFx2_ASAP7_75t_L g794 ( 
.A(n_578),
.Y(n_794)
);

AO22x2_ASAP7_75t_L g795 ( 
.A1(n_627),
.A2(n_435),
.B1(n_415),
.B2(n_244),
.Y(n_795)
);

AND2x6_ASAP7_75t_L g796 ( 
.A(n_618),
.B(n_417),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_635),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_618),
.B(n_489),
.Y(n_798)
);

INVx5_ASAP7_75t_L g799 ( 
.A(n_618),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_L g800 ( 
.A1(n_580),
.A2(n_499),
.B1(n_505),
.B2(n_497),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_713),
.B(n_452),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_781),
.B(n_630),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_790),
.A2(n_629),
.B1(n_313),
.B2(n_315),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_720),
.B(n_457),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_781),
.B(n_630),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_685),
.B(n_782),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_790),
.A2(n_313),
.B1(n_315),
.B2(n_288),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_782),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_721),
.B(n_630),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_668),
.Y(n_810)
);

OAI22xp33_ASAP7_75t_L g811 ( 
.A1(n_729),
.A2(n_592),
.B1(n_481),
.B2(n_490),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_652),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_723),
.B(n_417),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_691),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_653),
.B(n_630),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_685),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_723),
.B(n_580),
.Y(n_817)
);

NAND2xp33_ASAP7_75t_L g818 ( 
.A(n_711),
.B(n_318),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_691),
.Y(n_819)
);

AOI22xp5_ASAP7_75t_L g820 ( 
.A1(n_731),
.A2(n_477),
.B1(n_603),
.B2(n_441),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_728),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_726),
.B(n_603),
.Y(n_822)
);

NOR2x1p5_ASAP7_75t_L g823 ( 
.A(n_659),
.B(n_499),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_668),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_728),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_723),
.B(n_318),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_730),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_730),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_692),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_736),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_692),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_765),
.B(n_505),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_736),
.Y(n_833)
);

NAND2xp33_ASAP7_75t_L g834 ( 
.A(n_711),
.B(n_318),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_723),
.B(n_318),
.Y(n_835)
);

OAI221xp5_ASAP7_75t_L g836 ( 
.A1(n_664),
.A2(n_643),
.B1(n_639),
.B2(n_638),
.C(n_632),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_763),
.B(n_731),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_653),
.B(n_630),
.Y(n_838)
);

AND2x6_ASAP7_75t_SL g839 ( 
.A(n_665),
.B(n_233),
.Y(n_839)
);

NAND2xp33_ASAP7_75t_L g840 ( 
.A(n_711),
.B(n_318),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_654),
.B(n_510),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_748),
.A2(n_448),
.B1(n_449),
.B2(n_440),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_737),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_763),
.B(n_318),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_763),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_658),
.B(n_630),
.Y(n_846)
);

BUFx6f_ASAP7_75t_SL g847 ( 
.A(n_645),
.Y(n_847)
);

INVx5_ASAP7_75t_L g848 ( 
.A(n_796),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_748),
.B(n_627),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_696),
.Y(n_850)
);

INVx1_ASAP7_75t_SL g851 ( 
.A(n_684),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_737),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_763),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_738),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_750),
.A2(n_656),
.B1(n_747),
.B2(n_786),
.Y(n_855)
);

NAND3xp33_ASAP7_75t_L g856 ( 
.A(n_708),
.B(n_516),
.C(n_510),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_798),
.B(n_790),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_667),
.B(n_516),
.Y(n_858)
);

INVxp67_ASAP7_75t_SL g859 ( 
.A(n_652),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_658),
.B(n_630),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_790),
.A2(n_324),
.B1(n_327),
.B2(n_288),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_750),
.B(n_318),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_696),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_663),
.B(n_640),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_724),
.B(n_521),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_738),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_663),
.B(n_640),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_684),
.B(n_521),
.Y(n_868)
);

NAND2xp33_ASAP7_75t_L g869 ( 
.A(n_711),
.B(n_318),
.Y(n_869)
);

BUFx10_ASAP7_75t_L g870 ( 
.A(n_686),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_753),
.B(n_318),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_689),
.B(n_690),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_758),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_740),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_689),
.B(n_690),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_652),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_778),
.B(n_528),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_753),
.B(n_640),
.Y(n_878)
);

NAND3xp33_ASAP7_75t_L g879 ( 
.A(n_727),
.B(n_531),
.C(n_528),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_755),
.B(n_640),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_700),
.B(n_673),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_755),
.B(n_640),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_695),
.B(n_640),
.Y(n_883)
);

OA21x2_ASAP7_75t_L g884 ( 
.A1(n_759),
.A2(n_564),
.B(n_604),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_759),
.B(n_640),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_695),
.B(n_699),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_699),
.B(n_642),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_710),
.B(n_531),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_744),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_697),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_744),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_767),
.B(n_642),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_701),
.B(n_642),
.Y(n_893)
);

INVx4_ASAP7_75t_L g894 ( 
.A(n_785),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_694),
.B(n_532),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_749),
.Y(n_896)
);

NAND3xp33_ASAP7_75t_L g897 ( 
.A(n_792),
.B(n_547),
.C(n_532),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_792),
.Y(n_898)
);

OAI22xp33_ASAP7_75t_L g899 ( 
.A1(n_729),
.A2(n_548),
.B1(n_547),
.B2(n_327),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_709),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_749),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_697),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_659),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_701),
.B(n_642),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_657),
.B(n_631),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_702),
.B(n_642),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_702),
.B(n_642),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_751),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_800),
.B(n_548),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_751),
.Y(n_910)
);

INVx8_ASAP7_75t_L g911 ( 
.A(n_647),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_767),
.B(n_642),
.Y(n_912)
);

A2O1A1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_666),
.A2(n_564),
.B(n_274),
.C(n_277),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_703),
.B(n_625),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_647),
.A2(n_333),
.B1(n_337),
.B2(n_266),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_704),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_703),
.B(n_625),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_779),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_779),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_704),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_739),
.B(n_631),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_647),
.A2(n_353),
.B1(n_261),
.B2(n_269),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_657),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_791),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_709),
.Y(n_925)
);

NOR2xp67_ASAP7_75t_L g926 ( 
.A(n_693),
.B(n_632),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_718),
.A2(n_263),
.B1(n_271),
.B2(n_270),
.Y(n_927)
);

NOR3xp33_ASAP7_75t_L g928 ( 
.A(n_707),
.B(n_639),
.C(n_638),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_794),
.B(n_643),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_791),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_705),
.B(n_625),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_706),
.Y(n_932)
);

NAND2xp33_ASAP7_75t_L g933 ( 
.A(n_711),
.B(n_324),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_794),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_706),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_797),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_716),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_777),
.A2(n_380),
.B(n_274),
.C(n_277),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_L g939 ( 
.A1(n_705),
.A2(n_406),
.B1(n_393),
.B2(n_397),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_774),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_793),
.B(n_334),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_797),
.Y(n_942)
);

AO221x1_ASAP7_75t_L g943 ( 
.A1(n_677),
.A2(n_339),
.B1(n_429),
.B2(n_244),
.C(n_424),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_725),
.B(n_641),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_769),
.B(n_641),
.Y(n_945)
);

AO22x1_ASAP7_75t_L g946 ( 
.A1(n_756),
.A2(n_280),
.B1(n_294),
.B2(n_278),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_657),
.B(n_604),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_698),
.Y(n_948)
);

INVxp67_ASAP7_75t_L g949 ( 
.A(n_671),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_698),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_775),
.B(n_338),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_698),
.B(n_605),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_769),
.B(n_341),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_758),
.Y(n_954)
);

INVxp67_ASAP7_75t_L g955 ( 
.A(n_775),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_716),
.B(n_717),
.Y(n_956)
);

OR2x2_ASAP7_75t_L g957 ( 
.A(n_733),
.B(n_343),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_717),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_742),
.B(n_344),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_645),
.B(n_357),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_718),
.A2(n_331),
.B1(n_431),
.B2(n_273),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_719),
.B(n_605),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_719),
.B(n_560),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_734),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_648),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_734),
.B(n_272),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_768),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_645),
.B(n_403),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_735),
.B(n_560),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_735),
.B(n_567),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_718),
.B(n_352),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_741),
.B(n_275),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_865),
.B(n_645),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_929),
.B(n_733),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_913),
.A2(n_745),
.B(n_746),
.C(n_741),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_812),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_814),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_857),
.A2(n_760),
.B(n_772),
.Y(n_978)
);

HB1xp67_ASAP7_75t_L g979 ( 
.A(n_851),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_965),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_806),
.B(n_677),
.Y(n_981)
);

NAND2x1p5_ASAP7_75t_L g982 ( 
.A(n_853),
.B(n_655),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_898),
.B(n_682),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_857),
.A2(n_680),
.B(n_662),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_809),
.A2(n_680),
.B(n_662),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_881),
.A2(n_646),
.B1(n_677),
.B2(n_760),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_952),
.A2(n_680),
.B(n_662),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_868),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_806),
.B(n_677),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_855),
.A2(n_760),
.B1(n_772),
.B2(n_646),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_898),
.B(n_682),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_806),
.A2(n_646),
.B1(n_760),
.B2(n_732),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_802),
.A2(n_670),
.B(n_655),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_926),
.B(n_712),
.Y(n_994)
);

AOI22xp5_ASAP7_75t_L g995 ( 
.A1(n_877),
.A2(n_646),
.B1(n_760),
.B2(n_732),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_805),
.A2(n_670),
.B(n_655),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_934),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_947),
.A2(n_670),
.B(n_655),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_821),
.B(n_745),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_816),
.B(n_714),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_825),
.B(n_746),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_947),
.A2(n_675),
.B(n_670),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_R g1003 ( 
.A1(n_903),
.A2(n_355),
.B1(n_356),
.B2(n_354),
.Y(n_1003)
);

INVx1_ASAP7_75t_SL g1004 ( 
.A(n_940),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_918),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_816),
.B(n_752),
.Y(n_1006)
);

OA22x2_ASAP7_75t_L g1007 ( 
.A1(n_943),
.A2(n_810),
.B1(n_824),
.B2(n_900),
.Y(n_1007)
);

AOI33xp33_ASAP7_75t_L g1008 ( 
.A1(n_900),
.A2(n_776),
.A3(n_295),
.B1(n_371),
.B2(n_317),
.B3(n_424),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_814),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_913),
.A2(n_757),
.B(n_752),
.C(n_772),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_951),
.A2(n_832),
.B(n_921),
.C(n_941),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_859),
.A2(n_787),
.B(n_675),
.Y(n_1012)
);

INVx4_ASAP7_75t_L g1013 ( 
.A(n_812),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_919),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_849),
.B(n_757),
.Y(n_1015)
);

OA21x2_ASAP7_75t_L g1016 ( 
.A1(n_803),
.A2(n_789),
.B(n_771),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_827),
.B(n_828),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_830),
.B(n_768),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_963),
.A2(n_787),
.B(n_675),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_812),
.Y(n_1020)
);

INVx2_ASAP7_75t_SL g1021 ( 
.A(n_945),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_862),
.A2(n_962),
.B(n_956),
.Y(n_1022)
);

BUFx4f_ASAP7_75t_L g1023 ( 
.A(n_911),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_833),
.B(n_771),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_843),
.B(n_773),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_852),
.B(n_773),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_849),
.B(n_780),
.Y(n_1027)
);

AOI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_801),
.A2(n_711),
.B1(n_732),
.B2(n_780),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_969),
.A2(n_787),
.B(n_675),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_938),
.A2(n_772),
.B(n_574),
.C(n_571),
.Y(n_1030)
);

OR2x6_ASAP7_75t_L g1031 ( 
.A(n_911),
.B(n_681),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_813),
.A2(n_788),
.B(n_787),
.Y(n_1032)
);

INVx4_ASAP7_75t_L g1033 ( 
.A(n_812),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_862),
.A2(n_772),
.B(n_732),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_813),
.A2(n_788),
.B(n_649),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_854),
.B(n_784),
.Y(n_1036)
);

CKINVDCx10_ASAP7_75t_R g1037 ( 
.A(n_847),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_819),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_866),
.B(n_784),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_925),
.B(n_681),
.Y(n_1040)
);

INVxp67_ASAP7_75t_L g1041 ( 
.A(n_822),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_874),
.B(n_711),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_955),
.A2(n_783),
.B1(n_374),
.B2(n_393),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_894),
.A2(n_788),
.B(n_649),
.Y(n_1044)
);

NAND2x1p5_ASAP7_75t_L g1045 ( 
.A(n_853),
.B(n_788),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_894),
.A2(n_965),
.B(n_835),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_894),
.A2(n_649),
.B(n_648),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_849),
.B(n_283),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_962),
.A2(n_732),
.B(n_661),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_965),
.A2(n_649),
.B(n_648),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_965),
.A2(n_649),
.B(n_648),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_826),
.A2(n_722),
.B(n_715),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_835),
.A2(n_722),
.B(n_715),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_844),
.A2(n_722),
.B(n_715),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_SL g1055 ( 
.A1(n_844),
.A2(n_406),
.B(n_369),
.C(n_421),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_845),
.A2(n_722),
.B(n_715),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_889),
.B(n_732),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_888),
.B(n_795),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_949),
.B(n_411),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_804),
.B(n_414),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_842),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_845),
.A2(n_715),
.B(n_650),
.Y(n_1062)
);

OAI21xp33_ASAP7_75t_L g1063 ( 
.A1(n_909),
.A2(n_363),
.B(n_362),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_876),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_891),
.B(n_660),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_872),
.A2(n_715),
.B(n_650),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_808),
.A2(n_374),
.B1(n_397),
.B2(n_421),
.Y(n_1067)
);

OAI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_924),
.A2(n_661),
.B(n_660),
.Y(n_1068)
);

OAI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_930),
.A2(n_674),
.B(n_669),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_875),
.A2(n_743),
.B(n_650),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_886),
.A2(n_837),
.B(n_815),
.Y(n_1071)
);

NOR2x2_ASAP7_75t_L g1072 ( 
.A(n_839),
.B(n_811),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_936),
.A2(n_674),
.B(n_669),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_923),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_923),
.B(n_285),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_942),
.Y(n_1076)
);

BUFx2_ASAP7_75t_L g1077 ( 
.A(n_820),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_896),
.B(n_678),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_837),
.A2(n_743),
.B(n_650),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_838),
.A2(n_860),
.B(n_846),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_841),
.B(n_672),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_829),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_864),
.A2(n_743),
.B(n_650),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_876),
.A2(n_950),
.B1(n_861),
.B2(n_807),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_858),
.B(n_672),
.Y(n_1085)
);

INVxp67_ASAP7_75t_L g1086 ( 
.A(n_905),
.Y(n_1086)
);

AOI21x1_ASAP7_75t_L g1087 ( 
.A1(n_878),
.A2(n_651),
.B(n_789),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_923),
.B(n_290),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_901),
.B(n_678),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_953),
.B(n_795),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_923),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_950),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_908),
.B(n_679),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_867),
.A2(n_743),
.B(n_650),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_911),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_895),
.B(n_672),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_905),
.B(n_369),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_911),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_910),
.B(n_905),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_883),
.A2(n_799),
.B(n_743),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_829),
.Y(n_1101)
);

NOR3xp33_ASAP7_75t_L g1102 ( 
.A(n_897),
.B(n_428),
.C(n_367),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_887),
.A2(n_799),
.B(n_743),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_948),
.B(n_679),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_893),
.A2(n_687),
.B(n_683),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_831),
.B(n_683),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_959),
.A2(n_428),
.B(n_687),
.C(n_688),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_848),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_831),
.B(n_688),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_904),
.A2(n_799),
.B(n_762),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_906),
.A2(n_907),
.B(n_863),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_970),
.A2(n_848),
.B(n_914),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_848),
.A2(n_799),
.B(n_762),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_850),
.B(n_754),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_957),
.B(n_676),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_850),
.A2(n_890),
.B(n_863),
.Y(n_1116)
);

NOR2x1p5_ASAP7_75t_L g1117 ( 
.A(n_903),
.B(n_364),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_890),
.B(n_902),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_902),
.B(n_754),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_916),
.B(n_754),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_916),
.B(n_754),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_856),
.B(n_676),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_848),
.A2(n_931),
.B(n_917),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_920),
.A2(n_651),
.B(n_676),
.Y(n_1124)
);

NAND3xp33_ASAP7_75t_L g1125 ( 
.A(n_928),
.B(n_373),
.C(n_368),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_899),
.B(n_301),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_920),
.B(n_932),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_932),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_848),
.A2(n_799),
.B(n_764),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_935),
.B(n_761),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_935),
.A2(n_958),
.B(n_937),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_937),
.B(n_761),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_958),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_873),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_964),
.A2(n_764),
.B(n_762),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_873),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_964),
.B(n_761),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_954),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_967),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_944),
.A2(n_766),
.B(n_764),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_817),
.B(n_278),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_873),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_870),
.B(n_376),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_878),
.A2(n_770),
.B(n_766),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_871),
.Y(n_1145)
);

NOR2xp67_ASAP7_75t_L g1146 ( 
.A(n_879),
.B(n_302),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_880),
.A2(n_770),
.B(n_761),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_880),
.A2(n_770),
.B(n_573),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_882),
.A2(n_573),
.B(n_570),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_966),
.B(n_795),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_870),
.B(n_377),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_971),
.A2(n_415),
.B(n_385),
.C(n_289),
.Y(n_1152)
);

O2A1O1Ixp33_ASAP7_75t_SL g1153 ( 
.A1(n_871),
.A2(n_571),
.B(n_574),
.C(n_395),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_882),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_885),
.A2(n_796),
.B(n_572),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_966),
.B(n_795),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_870),
.B(n_378),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_885),
.A2(n_573),
.B(n_570),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_972),
.B(n_785),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_892),
.Y(n_1160)
);

NAND2x1p5_ASAP7_75t_L g1161 ( 
.A(n_892),
.B(n_912),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_972),
.B(n_939),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1011),
.B(n_884),
.Y(n_1163)
);

O2A1O1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_994),
.A2(n_817),
.B(n_836),
.C(n_938),
.Y(n_1164)
);

NAND3xp33_ASAP7_75t_L g1165 ( 
.A(n_1060),
.B(n_915),
.C(n_960),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_979),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_984),
.A2(n_933),
.B(n_834),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_973),
.B(n_988),
.Y(n_1168)
);

INVxp67_ASAP7_75t_SL g1169 ( 
.A(n_1074),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_SL g1170 ( 
.A1(n_1150),
.A2(n_912),
.B(n_922),
.C(n_961),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1021),
.B(n_884),
.Y(n_1171)
);

INVx4_ASAP7_75t_L g1172 ( 
.A(n_1095),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_995),
.A2(n_847),
.B1(n_968),
.B2(n_927),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1041),
.B(n_884),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_1095),
.B(n_823),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1082),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_979),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1101),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_985),
.A2(n_933),
.B(n_834),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_1060),
.B(n_847),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1041),
.B(n_946),
.Y(n_1181)
);

BUFx8_ASAP7_75t_SL g1182 ( 
.A(n_1061),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1133),
.Y(n_1183)
);

A2O1A1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1010),
.A2(n_869),
.B(n_840),
.C(n_818),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_R g1185 ( 
.A(n_1023),
.B(n_818),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1019),
.A2(n_869),
.B(n_840),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1017),
.B(n_785),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1086),
.B(n_785),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_1004),
.Y(n_1189)
);

NOR2x1_ASAP7_75t_SL g1190 ( 
.A(n_980),
.B(n_280),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_1074),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_1095),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1102),
.A2(n_282),
.B1(n_427),
.B2(n_426),
.Y(n_1193)
);

INVx1_ASAP7_75t_SL g1194 ( 
.A(n_997),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1029),
.A2(n_573),
.B(n_570),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_983),
.A2(n_360),
.B1(n_304),
.B2(n_316),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_991),
.A2(n_413),
.B1(n_323),
.B2(n_329),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_992),
.A2(n_317),
.B1(n_380),
.B2(n_379),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1005),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1014),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1010),
.A2(n_429),
.B(n_423),
.C(n_339),
.Y(n_1201)
);

NAND2x1p5_ASAP7_75t_L g1202 ( 
.A(n_1095),
.B(n_573),
.Y(n_1202)
);

O2A1O1Ixp5_ASAP7_75t_L g1203 ( 
.A1(n_1081),
.A2(n_289),
.B(n_385),
.C(n_295),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_1077),
.Y(n_1204)
);

INVx5_ASAP7_75t_L g1205 ( 
.A(n_1108),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1115),
.A2(n_395),
.B(n_394),
.C(n_294),
.Y(n_1206)
);

BUFx12f_ASAP7_75t_L g1207 ( 
.A(n_1031),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_974),
.B(n_383),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_977),
.Y(n_1209)
);

O2A1O1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_1000),
.A2(n_423),
.B(n_379),
.C(n_371),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1074),
.Y(n_1211)
);

AND2x4_ASAP7_75t_L g1212 ( 
.A(n_1098),
.B(n_346),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_R g1213 ( 
.A(n_1023),
.B(n_330),
.Y(n_1213)
);

NAND3xp33_ASAP7_75t_SL g1214 ( 
.A(n_1102),
.B(n_398),
.C(n_433),
.Y(n_1214)
);

INVx1_ASAP7_75t_SL g1215 ( 
.A(n_1040),
.Y(n_1215)
);

A2O1A1Ixp33_ASAP7_75t_SL g1216 ( 
.A1(n_1115),
.A2(n_572),
.B(n_586),
.C(n_581),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1076),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1086),
.A2(n_335),
.B1(n_342),
.B2(n_345),
.Y(n_1218)
);

OAI21xp33_ASAP7_75t_L g1219 ( 
.A1(n_1063),
.A2(n_399),
.B(n_432),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1090),
.A2(n_382),
.B1(n_347),
.B2(n_350),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1064),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1009),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1162),
.A2(n_394),
.B(n_346),
.C(n_358),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1044),
.A2(n_573),
.B(n_585),
.Y(n_1224)
);

CKINVDCx20_ASAP7_75t_R g1225 ( 
.A(n_1098),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1038),
.Y(n_1226)
);

AOI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1059),
.A2(n_389),
.B1(n_359),
.B2(n_366),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1081),
.B(n_796),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1059),
.B(n_386),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1058),
.B(n_387),
.Y(n_1230)
);

AO32x2_ASAP7_75t_L g1231 ( 
.A1(n_990),
.A2(n_358),
.A3(n_14),
.B1(n_15),
.B2(n_18),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_978),
.A2(n_573),
.B(n_585),
.Y(n_1232)
);

NAND2x2_ASAP7_75t_L g1233 ( 
.A(n_1117),
.B(n_391),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1098),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1087),
.A2(n_586),
.B(n_581),
.Y(n_1235)
);

AOI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1071),
.A2(n_579),
.B(n_586),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_1141),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_SL g1238 ( 
.A(n_1099),
.B(n_1064),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1030),
.A2(n_372),
.B(n_381),
.C(n_388),
.Y(n_1239)
);

A2O1A1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1030),
.A2(n_419),
.B(n_401),
.C(n_425),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1128),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1046),
.A2(n_585),
.B(n_576),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1096),
.A2(n_418),
.B(n_407),
.C(n_404),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_R g1244 ( 
.A(n_1098),
.B(n_400),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1085),
.B(n_796),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1141),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1085),
.B(n_796),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1034),
.A2(n_585),
.B(n_581),
.Y(n_1248)
);

O2A1O1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1126),
.A2(n_579),
.B(n_576),
.C(n_572),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1096),
.B(n_402),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1065),
.Y(n_1251)
);

BUFx12f_ASAP7_75t_L g1252 ( 
.A(n_1031),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1092),
.B(n_408),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_986),
.A2(n_410),
.B(n_412),
.C(n_416),
.Y(n_1254)
);

O2A1O1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1152),
.A2(n_567),
.B(n_576),
.C(n_579),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1012),
.A2(n_585),
.B(n_796),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_981),
.A2(n_436),
.B1(n_420),
.B2(n_585),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_987),
.A2(n_585),
.B(n_796),
.Y(n_1258)
);

INVx4_ASAP7_75t_L g1259 ( 
.A(n_1074),
.Y(n_1259)
);

INVxp33_ASAP7_75t_L g1260 ( 
.A(n_1143),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1151),
.B(n_13),
.Y(n_1261)
);

HB1xp67_ASAP7_75t_L g1262 ( 
.A(n_1097),
.Y(n_1262)
);

A2O1A1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1122),
.A2(n_1022),
.B(n_1125),
.C(n_1156),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_SL g1264 ( 
.A(n_1092),
.B(n_1157),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1097),
.B(n_19),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1145),
.B(n_221),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1154),
.B(n_220),
.Y(n_1267)
);

INVx8_ASAP7_75t_L g1268 ( 
.A(n_980),
.Y(n_1268)
);

INVx2_ASAP7_75t_SL g1269 ( 
.A(n_1037),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_989),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1032),
.A2(n_219),
.B(n_217),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_1031),
.B(n_1013),
.Y(n_1272)
);

AND2x2_ASAP7_75t_SL g1273 ( 
.A(n_1008),
.B(n_20),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1134),
.Y(n_1274)
);

CKINVDCx14_ASAP7_75t_R g1275 ( 
.A(n_1003),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1146),
.B(n_1013),
.Y(n_1276)
);

INVxp67_ASAP7_75t_L g1277 ( 
.A(n_1048),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_998),
.A2(n_215),
.B(n_214),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_980),
.Y(n_1279)
);

AOI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1084),
.A2(n_209),
.B1(n_207),
.B2(n_206),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1002),
.A2(n_184),
.B(n_178),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1078),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1134),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_SL g1284 ( 
.A(n_1033),
.B(n_175),
.Y(n_1284)
);

INVx4_ASAP7_75t_L g1285 ( 
.A(n_980),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1138),
.Y(n_1286)
);

O2A1O1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1067),
.A2(n_21),
.B(n_26),
.C(n_27),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1160),
.B(n_170),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_999),
.B(n_167),
.Y(n_1289)
);

CKINVDCx16_ASAP7_75t_R g1290 ( 
.A(n_1043),
.Y(n_1290)
);

O2A1O1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_1015),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_1291)
);

AOI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1080),
.A2(n_152),
.B(n_146),
.Y(n_1292)
);

INVx5_ASAP7_75t_L g1293 ( 
.A(n_1108),
.Y(n_1293)
);

AOI221xp5_ASAP7_75t_L g1294 ( 
.A1(n_1139),
.A2(n_28),
.B1(n_29),
.B2(n_32),
.C(n_33),
.Y(n_1294)
);

O2A1O1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1107),
.A2(n_29),
.B(n_32),
.C(n_34),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_976),
.Y(n_1296)
);

O2A1O1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1006),
.A2(n_1027),
.B(n_1001),
.C(n_1055),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1033),
.B(n_145),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1018),
.B(n_140),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_SL g1300 ( 
.A(n_1136),
.B(n_134),
.Y(n_1300)
);

A2O1A1Ixp33_ASAP7_75t_SL g1301 ( 
.A1(n_1122),
.A2(n_975),
.B(n_1135),
.C(n_1091),
.Y(n_1301)
);

A2O1A1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_975),
.A2(n_34),
.B(n_35),
.C(n_37),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1024),
.B(n_43),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1118),
.Y(n_1304)
);

A2O1A1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1028),
.A2(n_53),
.B(n_56),
.C(n_58),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1136),
.B(n_130),
.Y(n_1306)
);

BUFx6f_ASAP7_75t_L g1307 ( 
.A(n_1136),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_SL g1308 ( 
.A(n_1136),
.B(n_126),
.Y(n_1308)
);

INVx2_ASAP7_75t_SL g1309 ( 
.A(n_976),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1007),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_1310)
);

AND2x4_ASAP7_75t_L g1311 ( 
.A(n_1020),
.B(n_107),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_SL g1312 ( 
.A(n_1142),
.B(n_120),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_1007),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_1020),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1089),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1025),
.B(n_116),
.Y(n_1316)
);

INVx6_ASAP7_75t_L g1317 ( 
.A(n_1142),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_993),
.A2(n_996),
.B(n_1047),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1127),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1142),
.B(n_115),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1026),
.B(n_59),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1036),
.A2(n_61),
.B1(n_63),
.B2(n_65),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1142),
.Y(n_1323)
);

A2O1A1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1042),
.A2(n_61),
.B(n_63),
.C(n_65),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_1075),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1039),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1123),
.A2(n_109),
.B(n_106),
.Y(n_1327)
);

NAND2x1p5_ASAP7_75t_L g1328 ( 
.A(n_1108),
.B(n_97),
.Y(n_1328)
);

AO22x2_ASAP7_75t_L g1329 ( 
.A1(n_1310),
.A2(n_1072),
.B1(n_1159),
.B2(n_1057),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1199),
.Y(n_1330)
);

INVx2_ASAP7_75t_SL g1331 ( 
.A(n_1166),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1290),
.A2(n_1045),
.B1(n_982),
.B2(n_1093),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_1182),
.Y(n_1333)
);

AOI221x1_ASAP7_75t_L g1334 ( 
.A1(n_1261),
.A2(n_1111),
.B1(n_1112),
.B2(n_1124),
.C(n_1140),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1260),
.B(n_1088),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1235),
.A2(n_1116),
.B(n_1131),
.Y(n_1336)
);

OR2x6_ASAP7_75t_L g1337 ( 
.A(n_1268),
.B(n_982),
.Y(n_1337)
);

OAI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1263),
.A2(n_1049),
.B(n_1105),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1186),
.A2(n_1108),
.B(n_1035),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1286),
.Y(n_1340)
);

A2O1A1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1229),
.A2(n_1147),
.B(n_1144),
.C(n_1110),
.Y(n_1341)
);

A2O1A1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1164),
.A2(n_1104),
.B(n_1070),
.C(n_1066),
.Y(n_1342)
);

BUFx10_ASAP7_75t_L g1343 ( 
.A(n_1175),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_1189),
.Y(n_1344)
);

AOI221x1_ASAP7_75t_L g1345 ( 
.A1(n_1302),
.A2(n_1069),
.B1(n_1073),
.B2(n_1068),
.C(n_1062),
.Y(n_1345)
);

O2A1O1Ixp5_ASAP7_75t_L g1346 ( 
.A1(n_1203),
.A2(n_1079),
.B(n_1056),
.C(n_1052),
.Y(n_1346)
);

AO21x1_ASAP7_75t_L g1347 ( 
.A1(n_1310),
.A2(n_1161),
.B(n_1045),
.Y(n_1347)
);

AOI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1208),
.A2(n_1161),
.B1(n_1153),
.B2(n_1016),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1326),
.B(n_1109),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1236),
.A2(n_1148),
.B(n_1050),
.Y(n_1350)
);

O2A1O1Ixp5_ASAP7_75t_SL g1351 ( 
.A1(n_1270),
.A2(n_1155),
.B(n_1106),
.C(n_1121),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1163),
.A2(n_1120),
.B(n_1137),
.Y(n_1352)
);

AOI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1165),
.A2(n_1016),
.B1(n_1119),
.B2(n_1132),
.Y(n_1353)
);

AO31x2_ASAP7_75t_L g1354 ( 
.A1(n_1201),
.A2(n_1053),
.A3(n_1054),
.B(n_1051),
.Y(n_1354)
);

AO31x2_ASAP7_75t_L g1355 ( 
.A1(n_1239),
.A2(n_1240),
.A3(n_1318),
.B(n_1206),
.Y(n_1355)
);

AOI21xp33_ASAP7_75t_L g1356 ( 
.A1(n_1250),
.A2(n_1114),
.B(n_1130),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1184),
.A2(n_1158),
.B(n_1149),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1204),
.B(n_1103),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1195),
.A2(n_1100),
.B(n_1094),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1248),
.A2(n_1083),
.B(n_1113),
.Y(n_1360)
);

OAI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1167),
.A2(n_1129),
.B(n_95),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1258),
.A2(n_92),
.B(n_70),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1179),
.A2(n_67),
.B(n_70),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1251),
.B(n_1282),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1177),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1301),
.A2(n_72),
.B(n_73),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1313),
.A2(n_76),
.B1(n_78),
.B2(n_80),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1272),
.B(n_76),
.Y(n_1368)
);

AOI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1181),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_1369)
);

BUFx6f_ASAP7_75t_L g1370 ( 
.A(n_1192),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1242),
.A2(n_81),
.B(n_84),
.Y(n_1371)
);

O2A1O1Ixp33_ASAP7_75t_L g1372 ( 
.A1(n_1168),
.A2(n_87),
.B(n_88),
.C(n_1181),
.Y(n_1372)
);

A2O1A1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1303),
.A2(n_1254),
.B(n_1180),
.C(n_1297),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_1269),
.Y(n_1374)
);

AO31x2_ASAP7_75t_L g1375 ( 
.A1(n_1223),
.A2(n_87),
.A3(n_1198),
.B(n_1232),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1315),
.A2(n_1198),
.B1(n_1200),
.B2(n_1217),
.Y(n_1376)
);

INVx2_ASAP7_75t_SL g1377 ( 
.A(n_1194),
.Y(n_1377)
);

BUFx3_ASAP7_75t_L g1378 ( 
.A(n_1225),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1246),
.B(n_1230),
.Y(n_1379)
);

BUFx10_ASAP7_75t_L g1380 ( 
.A(n_1175),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1237),
.B(n_1262),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1209),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1304),
.B(n_1319),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1321),
.B(n_1277),
.Y(n_1384)
);

NAND3xp33_ASAP7_75t_SL g1385 ( 
.A(n_1193),
.B(n_1227),
.C(n_1325),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1176),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1228),
.A2(n_1247),
.B(n_1245),
.Y(n_1387)
);

AO31x2_ASAP7_75t_L g1388 ( 
.A1(n_1305),
.A2(n_1257),
.A3(n_1245),
.B(n_1228),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1289),
.A2(n_1299),
.B(n_1316),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1238),
.B(n_1264),
.Y(n_1390)
);

A2O1A1Ixp33_ASAP7_75t_L g1391 ( 
.A1(n_1280),
.A2(n_1214),
.B(n_1219),
.C(n_1299),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1224),
.A2(n_1256),
.B(n_1292),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1266),
.A2(n_1288),
.B(n_1267),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1265),
.B(n_1221),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1222),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1289),
.A2(n_1316),
.B(n_1247),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1187),
.A2(n_1266),
.B(n_1170),
.Y(n_1397)
);

INVx2_ASAP7_75t_SL g1398 ( 
.A(n_1215),
.Y(n_1398)
);

AOI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1173),
.A2(n_1273),
.B1(n_1294),
.B2(n_1270),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1173),
.B(n_1196),
.Y(n_1400)
);

O2A1O1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_1287),
.A2(n_1322),
.B(n_1324),
.C(n_1295),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1178),
.Y(n_1402)
);

INVx3_ASAP7_75t_SL g1403 ( 
.A(n_1212),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1183),
.Y(n_1404)
);

AND2x4_ASAP7_75t_L g1405 ( 
.A(n_1272),
.B(n_1296),
.Y(n_1405)
);

A2O1A1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1243),
.A2(n_1267),
.B(n_1288),
.C(n_1291),
.Y(n_1406)
);

AOI221x1_ASAP7_75t_L g1407 ( 
.A1(n_1322),
.A2(n_1257),
.B1(n_1281),
.B2(n_1278),
.C(n_1271),
.Y(n_1407)
);

INVxp67_ASAP7_75t_L g1408 ( 
.A(n_1212),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1187),
.A2(n_1174),
.B(n_1293),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1249),
.A2(n_1255),
.B(n_1171),
.Y(n_1410)
);

A2O1A1Ixp33_ASAP7_75t_L g1411 ( 
.A1(n_1210),
.A2(n_1253),
.B(n_1327),
.C(n_1220),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_SL g1412 ( 
.A1(n_1190),
.A2(n_1174),
.B(n_1171),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1188),
.A2(n_1202),
.B(n_1276),
.Y(n_1413)
);

NAND2xp33_ASAP7_75t_L g1414 ( 
.A(n_1185),
.B(n_1234),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1197),
.B(n_1244),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1205),
.A2(n_1293),
.B(n_1216),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1188),
.A2(n_1241),
.B(n_1226),
.Y(n_1417)
);

AOI221xp5_ASAP7_75t_L g1418 ( 
.A1(n_1275),
.A2(n_1284),
.B1(n_1298),
.B2(n_1308),
.C(n_1306),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1311),
.A2(n_1283),
.B1(n_1274),
.B2(n_1320),
.Y(n_1419)
);

BUFx6f_ASAP7_75t_L g1420 ( 
.A(n_1192),
.Y(n_1420)
);

BUFx2_ASAP7_75t_L g1421 ( 
.A(n_1314),
.Y(n_1421)
);

XNOR2xp5_ASAP7_75t_L g1422 ( 
.A(n_1218),
.B(n_1311),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1320),
.B(n_1169),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1309),
.B(n_1323),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1202),
.A2(n_1211),
.B(n_1191),
.Y(n_1425)
);

AO31x2_ASAP7_75t_L g1426 ( 
.A1(n_1231),
.A2(n_1259),
.A3(n_1285),
.B(n_1172),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1205),
.A2(n_1293),
.B(n_1312),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1191),
.B(n_1211),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1279),
.Y(n_1429)
);

INVx1_ASAP7_75t_SL g1430 ( 
.A(n_1317),
.Y(n_1430)
);

INVx1_ASAP7_75t_SL g1431 ( 
.A(n_1317),
.Y(n_1431)
);

OAI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1300),
.A2(n_1328),
.B(n_1259),
.Y(n_1432)
);

AOI221x1_ASAP7_75t_L g1433 ( 
.A1(n_1231),
.A2(n_1285),
.B1(n_1307),
.B2(n_1279),
.C(n_1172),
.Y(n_1433)
);

OA21x2_ASAP7_75t_L g1434 ( 
.A1(n_1231),
.A2(n_1328),
.B(n_1317),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1205),
.A2(n_1293),
.B(n_1268),
.Y(n_1435)
);

INVx6_ASAP7_75t_SL g1436 ( 
.A(n_1233),
.Y(n_1436)
);

AOI221x1_ASAP7_75t_L g1437 ( 
.A1(n_1307),
.A2(n_1279),
.B1(n_1234),
.B2(n_1207),
.C(n_1252),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1205),
.A2(n_1268),
.B(n_1307),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1213),
.B(n_973),
.Y(n_1439)
);

AO221x2_ASAP7_75t_L g1440 ( 
.A1(n_1270),
.A2(n_1322),
.B1(n_1310),
.B2(n_899),
.C(n_1165),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1186),
.A2(n_1011),
.B(n_1318),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1192),
.Y(n_1442)
);

OA21x2_ASAP7_75t_L g1443 ( 
.A1(n_1163),
.A2(n_1263),
.B(n_1203),
.Y(n_1443)
);

INVx2_ASAP7_75t_SL g1444 ( 
.A(n_1166),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1204),
.B(n_988),
.Y(n_1445)
);

A2O1A1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1261),
.A2(n_1011),
.B(n_881),
.C(n_1060),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1186),
.A2(n_1011),
.B(n_1318),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1186),
.A2(n_1011),
.B(n_1318),
.Y(n_1448)
);

NAND2x1_ASAP7_75t_L g1449 ( 
.A(n_1172),
.B(n_1013),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1326),
.B(n_973),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1186),
.A2(n_1011),
.B(n_1318),
.Y(n_1451)
);

INVxp67_ASAP7_75t_L g1452 ( 
.A(n_1166),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1186),
.A2(n_1011),
.B(n_1318),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1186),
.A2(n_1011),
.B(n_1318),
.Y(n_1454)
);

O2A1O1Ixp33_ASAP7_75t_SL g1455 ( 
.A1(n_1305),
.A2(n_1011),
.B(n_1184),
.C(n_1263),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1272),
.B(n_1175),
.Y(n_1456)
);

A2O1A1Ixp33_ASAP7_75t_L g1457 ( 
.A1(n_1261),
.A2(n_1011),
.B(n_881),
.C(n_1060),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1235),
.A2(n_1236),
.B(n_1318),
.Y(n_1458)
);

AO31x2_ASAP7_75t_L g1459 ( 
.A1(n_1163),
.A2(n_1201),
.A3(n_990),
.B(n_1263),
.Y(n_1459)
);

AO31x2_ASAP7_75t_L g1460 ( 
.A1(n_1163),
.A2(n_1201),
.A3(n_990),
.B(n_1263),
.Y(n_1460)
);

OAI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1263),
.A2(n_1011),
.B(n_1163),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1326),
.B(n_973),
.Y(n_1462)
);

OAI22x1_ASAP7_75t_L g1463 ( 
.A1(n_1261),
.A2(n_1060),
.B1(n_1165),
.B2(n_881),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1186),
.A2(n_1011),
.B(n_1318),
.Y(n_1464)
);

INVx3_ASAP7_75t_L g1465 ( 
.A(n_1307),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_L g1466 ( 
.A(n_1192),
.Y(n_1466)
);

NAND2x2_ASAP7_75t_L g1467 ( 
.A(n_1269),
.B(n_681),
.Y(n_1467)
);

AO31x2_ASAP7_75t_L g1468 ( 
.A1(n_1163),
.A2(n_1201),
.A3(n_990),
.B(n_1263),
.Y(n_1468)
);

AO21x1_ASAP7_75t_L g1469 ( 
.A1(n_1261),
.A2(n_990),
.B(n_1310),
.Y(n_1469)
);

O2A1O1Ixp33_ASAP7_75t_SL g1470 ( 
.A1(n_1305),
.A2(n_1011),
.B(n_1184),
.C(n_1263),
.Y(n_1470)
);

NAND3xp33_ASAP7_75t_SL g1471 ( 
.A(n_1261),
.B(n_1011),
.C(n_1060),
.Y(n_1471)
);

AO31x2_ASAP7_75t_L g1472 ( 
.A1(n_1163),
.A2(n_1201),
.A3(n_990),
.B(n_1263),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1261),
.A2(n_1060),
.B1(n_881),
.B2(n_1229),
.Y(n_1473)
);

OAI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1263),
.A2(n_1011),
.B(n_1163),
.Y(n_1474)
);

AOI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1186),
.A2(n_1011),
.B(n_1318),
.Y(n_1475)
);

AOI221xp5_ASAP7_75t_SL g1476 ( 
.A1(n_1310),
.A2(n_1011),
.B1(n_1270),
.B2(n_1198),
.C(n_1322),
.Y(n_1476)
);

A2O1A1Ixp33_ASAP7_75t_L g1477 ( 
.A1(n_1261),
.A2(n_1011),
.B(n_881),
.C(n_1060),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1260),
.B(n_1060),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1326),
.B(n_973),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1326),
.B(n_973),
.Y(n_1480)
);

AO31x2_ASAP7_75t_L g1481 ( 
.A1(n_1163),
.A2(n_1201),
.A3(n_990),
.B(n_1263),
.Y(n_1481)
);

AOI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1186),
.A2(n_1011),
.B(n_1318),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1326),
.B(n_973),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1199),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1208),
.B(n_974),
.Y(n_1485)
);

CKINVDCx11_ASAP7_75t_R g1486 ( 
.A(n_1233),
.Y(n_1486)
);

AOI221xp5_ASAP7_75t_L g1487 ( 
.A1(n_1261),
.A2(n_1060),
.B1(n_881),
.B2(n_865),
.C(n_899),
.Y(n_1487)
);

A2O1A1Ixp33_ASAP7_75t_L g1488 ( 
.A1(n_1261),
.A2(n_1011),
.B(n_881),
.C(n_1060),
.Y(n_1488)
);

AO32x2_ASAP7_75t_L g1489 ( 
.A1(n_1198),
.A2(n_1310),
.A3(n_990),
.B1(n_1270),
.B2(n_1322),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1326),
.B(n_973),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_SL g1491 ( 
.A(n_1290),
.B(n_1011),
.Y(n_1491)
);

CKINVDCx20_ASAP7_75t_R g1492 ( 
.A(n_1225),
.Y(n_1492)
);

INVx2_ASAP7_75t_SL g1493 ( 
.A(n_1166),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1286),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1260),
.B(n_1060),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1326),
.B(n_973),
.Y(n_1496)
);

INVx6_ASAP7_75t_L g1497 ( 
.A(n_1343),
.Y(n_1497)
);

INVx6_ASAP7_75t_L g1498 ( 
.A(n_1343),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1330),
.Y(n_1499)
);

CKINVDCx11_ASAP7_75t_R g1500 ( 
.A(n_1492),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1487),
.A2(n_1440),
.B1(n_1473),
.B2(n_1471),
.Y(n_1501)
);

CKINVDCx20_ASAP7_75t_R g1502 ( 
.A(n_1333),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_SL g1503 ( 
.A1(n_1400),
.A2(n_1440),
.B1(n_1415),
.B2(n_1478),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1469),
.A2(n_1491),
.B1(n_1399),
.B2(n_1463),
.Y(n_1504)
);

BUFx8_ASAP7_75t_SL g1505 ( 
.A(n_1374),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1446),
.A2(n_1457),
.B1(n_1477),
.B2(n_1488),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1385),
.A2(n_1495),
.B1(n_1485),
.B2(n_1335),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1484),
.Y(n_1508)
);

OAI22xp33_ASAP7_75t_SL g1509 ( 
.A1(n_1369),
.A2(n_1399),
.B1(n_1367),
.B2(n_1496),
.Y(n_1509)
);

BUFx3_ASAP7_75t_L g1510 ( 
.A(n_1344),
.Y(n_1510)
);

CKINVDCx20_ASAP7_75t_R g1511 ( 
.A(n_1486),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1405),
.Y(n_1512)
);

BUFx3_ASAP7_75t_L g1513 ( 
.A(n_1405),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1329),
.A2(n_1367),
.B1(n_1369),
.B2(n_1347),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1329),
.A2(n_1474),
.B1(n_1461),
.B2(n_1439),
.Y(n_1515)
);

BUFx4_ASAP7_75t_SL g1516 ( 
.A(n_1378),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_1436),
.Y(n_1517)
);

OAI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1433),
.A2(n_1462),
.B1(n_1490),
.B2(n_1483),
.Y(n_1518)
);

CKINVDCx20_ASAP7_75t_R g1519 ( 
.A(n_1403),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1450),
.A2(n_1479),
.B1(n_1480),
.B2(n_1384),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1377),
.Y(n_1521)
);

INVx8_ASAP7_75t_L g1522 ( 
.A(n_1337),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1402),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1364),
.B(n_1383),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1375),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1404),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1340),
.Y(n_1527)
);

INVx6_ASAP7_75t_L g1528 ( 
.A(n_1380),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1375),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1461),
.A2(n_1474),
.B1(n_1418),
.B2(n_1422),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1376),
.A2(n_1366),
.B1(n_1338),
.B2(n_1379),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1494),
.Y(n_1532)
);

CKINVDCx20_ASAP7_75t_R g1533 ( 
.A(n_1380),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1382),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1395),
.Y(n_1535)
);

BUFx4f_ASAP7_75t_SL g1536 ( 
.A(n_1436),
.Y(n_1536)
);

CKINVDCx11_ASAP7_75t_R g1537 ( 
.A(n_1467),
.Y(n_1537)
);

CKINVDCx20_ASAP7_75t_R g1538 ( 
.A(n_1445),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1443),
.Y(n_1539)
);

CKINVDCx11_ASAP7_75t_R g1540 ( 
.A(n_1421),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1376),
.A2(n_1338),
.B1(n_1363),
.B2(n_1408),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_1365),
.Y(n_1542)
);

INVx4_ASAP7_75t_L g1543 ( 
.A(n_1370),
.Y(n_1543)
);

NAND2x1p5_ASAP7_75t_L g1544 ( 
.A(n_1435),
.B(n_1449),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1390),
.A2(n_1368),
.B1(n_1349),
.B2(n_1434),
.Y(n_1545)
);

NAND2x1p5_ASAP7_75t_L g1546 ( 
.A(n_1358),
.B(n_1425),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1394),
.B(n_1493),
.Y(n_1547)
);

CKINVDCx11_ASAP7_75t_R g1548 ( 
.A(n_1368),
.Y(n_1548)
);

CKINVDCx11_ASAP7_75t_R g1549 ( 
.A(n_1456),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1424),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1398),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1434),
.A2(n_1476),
.B1(n_1387),
.B2(n_1389),
.Y(n_1552)
);

CKINVDCx20_ASAP7_75t_R g1553 ( 
.A(n_1452),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1476),
.A2(n_1387),
.B1(n_1361),
.B2(n_1443),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1429),
.Y(n_1555)
);

INVxp67_ASAP7_75t_SL g1556 ( 
.A(n_1417),
.Y(n_1556)
);

AOI22xp5_ASAP7_75t_SL g1557 ( 
.A1(n_1456),
.A2(n_1331),
.B1(n_1444),
.B2(n_1381),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1428),
.Y(n_1558)
);

BUFx6f_ASAP7_75t_L g1559 ( 
.A(n_1370),
.Y(n_1559)
);

CKINVDCx20_ASAP7_75t_R g1560 ( 
.A(n_1430),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1417),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1361),
.A2(n_1453),
.B1(n_1482),
.B2(n_1475),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_SL g1563 ( 
.A1(n_1332),
.A2(n_1423),
.B1(n_1489),
.B2(n_1432),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1426),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1373),
.B(n_1419),
.Y(n_1565)
);

AOI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1332),
.A2(n_1391),
.B1(n_1414),
.B2(n_1411),
.Y(n_1566)
);

BUFx3_ASAP7_75t_L g1567 ( 
.A(n_1420),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_SL g1568 ( 
.A1(n_1489),
.A2(n_1432),
.B1(n_1451),
.B2(n_1448),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_SL g1569 ( 
.A1(n_1489),
.A2(n_1454),
.B1(n_1447),
.B2(n_1464),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1406),
.A2(n_1348),
.B1(n_1401),
.B2(n_1337),
.Y(n_1570)
);

BUFx2_ASAP7_75t_L g1571 ( 
.A(n_1465),
.Y(n_1571)
);

BUFx2_ASAP7_75t_SL g1572 ( 
.A(n_1442),
.Y(n_1572)
);

INVx2_ASAP7_75t_SL g1573 ( 
.A(n_1442),
.Y(n_1573)
);

OAI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1407),
.A2(n_1348),
.B1(n_1437),
.B2(n_1353),
.Y(n_1574)
);

INVx1_ASAP7_75t_SL g1575 ( 
.A(n_1430),
.Y(n_1575)
);

BUFx8_ASAP7_75t_L g1576 ( 
.A(n_1442),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_SL g1577 ( 
.A1(n_1441),
.A2(n_1393),
.B1(n_1371),
.B2(n_1362),
.Y(n_1577)
);

INVx3_ASAP7_75t_L g1578 ( 
.A(n_1337),
.Y(n_1578)
);

BUFx3_ASAP7_75t_L g1579 ( 
.A(n_1466),
.Y(n_1579)
);

INVx3_ASAP7_75t_L g1580 ( 
.A(n_1466),
.Y(n_1580)
);

INVx6_ASAP7_75t_L g1581 ( 
.A(n_1466),
.Y(n_1581)
);

INVx1_ASAP7_75t_SL g1582 ( 
.A(n_1431),
.Y(n_1582)
);

AOI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1455),
.A2(n_1470),
.B1(n_1353),
.B2(n_1397),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1375),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1412),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1356),
.A2(n_1396),
.B1(n_1357),
.B2(n_1352),
.Y(n_1586)
);

CKINVDCx11_ASAP7_75t_R g1587 ( 
.A(n_1372),
.Y(n_1587)
);

BUFx10_ASAP7_75t_L g1588 ( 
.A(n_1438),
.Y(n_1588)
);

CKINVDCx20_ASAP7_75t_R g1589 ( 
.A(n_1427),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1459),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_SL g1591 ( 
.A1(n_1357),
.A2(n_1413),
.B1(n_1409),
.B2(n_1352),
.Y(n_1591)
);

AOI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1341),
.A2(n_1342),
.B1(n_1416),
.B2(n_1339),
.Y(n_1592)
);

CKINVDCx20_ASAP7_75t_R g1593 ( 
.A(n_1388),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1388),
.B(n_1460),
.Y(n_1594)
);

AOI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1410),
.A2(n_1392),
.B1(n_1360),
.B2(n_1359),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1351),
.A2(n_1336),
.B1(n_1481),
.B2(n_1472),
.Y(n_1596)
);

NAND2x1p5_ASAP7_75t_L g1597 ( 
.A(n_1350),
.B(n_1458),
.Y(n_1597)
);

CKINVDCx11_ASAP7_75t_R g1598 ( 
.A(n_1388),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1460),
.B(n_1481),
.Y(n_1599)
);

INVx6_ASAP7_75t_L g1600 ( 
.A(n_1354),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1354),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_SL g1602 ( 
.A1(n_1355),
.A2(n_1468),
.B1(n_1472),
.B2(n_1481),
.Y(n_1602)
);

CKINVDCx11_ASAP7_75t_R g1603 ( 
.A(n_1334),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1345),
.A2(n_1355),
.B1(n_1346),
.B2(n_1354),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1355),
.A2(n_1487),
.B1(n_1440),
.B2(n_1473),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1330),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1485),
.B(n_1208),
.Y(n_1607)
);

CKINVDCx6p67_ASAP7_75t_R g1608 ( 
.A(n_1344),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1330),
.Y(n_1609)
);

BUFx6f_ASAP7_75t_L g1610 ( 
.A(n_1370),
.Y(n_1610)
);

CKINVDCx11_ASAP7_75t_R g1611 ( 
.A(n_1492),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1344),
.Y(n_1612)
);

AOI22x1_ASAP7_75t_L g1613 ( 
.A1(n_1463),
.A2(n_1329),
.B1(n_1290),
.B2(n_1389),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_SL g1614 ( 
.A1(n_1400),
.A2(n_1060),
.B1(n_775),
.B2(n_729),
.Y(n_1614)
);

INVx6_ASAP7_75t_L g1615 ( 
.A(n_1343),
.Y(n_1615)
);

BUFx3_ASAP7_75t_L g1616 ( 
.A(n_1344),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1487),
.A2(n_1440),
.B1(n_1473),
.B2(n_1471),
.Y(n_1617)
);

INVx6_ASAP7_75t_L g1618 ( 
.A(n_1343),
.Y(n_1618)
);

OAI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1473),
.A2(n_1011),
.B1(n_1487),
.B2(n_1457),
.Y(n_1619)
);

AO22x1_ASAP7_75t_L g1620 ( 
.A1(n_1367),
.A2(n_973),
.B1(n_1060),
.B2(n_1261),
.Y(n_1620)
);

BUFx3_ASAP7_75t_L g1621 ( 
.A(n_1344),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_SL g1622 ( 
.A1(n_1400),
.A2(n_1060),
.B1(n_775),
.B2(n_729),
.Y(n_1622)
);

INVx1_ASAP7_75t_SL g1623 ( 
.A(n_1445),
.Y(n_1623)
);

BUFx10_ASAP7_75t_L g1624 ( 
.A(n_1333),
.Y(n_1624)
);

BUFx12f_ASAP7_75t_L g1625 ( 
.A(n_1486),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1487),
.A2(n_1440),
.B1(n_1473),
.B2(n_1471),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1330),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1330),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1330),
.Y(n_1629)
);

CKINVDCx6p67_ASAP7_75t_R g1630 ( 
.A(n_1344),
.Y(n_1630)
);

BUFx12f_ASAP7_75t_L g1631 ( 
.A(n_1486),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1487),
.A2(n_1440),
.B1(n_1473),
.B2(n_1471),
.Y(n_1632)
);

OAI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1473),
.A2(n_1011),
.B1(n_1487),
.B2(n_1457),
.Y(n_1633)
);

CKINVDCx20_ASAP7_75t_R g1634 ( 
.A(n_1492),
.Y(n_1634)
);

INVx8_ASAP7_75t_L g1635 ( 
.A(n_1337),
.Y(n_1635)
);

BUFx8_ASAP7_75t_SL g1636 ( 
.A(n_1492),
.Y(n_1636)
);

OAI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1473),
.A2(n_1011),
.B1(n_1487),
.B2(n_1457),
.Y(n_1637)
);

BUFx2_ASAP7_75t_SL g1638 ( 
.A(n_1492),
.Y(n_1638)
);

INVx8_ASAP7_75t_L g1639 ( 
.A(n_1337),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1330),
.Y(n_1640)
);

INVx3_ASAP7_75t_L g1641 ( 
.A(n_1435),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1330),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_SL g1643 ( 
.A1(n_1400),
.A2(n_1060),
.B1(n_775),
.B2(n_729),
.Y(n_1643)
);

INVx3_ASAP7_75t_L g1644 ( 
.A(n_1435),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1330),
.Y(n_1645)
);

INVx3_ASAP7_75t_L g1646 ( 
.A(n_1435),
.Y(n_1646)
);

OAI21xp5_ASAP7_75t_SL g1647 ( 
.A1(n_1473),
.A2(n_1060),
.B(n_682),
.Y(n_1647)
);

AOI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1441),
.A2(n_1448),
.B(n_1447),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1330),
.Y(n_1649)
);

BUFx5_ASAP7_75t_L g1650 ( 
.A(n_1386),
.Y(n_1650)
);

INVx2_ASAP7_75t_SL g1651 ( 
.A(n_1344),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1473),
.A2(n_1011),
.B1(n_1487),
.B2(n_1457),
.Y(n_1652)
);

INVx6_ASAP7_75t_L g1653 ( 
.A(n_1343),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1330),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1330),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1485),
.B(n_1208),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1584),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1539),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1564),
.Y(n_1659)
);

BUFx2_ASAP7_75t_SL g1660 ( 
.A(n_1589),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1539),
.Y(n_1661)
);

INVxp67_ASAP7_75t_L g1662 ( 
.A(n_1547),
.Y(n_1662)
);

BUFx12f_ASAP7_75t_L g1663 ( 
.A(n_1500),
.Y(n_1663)
);

BUFx3_ASAP7_75t_L g1664 ( 
.A(n_1522),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1594),
.B(n_1515),
.Y(n_1665)
);

INVx4_ASAP7_75t_SL g1666 ( 
.A(n_1600),
.Y(n_1666)
);

OAI21xp33_ASAP7_75t_SL g1667 ( 
.A1(n_1530),
.A2(n_1583),
.B(n_1501),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1647),
.B(n_1538),
.Y(n_1668)
);

NAND2x1p5_ASAP7_75t_L g1669 ( 
.A(n_1566),
.B(n_1641),
.Y(n_1669)
);

INVx3_ASAP7_75t_L g1670 ( 
.A(n_1546),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1515),
.B(n_1593),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1605),
.B(n_1556),
.Y(n_1672)
);

BUFx3_ASAP7_75t_L g1673 ( 
.A(n_1522),
.Y(n_1673)
);

OAI21x1_ASAP7_75t_L g1674 ( 
.A1(n_1648),
.A2(n_1597),
.B(n_1595),
.Y(n_1674)
);

BUFx6f_ASAP7_75t_L g1675 ( 
.A(n_1600),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1599),
.B(n_1590),
.Y(n_1676)
);

AOI21xp33_ASAP7_75t_L g1677 ( 
.A1(n_1619),
.A2(n_1637),
.B(n_1633),
.Y(n_1677)
);

AO21x2_ASAP7_75t_L g1678 ( 
.A1(n_1574),
.A2(n_1592),
.B(n_1604),
.Y(n_1678)
);

AND2x4_ASAP7_75t_L g1679 ( 
.A(n_1585),
.B(n_1578),
.Y(n_1679)
);

OA21x2_ASAP7_75t_L g1680 ( 
.A1(n_1596),
.A2(n_1562),
.B(n_1586),
.Y(n_1680)
);

INVxp67_ASAP7_75t_SL g1681 ( 
.A(n_1524),
.Y(n_1681)
);

BUFx3_ASAP7_75t_L g1682 ( 
.A(n_1522),
.Y(n_1682)
);

CKINVDCx20_ASAP7_75t_R g1683 ( 
.A(n_1505),
.Y(n_1683)
);

AOI21x1_ASAP7_75t_L g1684 ( 
.A1(n_1525),
.A2(n_1529),
.B(n_1620),
.Y(n_1684)
);

INVx1_ASAP7_75t_SL g1685 ( 
.A(n_1542),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1525),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1529),
.Y(n_1687)
);

OAI21x1_ASAP7_75t_L g1688 ( 
.A1(n_1597),
.A2(n_1601),
.B(n_1562),
.Y(n_1688)
);

INVx3_ASAP7_75t_L g1689 ( 
.A(n_1546),
.Y(n_1689)
);

AOI22xp33_ASAP7_75t_L g1690 ( 
.A1(n_1587),
.A2(n_1530),
.B1(n_1614),
.B2(n_1622),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1605),
.B(n_1556),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1563),
.B(n_1598),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1598),
.B(n_1504),
.Y(n_1693)
);

INVx3_ASAP7_75t_L g1694 ( 
.A(n_1600),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1504),
.B(n_1602),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1503),
.B(n_1603),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1561),
.B(n_1545),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1650),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_1636),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1650),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1643),
.A2(n_1626),
.B1(n_1632),
.B2(n_1501),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1650),
.Y(n_1702)
);

BUFx2_ASAP7_75t_L g1703 ( 
.A(n_1650),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1520),
.B(n_1623),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1650),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1578),
.B(n_1644),
.Y(n_1706)
);

INVx4_ASAP7_75t_L g1707 ( 
.A(n_1635),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1508),
.Y(n_1708)
);

OAI21x1_ASAP7_75t_L g1709 ( 
.A1(n_1601),
.A2(n_1586),
.B(n_1596),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1526),
.B(n_1628),
.Y(n_1710)
);

INVx2_ASAP7_75t_SL g1711 ( 
.A(n_1635),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1545),
.B(n_1552),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1628),
.Y(n_1713)
);

AOI21x1_ASAP7_75t_L g1714 ( 
.A1(n_1506),
.A2(n_1652),
.B(n_1570),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1617),
.A2(n_1632),
.B1(n_1626),
.B2(n_1509),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1640),
.Y(n_1716)
);

BUFx2_ASAP7_75t_L g1717 ( 
.A(n_1649),
.Y(n_1717)
);

BUFx3_ASAP7_75t_L g1718 ( 
.A(n_1635),
.Y(n_1718)
);

OAI21x1_ASAP7_75t_L g1719 ( 
.A1(n_1646),
.A2(n_1554),
.B(n_1544),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1617),
.A2(n_1613),
.B1(n_1514),
.B2(n_1607),
.Y(n_1720)
);

AO21x1_ASAP7_75t_L g1721 ( 
.A1(n_1574),
.A2(n_1518),
.B(n_1565),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1552),
.B(n_1554),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1655),
.Y(n_1723)
);

BUFx2_ASAP7_75t_L g1724 ( 
.A(n_1499),
.Y(n_1724)
);

OAI21x1_ASAP7_75t_L g1725 ( 
.A1(n_1544),
.A2(n_1541),
.B(n_1531),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1568),
.B(n_1569),
.Y(n_1726)
);

INVx2_ASAP7_75t_SL g1727 ( 
.A(n_1639),
.Y(n_1727)
);

INVx2_ASAP7_75t_SL g1728 ( 
.A(n_1639),
.Y(n_1728)
);

INVx3_ASAP7_75t_L g1729 ( 
.A(n_1588),
.Y(n_1729)
);

BUFx2_ASAP7_75t_SL g1730 ( 
.A(n_1533),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1523),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1606),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1609),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1627),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1629),
.Y(n_1735)
);

OAI21x1_ASAP7_75t_L g1736 ( 
.A1(n_1541),
.A2(n_1531),
.B(n_1654),
.Y(n_1736)
);

INVx1_ASAP7_75t_SL g1737 ( 
.A(n_1560),
.Y(n_1737)
);

AOI21x1_ASAP7_75t_L g1738 ( 
.A1(n_1642),
.A2(n_1645),
.B(n_1555),
.Y(n_1738)
);

BUFx4f_ASAP7_75t_L g1739 ( 
.A(n_1639),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1558),
.B(n_1514),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1575),
.Y(n_1741)
);

BUFx2_ASAP7_75t_L g1742 ( 
.A(n_1571),
.Y(n_1742)
);

BUFx8_ASAP7_75t_L g1743 ( 
.A(n_1625),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1591),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1534),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1535),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1527),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1532),
.B(n_1550),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1588),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1559),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1518),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_1611),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1507),
.B(n_1656),
.Y(n_1753)
);

OAI21x1_ASAP7_75t_L g1754 ( 
.A1(n_1577),
.A2(n_1580),
.B(n_1557),
.Y(n_1754)
);

NOR2x1_ASAP7_75t_SL g1755 ( 
.A(n_1572),
.B(n_1610),
.Y(n_1755)
);

INVx2_ASAP7_75t_SL g1756 ( 
.A(n_1497),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1582),
.B(n_1513),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1512),
.B(n_1513),
.Y(n_1758)
);

INVx2_ASAP7_75t_SL g1759 ( 
.A(n_1497),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1512),
.B(n_1580),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1559),
.B(n_1610),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1553),
.B(n_1634),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1567),
.Y(n_1763)
);

BUFx3_ASAP7_75t_L g1764 ( 
.A(n_1576),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1567),
.Y(n_1765)
);

AND2x4_ASAP7_75t_L g1766 ( 
.A(n_1579),
.B(n_1621),
.Y(n_1766)
);

BUFx2_ASAP7_75t_L g1767 ( 
.A(n_1551),
.Y(n_1767)
);

BUFx3_ASAP7_75t_L g1768 ( 
.A(n_1576),
.Y(n_1768)
);

BUFx2_ASAP7_75t_L g1769 ( 
.A(n_1521),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1638),
.B(n_1612),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1581),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1498),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1498),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1498),
.Y(n_1774)
);

OA21x2_ASAP7_75t_L g1775 ( 
.A1(n_1573),
.A2(n_1651),
.B(n_1517),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1757),
.B(n_1621),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1757),
.B(n_1616),
.Y(n_1777)
);

O2A1O1Ixp33_ASAP7_75t_L g1778 ( 
.A1(n_1677),
.A2(n_1510),
.B(n_1519),
.C(n_1511),
.Y(n_1778)
);

CKINVDCx10_ASAP7_75t_R g1779 ( 
.A(n_1743),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1693),
.B(n_1510),
.Y(n_1780)
);

OAI21x1_ASAP7_75t_SL g1781 ( 
.A1(n_1714),
.A2(n_1543),
.B(n_1516),
.Y(n_1781)
);

OR2x6_ASAP7_75t_L g1782 ( 
.A(n_1725),
.B(n_1669),
.Y(n_1782)
);

AOI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1690),
.A2(n_1537),
.B1(n_1548),
.B2(n_1549),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1693),
.B(n_1608),
.Y(n_1784)
);

BUFx3_ASAP7_75t_L g1785 ( 
.A(n_1766),
.Y(n_1785)
);

OA21x2_ASAP7_75t_L g1786 ( 
.A1(n_1709),
.A2(n_1615),
.B(n_1618),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1692),
.B(n_1630),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1679),
.B(n_1502),
.Y(n_1788)
);

OAI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1701),
.A2(n_1615),
.B1(n_1528),
.B2(n_1618),
.Y(n_1789)
);

A2O1A1Ixp33_ASAP7_75t_L g1790 ( 
.A1(n_1667),
.A2(n_1615),
.B(n_1528),
.C(n_1618),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_L g1791 ( 
.A(n_1667),
.B(n_1653),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1724),
.Y(n_1792)
);

A2O1A1Ixp33_ASAP7_75t_L g1793 ( 
.A1(n_1715),
.A2(n_1696),
.B(n_1725),
.C(n_1720),
.Y(n_1793)
);

OR2x6_ASAP7_75t_L g1794 ( 
.A(n_1669),
.B(n_1653),
.Y(n_1794)
);

AND2x4_ASAP7_75t_L g1795 ( 
.A(n_1679),
.B(n_1540),
.Y(n_1795)
);

OAI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1714),
.A2(n_1736),
.B(n_1751),
.Y(n_1796)
);

OAI21x1_ASAP7_75t_L g1797 ( 
.A1(n_1674),
.A2(n_1536),
.B(n_1624),
.Y(n_1797)
);

AOI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1696),
.A2(n_1631),
.B1(n_1536),
.B2(n_1624),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1686),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1738),
.Y(n_1800)
);

HB1xp67_ASAP7_75t_L g1801 ( 
.A(n_1686),
.Y(n_1801)
);

AO21x2_ASAP7_75t_L g1802 ( 
.A1(n_1721),
.A2(n_1684),
.B(n_1751),
.Y(n_1802)
);

AOI21xp5_ASAP7_75t_L g1803 ( 
.A1(n_1678),
.A2(n_1681),
.B(n_1680),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1692),
.B(n_1671),
.Y(n_1804)
);

AOI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1660),
.A2(n_1668),
.B1(n_1721),
.B2(n_1753),
.Y(n_1805)
);

AOI22xp33_ASAP7_75t_L g1806 ( 
.A1(n_1671),
.A2(n_1704),
.B1(n_1726),
.B2(n_1678),
.Y(n_1806)
);

O2A1O1Ixp33_ASAP7_75t_L g1807 ( 
.A1(n_1744),
.A2(n_1741),
.B(n_1678),
.C(n_1726),
.Y(n_1807)
);

A2O1A1Ixp33_ASAP7_75t_L g1808 ( 
.A1(n_1736),
.A2(n_1695),
.B(n_1744),
.C(n_1712),
.Y(n_1808)
);

CKINVDCx5p33_ASAP7_75t_R g1809 ( 
.A(n_1699),
.Y(n_1809)
);

AOI221xp5_ASAP7_75t_L g1810 ( 
.A1(n_1695),
.A2(n_1691),
.B1(n_1672),
.B2(n_1662),
.C(n_1740),
.Y(n_1810)
);

NOR2x1_ASAP7_75t_SL g1811 ( 
.A(n_1660),
.B(n_1675),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1672),
.B(n_1691),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1738),
.Y(n_1813)
);

OAI211xp5_ASAP7_75t_L g1814 ( 
.A1(n_1712),
.A2(n_1740),
.B(n_1684),
.C(n_1722),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1665),
.B(n_1710),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1697),
.B(n_1717),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1717),
.B(n_1713),
.Y(n_1817)
);

OAI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1669),
.A2(n_1749),
.B(n_1754),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1685),
.B(n_1737),
.Y(n_1819)
);

A2O1A1Ixp33_ASAP7_75t_L g1820 ( 
.A1(n_1739),
.A2(n_1722),
.B(n_1754),
.C(n_1768),
.Y(n_1820)
);

AOI22xp5_ASAP7_75t_SL g1821 ( 
.A1(n_1730),
.A2(n_1752),
.B1(n_1764),
.B2(n_1768),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_L g1822 ( 
.A(n_1770),
.B(n_1762),
.Y(n_1822)
);

OAI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1764),
.A2(n_1768),
.B1(n_1739),
.B2(n_1769),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1713),
.B(n_1716),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1767),
.B(n_1769),
.Y(n_1825)
);

NOR2xp33_ASAP7_75t_L g1826 ( 
.A(n_1770),
.B(n_1730),
.Y(n_1826)
);

AOI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1680),
.A2(n_1674),
.B(n_1688),
.Y(n_1827)
);

OAI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1749),
.A2(n_1680),
.B(n_1729),
.Y(n_1828)
);

O2A1O1Ixp33_ASAP7_75t_L g1829 ( 
.A1(n_1767),
.A2(n_1749),
.B(n_1774),
.C(n_1773),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1742),
.B(n_1758),
.Y(n_1830)
);

OA21x2_ASAP7_75t_L g1831 ( 
.A1(n_1719),
.A2(n_1657),
.B(n_1687),
.Y(n_1831)
);

AND2x4_ASAP7_75t_SL g1832 ( 
.A(n_1766),
.B(n_1683),
.Y(n_1832)
);

AOI22xp33_ASAP7_75t_L g1833 ( 
.A1(n_1663),
.A2(n_1680),
.B1(n_1743),
.B2(n_1748),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1758),
.B(n_1763),
.Y(n_1834)
);

AND2x4_ASAP7_75t_L g1835 ( 
.A(n_1679),
.B(n_1706),
.Y(n_1835)
);

NAND2xp33_ASAP7_75t_R g1836 ( 
.A(n_1766),
.B(n_1775),
.Y(n_1836)
);

OA21x2_ASAP7_75t_L g1837 ( 
.A1(n_1657),
.A2(n_1687),
.B(n_1698),
.Y(n_1837)
);

NOR2x1_ASAP7_75t_SL g1838 ( 
.A(n_1675),
.B(n_1698),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1679),
.B(n_1706),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1765),
.B(n_1761),
.Y(n_1840)
);

NAND4xp25_ASAP7_75t_L g1841 ( 
.A(n_1745),
.B(n_1734),
.C(n_1732),
.D(n_1733),
.Y(n_1841)
);

BUFx12f_ASAP7_75t_L g1842 ( 
.A(n_1663),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1761),
.B(n_1760),
.Y(n_1843)
);

OAI221xp5_ASAP7_75t_L g1844 ( 
.A1(n_1739),
.A2(n_1727),
.B1(n_1711),
.B2(n_1728),
.C(n_1764),
.Y(n_1844)
);

CKINVDCx20_ASAP7_75t_R g1845 ( 
.A(n_1743),
.Y(n_1845)
);

AO32x2_ASAP7_75t_L g1846 ( 
.A1(n_1711),
.A2(n_1727),
.A3(n_1728),
.B1(n_1759),
.B2(n_1756),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1731),
.B(n_1733),
.Y(n_1847)
);

NAND2xp33_ASAP7_75t_L g1848 ( 
.A(n_1756),
.B(n_1759),
.Y(n_1848)
);

AND2x4_ASAP7_75t_L g1849 ( 
.A(n_1706),
.B(n_1666),
.Y(n_1849)
);

NAND4xp25_ASAP7_75t_L g1850 ( 
.A(n_1735),
.B(n_1746),
.C(n_1747),
.D(n_1723),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1775),
.B(n_1750),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1799),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1799),
.Y(n_1853)
);

BUFx3_ASAP7_75t_L g1854 ( 
.A(n_1842),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1815),
.B(n_1851),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1801),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1840),
.B(n_1703),
.Y(n_1857)
);

INVx3_ASAP7_75t_L g1858 ( 
.A(n_1835),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1834),
.B(n_1700),
.Y(n_1859)
);

INVxp67_ASAP7_75t_L g1860 ( 
.A(n_1825),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1837),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1801),
.Y(n_1862)
);

OAI21xp5_ASAP7_75t_SL g1863 ( 
.A1(n_1805),
.A2(n_1772),
.B(n_1743),
.Y(n_1863)
);

AND2x4_ASAP7_75t_L g1864 ( 
.A(n_1835),
.B(n_1706),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1816),
.B(n_1676),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1812),
.B(n_1658),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1812),
.B(n_1700),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1839),
.B(n_1702),
.Y(n_1868)
);

INVx3_ASAP7_75t_L g1869 ( 
.A(n_1839),
.Y(n_1869)
);

BUFx2_ASAP7_75t_L g1870 ( 
.A(n_1846),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1843),
.B(n_1702),
.Y(n_1871)
);

AOI21xp5_ASAP7_75t_SL g1872 ( 
.A1(n_1790),
.A2(n_1755),
.B(n_1775),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1800),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1813),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1810),
.B(n_1708),
.Y(n_1875)
);

HB1xp67_ASAP7_75t_L g1876 ( 
.A(n_1792),
.Y(n_1876)
);

AOI22xp33_ASAP7_75t_L g1877 ( 
.A1(n_1806),
.A2(n_1707),
.B1(n_1682),
.B2(n_1664),
.Y(n_1877)
);

AND2x2_ASAP7_75t_SL g1878 ( 
.A(n_1806),
.B(n_1675),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1817),
.B(n_1661),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1810),
.B(n_1708),
.Y(n_1880)
);

OAI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1793),
.A2(n_1682),
.B1(n_1673),
.B2(n_1718),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1817),
.B(n_1661),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1847),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1791),
.A2(n_1707),
.B1(n_1664),
.B2(n_1718),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1804),
.B(n_1830),
.Y(n_1885)
);

OAI221xp5_ASAP7_75t_SL g1886 ( 
.A1(n_1807),
.A2(n_1673),
.B1(n_1682),
.B2(n_1718),
.C(n_1664),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1828),
.B(n_1705),
.Y(n_1887)
);

AND2x4_ASAP7_75t_L g1888 ( 
.A(n_1849),
.B(n_1785),
.Y(n_1888)
);

AND2x4_ASAP7_75t_L g1889 ( 
.A(n_1849),
.B(n_1689),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1824),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1824),
.Y(n_1891)
);

BUFx2_ASAP7_75t_L g1892 ( 
.A(n_1846),
.Y(n_1892)
);

AOI22xp33_ASAP7_75t_L g1893 ( 
.A1(n_1791),
.A2(n_1826),
.B1(n_1789),
.B2(n_1822),
.Y(n_1893)
);

OR2x2_ASAP7_75t_L g1894 ( 
.A(n_1803),
.B(n_1659),
.Y(n_1894)
);

BUFx2_ASAP7_75t_L g1895 ( 
.A(n_1846),
.Y(n_1895)
);

AOI22xp5_ASAP7_75t_L g1896 ( 
.A1(n_1789),
.A2(n_1707),
.B1(n_1673),
.B2(n_1694),
.Y(n_1896)
);

INVxp67_ASAP7_75t_SL g1897 ( 
.A(n_1829),
.Y(n_1897)
);

AOI22xp33_ASAP7_75t_L g1898 ( 
.A1(n_1780),
.A2(n_1694),
.B1(n_1689),
.B2(n_1670),
.Y(n_1898)
);

AND2x4_ASAP7_75t_L g1899 ( 
.A(n_1887),
.B(n_1838),
.Y(n_1899)
);

INVx4_ASAP7_75t_L g1900 ( 
.A(n_1854),
.Y(n_1900)
);

BUFx2_ASAP7_75t_L g1901 ( 
.A(n_1870),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1855),
.B(n_1782),
.Y(n_1902)
);

OR2x2_ASAP7_75t_L g1903 ( 
.A(n_1865),
.B(n_1803),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1867),
.B(n_1802),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1873),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1867),
.B(n_1802),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1870),
.B(n_1782),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1873),
.Y(n_1908)
);

INVx3_ASAP7_75t_L g1909 ( 
.A(n_1861),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1868),
.B(n_1786),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1887),
.B(n_1797),
.Y(n_1911)
);

INVx1_ASAP7_75t_SL g1912 ( 
.A(n_1865),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1874),
.Y(n_1913)
);

INVx4_ASAP7_75t_L g1914 ( 
.A(n_1854),
.Y(n_1914)
);

OR2x2_ASAP7_75t_L g1915 ( 
.A(n_1866),
.B(n_1828),
.Y(n_1915)
);

AOI22xp33_ASAP7_75t_SL g1916 ( 
.A1(n_1878),
.A2(n_1814),
.B1(n_1821),
.B2(n_1811),
.Y(n_1916)
);

AO21x2_ASAP7_75t_L g1917 ( 
.A1(n_1897),
.A2(n_1827),
.B(n_1818),
.Y(n_1917)
);

AOI21xp5_ASAP7_75t_L g1918 ( 
.A1(n_1872),
.A2(n_1807),
.B(n_1827),
.Y(n_1918)
);

AO21x2_ASAP7_75t_L g1919 ( 
.A1(n_1894),
.A2(n_1818),
.B(n_1796),
.Y(n_1919)
);

NAND3xp33_ASAP7_75t_L g1920 ( 
.A(n_1893),
.B(n_1814),
.C(n_1808),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1858),
.B(n_1833),
.Y(n_1921)
);

INVxp67_ASAP7_75t_L g1922 ( 
.A(n_1852),
.Y(n_1922)
);

INVx1_ASAP7_75t_SL g1923 ( 
.A(n_1879),
.Y(n_1923)
);

BUFx2_ASAP7_75t_L g1924 ( 
.A(n_1892),
.Y(n_1924)
);

OAI21xp5_ASAP7_75t_L g1925 ( 
.A1(n_1881),
.A2(n_1820),
.B(n_1833),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1892),
.B(n_1831),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1852),
.Y(n_1927)
);

AOI221x1_ASAP7_75t_L g1928 ( 
.A1(n_1872),
.A2(n_1841),
.B1(n_1823),
.B2(n_1850),
.C(n_1781),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1853),
.Y(n_1929)
);

CKINVDCx5p33_ASAP7_75t_R g1930 ( 
.A(n_1860),
.Y(n_1930)
);

OAI21xp33_ASAP7_75t_L g1931 ( 
.A1(n_1878),
.A2(n_1863),
.B(n_1886),
.Y(n_1931)
);

AND2x4_ASAP7_75t_L g1932 ( 
.A(n_1869),
.B(n_1795),
.Y(n_1932)
);

OR2x2_ASAP7_75t_L g1933 ( 
.A(n_1895),
.B(n_1796),
.Y(n_1933)
);

AOI21xp5_ASAP7_75t_L g1934 ( 
.A1(n_1894),
.A2(n_1829),
.B(n_1848),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1885),
.B(n_1776),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1885),
.B(n_1777),
.Y(n_1936)
);

INVx3_ASAP7_75t_L g1937 ( 
.A(n_1864),
.Y(n_1937)
);

INVx3_ASAP7_75t_L g1938 ( 
.A(n_1864),
.Y(n_1938)
);

BUFx2_ASAP7_75t_L g1939 ( 
.A(n_1864),
.Y(n_1939)
);

HB1xp67_ASAP7_75t_L g1940 ( 
.A(n_1856),
.Y(n_1940)
);

AOI22xp33_ASAP7_75t_L g1941 ( 
.A1(n_1877),
.A2(n_1783),
.B1(n_1795),
.B2(n_1788),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1901),
.B(n_1883),
.Y(n_1942)
);

NOR2xp67_ASAP7_75t_SL g1943 ( 
.A(n_1920),
.B(n_1844),
.Y(n_1943)
);

BUFx3_ASAP7_75t_L g1944 ( 
.A(n_1900),
.Y(n_1944)
);

NAND2xp33_ASAP7_75t_R g1945 ( 
.A(n_1918),
.B(n_1809),
.Y(n_1945)
);

INVx1_ASAP7_75t_SL g1946 ( 
.A(n_1912),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1937),
.B(n_1871),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1904),
.B(n_1876),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1937),
.B(n_1871),
.Y(n_1949)
);

NOR2xp33_ASAP7_75t_L g1950 ( 
.A(n_1900),
.B(n_1787),
.Y(n_1950)
);

INVxp67_ASAP7_75t_L g1951 ( 
.A(n_1940),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1937),
.B(n_1889),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1909),
.Y(n_1953)
);

BUFx2_ASAP7_75t_L g1954 ( 
.A(n_1939),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1937),
.B(n_1889),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1938),
.B(n_1889),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1905),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1905),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_SL g1959 ( 
.A(n_1916),
.B(n_1788),
.Y(n_1959)
);

OR2x6_ASAP7_75t_L g1960 ( 
.A(n_1918),
.B(n_1934),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1939),
.B(n_1907),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1904),
.B(n_1882),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1908),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1909),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1908),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1913),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1907),
.B(n_1859),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1913),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1907),
.B(n_1857),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1906),
.B(n_1890),
.Y(n_1970)
);

OAI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1920),
.A2(n_1896),
.B1(n_1884),
.B2(n_1798),
.Y(n_1971)
);

BUFx2_ASAP7_75t_L g1972 ( 
.A(n_1899),
.Y(n_1972)
);

AOI22xp33_ASAP7_75t_L g1973 ( 
.A1(n_1931),
.A2(n_1880),
.B1(n_1875),
.B2(n_1784),
.Y(n_1973)
);

INVx3_ASAP7_75t_R g1974 ( 
.A(n_1932),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1940),
.Y(n_1975)
);

NOR2xp67_ASAP7_75t_L g1976 ( 
.A(n_1934),
.B(n_1862),
.Y(n_1976)
);

NAND2xp67_ASAP7_75t_L g1977 ( 
.A(n_1921),
.B(n_1832),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1927),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1927),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1906),
.B(n_1890),
.Y(n_1980)
);

OR2x2_ASAP7_75t_L g1981 ( 
.A(n_1933),
.B(n_1882),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1922),
.B(n_1891),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1922),
.B(n_1891),
.Y(n_1983)
);

CKINVDCx20_ASAP7_75t_R g1984 ( 
.A(n_1930),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1910),
.B(n_1888),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1910),
.B(n_1888),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1901),
.B(n_1888),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1929),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1953),
.Y(n_1989)
);

OR2x2_ASAP7_75t_L g1990 ( 
.A(n_1948),
.B(n_1981),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1957),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1973),
.B(n_1912),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1957),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1961),
.B(n_1924),
.Y(n_1994)
);

INVx2_ASAP7_75t_SL g1995 ( 
.A(n_1987),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1958),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1958),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1973),
.B(n_1943),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1961),
.B(n_1924),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1963),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1972),
.B(n_1899),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1963),
.Y(n_2002)
);

NAND2x1_ASAP7_75t_L g2003 ( 
.A(n_1960),
.B(n_1899),
.Y(n_2003)
);

NAND2x1p5_ASAP7_75t_L g2004 ( 
.A(n_1976),
.B(n_1900),
.Y(n_2004)
);

OR2x6_ASAP7_75t_L g2005 ( 
.A(n_1960),
.B(n_1959),
.Y(n_2005)
);

HB1xp67_ASAP7_75t_L g2006 ( 
.A(n_1946),
.Y(n_2006)
);

INVxp67_ASAP7_75t_L g2007 ( 
.A(n_1943),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1965),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1972),
.B(n_1952),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1965),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1966),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1966),
.Y(n_2012)
);

AOI211xp5_ASAP7_75t_L g2013 ( 
.A1(n_1971),
.A2(n_1931),
.B(n_1925),
.C(n_1778),
.Y(n_2013)
);

AND2x4_ASAP7_75t_L g2014 ( 
.A(n_1944),
.B(n_1928),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1952),
.B(n_1899),
.Y(n_2015)
);

HB1xp67_ASAP7_75t_L g2016 ( 
.A(n_1946),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1968),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1953),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1971),
.B(n_1935),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1968),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1950),
.B(n_1935),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1953),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1978),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1978),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1979),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1955),
.B(n_1902),
.Y(n_2026)
);

OR2x2_ASAP7_75t_L g2027 ( 
.A(n_1948),
.B(n_1903),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1950),
.B(n_1936),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1979),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1969),
.B(n_1936),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1988),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1988),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1975),
.Y(n_2033)
);

AOI21xp5_ASAP7_75t_L g2034 ( 
.A1(n_1960),
.A2(n_1928),
.B(n_1925),
.Y(n_2034)
);

BUFx2_ASAP7_75t_L g2035 ( 
.A(n_1960),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1969),
.B(n_1923),
.Y(n_2036)
);

INVxp67_ASAP7_75t_L g2037 ( 
.A(n_1944),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1944),
.B(n_1923),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1960),
.B(n_1915),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_2013),
.B(n_1967),
.Y(n_2040)
);

OAI21xp33_ASAP7_75t_L g2041 ( 
.A1(n_1998),
.A2(n_1916),
.B(n_1941),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1994),
.B(n_1954),
.Y(n_2042)
);

INVxp67_ASAP7_75t_SL g2043 ( 
.A(n_2006),
.Y(n_2043)
);

OR2x2_ASAP7_75t_L g2044 ( 
.A(n_1990),
.B(n_2016),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_2007),
.B(n_1967),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_SL g2046 ( 
.A(n_2034),
.B(n_1900),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1994),
.B(n_1954),
.Y(n_2047)
);

OR2x2_ASAP7_75t_L g2048 ( 
.A(n_1990),
.B(n_1970),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_2019),
.B(n_1987),
.Y(n_2049)
);

OR2x2_ASAP7_75t_L g2050 ( 
.A(n_2027),
.B(n_1970),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1999),
.Y(n_2051)
);

OR2x2_ASAP7_75t_L g2052 ( 
.A(n_2027),
.B(n_1980),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1999),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_2037),
.B(n_1985),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1997),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1992),
.B(n_1985),
.Y(n_2056)
);

NAND2x1p5_ASAP7_75t_L g2057 ( 
.A(n_2014),
.B(n_1976),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_2021),
.B(n_1986),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_2026),
.B(n_1955),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_2026),
.B(n_1956),
.Y(n_2060)
);

INVx2_ASAP7_75t_SL g2061 ( 
.A(n_2009),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_2009),
.B(n_1956),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_2028),
.B(n_1986),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_2005),
.B(n_1947),
.Y(n_2064)
);

OR2x2_ASAP7_75t_L g2065 ( 
.A(n_2030),
.B(n_1980),
.Y(n_2065)
);

INVxp67_ASAP7_75t_L g2066 ( 
.A(n_2014),
.Y(n_2066)
);

OR2x6_ASAP7_75t_L g2067 ( 
.A(n_2005),
.B(n_1914),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_2005),
.B(n_1947),
.Y(n_2068)
);

OR2x2_ASAP7_75t_L g2069 ( 
.A(n_1995),
.B(n_1962),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1989),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1997),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2000),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1989),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2000),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_2014),
.B(n_1914),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_2005),
.B(n_1949),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_2015),
.B(n_2001),
.Y(n_2077)
);

AOI22xp5_ASAP7_75t_L g2078 ( 
.A1(n_2035),
.A2(n_1945),
.B1(n_1941),
.B2(n_1823),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2002),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_2077),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_2077),
.B(n_1995),
.Y(n_2081)
);

AOI22xp5_ASAP7_75t_L g2082 ( 
.A1(n_2041),
.A2(n_1945),
.B1(n_2035),
.B2(n_2039),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2055),
.Y(n_2083)
);

AOI22xp5_ASAP7_75t_L g2084 ( 
.A1(n_2041),
.A2(n_2003),
.B1(n_1917),
.B2(n_2001),
.Y(n_2084)
);

AOI211xp5_ASAP7_75t_L g2085 ( 
.A1(n_2046),
.A2(n_1778),
.B(n_2038),
.C(n_2033),
.Y(n_2085)
);

OAI21xp33_ASAP7_75t_SL g2086 ( 
.A1(n_2040),
.A2(n_2015),
.B(n_2036),
.Y(n_2086)
);

NOR2xp33_ASAP7_75t_L g2087 ( 
.A(n_2066),
.B(n_1914),
.Y(n_2087)
);

NAND2xp33_ASAP7_75t_L g2088 ( 
.A(n_2044),
.B(n_2004),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_2043),
.B(n_1914),
.Y(n_2089)
);

INVx1_ASAP7_75t_SL g2090 ( 
.A(n_2044),
.Y(n_2090)
);

OAI221xp5_ASAP7_75t_L g2091 ( 
.A1(n_2078),
.A2(n_2003),
.B1(n_2004),
.B2(n_1933),
.C(n_1903),
.Y(n_2091)
);

AOI21xp5_ASAP7_75t_L g2092 ( 
.A1(n_2078),
.A2(n_2004),
.B(n_1984),
.Y(n_2092)
);

AOI21xp33_ASAP7_75t_L g2093 ( 
.A1(n_2067),
.A2(n_1917),
.B(n_2002),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2055),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2071),
.Y(n_2095)
);

NOR2x1_ASAP7_75t_L g2096 ( 
.A(n_2067),
.B(n_1845),
.Y(n_2096)
);

AOI22xp5_ASAP7_75t_L g2097 ( 
.A1(n_2061),
.A2(n_1917),
.B1(n_1919),
.B2(n_1911),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2071),
.Y(n_2098)
);

NOR2xp33_ASAP7_75t_L g2099 ( 
.A(n_2049),
.B(n_2045),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2061),
.B(n_1991),
.Y(n_2100)
);

INVxp67_ASAP7_75t_SL g2101 ( 
.A(n_2057),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2072),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_2042),
.B(n_1993),
.Y(n_2103)
);

OAI22xp33_ASAP7_75t_L g2104 ( 
.A1(n_2067),
.A2(n_1951),
.B1(n_1926),
.B2(n_1844),
.Y(n_2104)
);

AOI21xp5_ASAP7_75t_SL g2105 ( 
.A1(n_2067),
.A2(n_1779),
.B(n_1951),
.Y(n_2105)
);

AOI221x1_ASAP7_75t_L g2106 ( 
.A1(n_2075),
.A2(n_1975),
.B1(n_2031),
.B2(n_2029),
.C(n_2008),
.Y(n_2106)
);

OAI22xp5_ASAP7_75t_L g2107 ( 
.A1(n_2057),
.A2(n_1926),
.B1(n_1911),
.B2(n_1932),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_SL g2108 ( 
.A(n_2042),
.B(n_1932),
.Y(n_2108)
);

OAI22xp33_ASAP7_75t_L g2109 ( 
.A1(n_2067),
.A2(n_1836),
.B1(n_1794),
.B2(n_1915),
.Y(n_2109)
);

INVx2_ASAP7_75t_SL g2110 ( 
.A(n_2081),
.Y(n_2110)
);

AOI22xp33_ASAP7_75t_SL g2111 ( 
.A1(n_2090),
.A2(n_2057),
.B1(n_2047),
.B2(n_2053),
.Y(n_2111)
);

AOI22xp5_ASAP7_75t_L g2112 ( 
.A1(n_2082),
.A2(n_2064),
.B1(n_2076),
.B2(n_2068),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_2099),
.B(n_2047),
.Y(n_2113)
);

AOI21xp5_ASAP7_75t_L g2114 ( 
.A1(n_2105),
.A2(n_2056),
.B(n_2072),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2083),
.Y(n_2115)
);

OAI21xp33_ASAP7_75t_L g2116 ( 
.A1(n_2096),
.A2(n_2054),
.B(n_2064),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_2080),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2094),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_2087),
.B(n_2051),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2095),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2098),
.Y(n_2121)
);

INVxp67_ASAP7_75t_SL g2122 ( 
.A(n_2101),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2102),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_2099),
.B(n_2051),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_2087),
.B(n_2051),
.Y(n_2125)
);

OAI22xp5_ASAP7_75t_L g2126 ( 
.A1(n_2084),
.A2(n_2053),
.B1(n_2063),
.B2(n_2058),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2089),
.B(n_2053),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2100),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2103),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2106),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2108),
.Y(n_2131)
);

AOI21xp33_ASAP7_75t_L g2132 ( 
.A1(n_2088),
.A2(n_2076),
.B(n_2068),
.Y(n_2132)
);

AND2x4_ASAP7_75t_L g2133 ( 
.A(n_2092),
.B(n_2062),
.Y(n_2133)
);

NOR4xp25_ASAP7_75t_SL g2134 ( 
.A(n_2091),
.B(n_2079),
.C(n_2074),
.D(n_2008),
.Y(n_2134)
);

HB1xp67_ASAP7_75t_L g2135 ( 
.A(n_2122),
.Y(n_2135)
);

INVxp67_ASAP7_75t_L g2136 ( 
.A(n_2122),
.Y(n_2136)
);

OAI22xp33_ASAP7_75t_SL g2137 ( 
.A1(n_2130),
.A2(n_2097),
.B1(n_2107),
.B2(n_2069),
.Y(n_2137)
);

NAND2xp33_ASAP7_75t_SL g2138 ( 
.A(n_2134),
.B(n_1974),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_2110),
.Y(n_2139)
);

OAI321xp33_ASAP7_75t_L g2140 ( 
.A1(n_2126),
.A2(n_2104),
.A3(n_2109),
.B1(n_2085),
.B2(n_2069),
.C(n_2052),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2133),
.B(n_2062),
.Y(n_2141)
);

NAND3xp33_ASAP7_75t_L g2142 ( 
.A(n_2111),
.B(n_2086),
.C(n_2093),
.Y(n_2142)
);

NOR2x1_ASAP7_75t_L g2143 ( 
.A(n_2114),
.B(n_2104),
.Y(n_2143)
);

INVx1_ASAP7_75t_SL g2144 ( 
.A(n_2133),
.Y(n_2144)
);

O2A1O1Ixp33_ASAP7_75t_L g2145 ( 
.A1(n_2114),
.A2(n_2109),
.B(n_2079),
.C(n_2074),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2117),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2117),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2115),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_SL g2149 ( 
.A(n_2111),
.B(n_2048),
.Y(n_2149)
);

NAND3xp33_ASAP7_75t_L g2150 ( 
.A(n_2143),
.B(n_2112),
.C(n_2132),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2135),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_SL g2152 ( 
.A(n_2140),
.B(n_2113),
.Y(n_2152)
);

NOR2xp67_ASAP7_75t_L g2153 ( 
.A(n_2136),
.B(n_2131),
.Y(n_2153)
);

NOR2x1_ASAP7_75t_L g2154 ( 
.A(n_2149),
.B(n_2118),
.Y(n_2154)
);

OAI21xp5_ASAP7_75t_L g2155 ( 
.A1(n_2142),
.A2(n_2116),
.B(n_2124),
.Y(n_2155)
);

CKINVDCx20_ASAP7_75t_R g2156 ( 
.A(n_2144),
.Y(n_2156)
);

INVxp67_ASAP7_75t_L g2157 ( 
.A(n_2149),
.Y(n_2157)
);

NAND4xp25_ASAP7_75t_L g2158 ( 
.A(n_2141),
.B(n_2129),
.C(n_2125),
.D(n_2127),
.Y(n_2158)
);

NAND4xp25_ASAP7_75t_SL g2159 ( 
.A(n_2145),
.B(n_2119),
.C(n_2128),
.D(n_2121),
.Y(n_2159)
);

O2A1O1Ixp5_ASAP7_75t_L g2160 ( 
.A1(n_2138),
.A2(n_2123),
.B(n_2120),
.C(n_2073),
.Y(n_2160)
);

OAI21xp5_ASAP7_75t_L g2161 ( 
.A1(n_2157),
.A2(n_2138),
.B(n_2137),
.Y(n_2161)
);

OAI221xp5_ASAP7_75t_L g2162 ( 
.A1(n_2154),
.A2(n_2139),
.B1(n_2147),
.B2(n_2146),
.C(n_2148),
.Y(n_2162)
);

O2A1O1Ixp33_ASAP7_75t_L g2163 ( 
.A1(n_2152),
.A2(n_2139),
.B(n_2048),
.C(n_2052),
.Y(n_2163)
);

CKINVDCx16_ASAP7_75t_R g2164 ( 
.A(n_2156),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2153),
.B(n_2059),
.Y(n_2165)
);

AOI222xp33_ASAP7_75t_L g2166 ( 
.A1(n_2155),
.A2(n_2073),
.B1(n_2070),
.B2(n_2060),
.C1(n_2059),
.C2(n_2029),
.Y(n_2166)
);

AOI221xp5_ASAP7_75t_L g2167 ( 
.A1(n_2150),
.A2(n_2073),
.B1(n_2070),
.B2(n_2050),
.C(n_2060),
.Y(n_2167)
);

INVx1_ASAP7_75t_SL g2168 ( 
.A(n_2164),
.Y(n_2168)
);

NAND3xp33_ASAP7_75t_SL g2169 ( 
.A(n_2161),
.B(n_2160),
.C(n_2151),
.Y(n_2169)
);

O2A1O1Ixp33_ASAP7_75t_L g2170 ( 
.A1(n_2162),
.A2(n_2158),
.B(n_2159),
.C(n_2050),
.Y(n_2170)
);

OAI21xp33_ASAP7_75t_L g2171 ( 
.A1(n_2165),
.A2(n_2070),
.B(n_2065),
.Y(n_2171)
);

AO22x2_ASAP7_75t_L g2172 ( 
.A1(n_2163),
.A2(n_2031),
.B1(n_2032),
.B2(n_2017),
.Y(n_2172)
);

O2A1O1Ixp33_ASAP7_75t_L g2173 ( 
.A1(n_2167),
.A2(n_2065),
.B(n_1819),
.C(n_2032),
.Y(n_2173)
);

INVx1_ASAP7_75t_SL g2174 ( 
.A(n_2166),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2168),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_2174),
.B(n_1996),
.Y(n_2176)
);

AND2x4_ASAP7_75t_L g2177 ( 
.A(n_2169),
.B(n_2025),
.Y(n_2177)
);

OAI22xp5_ASAP7_75t_L g2178 ( 
.A1(n_2170),
.A2(n_2024),
.B1(n_2023),
.B2(n_2010),
.Y(n_2178)
);

AND2x4_ASAP7_75t_L g2179 ( 
.A(n_2172),
.B(n_2011),
.Y(n_2179)
);

OAI221xp5_ASAP7_75t_L g2180 ( 
.A1(n_2175),
.A2(n_2171),
.B1(n_2173),
.B2(n_2012),
.C(n_2020),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_2177),
.B(n_2018),
.Y(n_2181)
);

AND2x4_ASAP7_75t_L g2182 ( 
.A(n_2179),
.B(n_2018),
.Y(n_2182)
);

XNOR2xp5_ASAP7_75t_L g2183 ( 
.A(n_2180),
.B(n_2178),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2183),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2184),
.B(n_2176),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2184),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2185),
.Y(n_2187)
);

BUFx2_ASAP7_75t_L g2188 ( 
.A(n_2186),
.Y(n_2188)
);

AOI22xp5_ASAP7_75t_L g2189 ( 
.A1(n_2188),
.A2(n_2181),
.B1(n_2182),
.B2(n_2022),
.Y(n_2189)
);

AOI22xp5_ASAP7_75t_L g2190 ( 
.A1(n_2187),
.A2(n_2022),
.B1(n_1964),
.B2(n_1942),
.Y(n_2190)
);

OAI21xp5_ASAP7_75t_SL g2191 ( 
.A1(n_2189),
.A2(n_1911),
.B(n_1921),
.Y(n_2191)
);

AOI21xp5_ASAP7_75t_L g2192 ( 
.A1(n_2191),
.A2(n_2190),
.B(n_1983),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2192),
.Y(n_2193)
);

OAI221xp5_ASAP7_75t_R g2194 ( 
.A1(n_2193),
.A2(n_1974),
.B1(n_1977),
.B2(n_1898),
.C(n_1982),
.Y(n_2194)
);

AOI211xp5_ASAP7_75t_L g2195 ( 
.A1(n_2194),
.A2(n_1983),
.B(n_1982),
.C(n_1771),
.Y(n_2195)
);


endmodule