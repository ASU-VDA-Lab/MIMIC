module fake_jpeg_26191_n_168 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_168);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_34),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_33),
.Y(n_39)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_22),
.Y(n_49)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_37),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_36),
.B(n_18),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_14),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_20),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_37),
.B(n_22),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_50),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_14),
.Y(n_58)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_26),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_57),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_23),
.B1(n_46),
.B2(n_32),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_69),
.B1(n_31),
.B2(n_39),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_23),
.B1(n_18),
.B2(n_25),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_54),
.Y(n_93)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

OAI21xp33_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_23),
.B(n_16),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_21),
.B(n_19),
.C(n_27),
.Y(n_80)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_58),
.B(n_16),
.Y(n_75)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_61),
.Y(n_86)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_33),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_66),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_26),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_65),
.B(n_68),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_33),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_48),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_47),
.A2(n_32),
.B1(n_30),
.B2(n_34),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_40),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_70),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_50),
.B(n_25),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_21),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_39),
.A2(n_27),
.B(n_3),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_2),
.B(n_3),
.Y(n_84)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_75),
.B(n_85),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_34),
.B1(n_31),
.B2(n_27),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_84),
.B1(n_72),
.B2(n_93),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_55),
.B1(n_67),
.B2(n_70),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_92),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_33),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_81),
.Y(n_104)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_90),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_28),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_59),
.B(n_64),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_89),
.Y(n_102)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_27),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_66),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_33),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_61),
.C(n_66),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_89),
.C(n_90),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_107),
.B1(n_77),
.B2(n_91),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_111),
.B1(n_80),
.B2(n_83),
.Y(n_126)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_105),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_77),
.Y(n_101)
);

NOR3xp33_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_108),
.C(n_86),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_60),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_106),
.B(n_86),
.Y(n_127)
);

OAI22x1_ASAP7_75t_L g107 ( 
.A1(n_93),
.A2(n_19),
.B1(n_69),
.B2(n_39),
.Y(n_107)
);

NOR3xp33_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_76),
.C(n_60),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_110),
.Y(n_122)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_87),
.A2(n_68),
.B1(n_71),
.B2(n_62),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_87),
.B(n_92),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_125),
.Y(n_133)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

AO21x1_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_92),
.B(n_81),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_117),
.Y(n_129)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_118),
.A2(n_124),
.B1(n_48),
.B2(n_40),
.Y(n_139)
);

NAND3xp33_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_127),
.C(n_58),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_126),
.C(n_102),
.Y(n_131)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

INVxp33_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_98),
.A2(n_87),
.B(n_81),
.Y(n_125)
);

A2O1A1O1Ixp25_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_104),
.B(n_102),
.C(n_94),
.D(n_111),
.Y(n_130)
);

AOI321xp33_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_62),
.A3(n_21),
.B1(n_19),
.B2(n_28),
.C(n_13),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_21),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_104),
.C(n_96),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_137),
.C(n_133),
.Y(n_149)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_122),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_96),
.C(n_103),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_139),
.A2(n_117),
.B1(n_122),
.B2(n_121),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_73),
.Y(n_146)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_142),
.A2(n_144),
.B(n_146),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_133),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_148),
.C(n_149),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_126),
.B1(n_116),
.B2(n_123),
.Y(n_144)
);

AOI322xp5_ASAP7_75t_L g145 ( 
.A1(n_130),
.A2(n_115),
.A3(n_116),
.B1(n_73),
.B2(n_79),
.C1(n_75),
.C2(n_58),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_145),
.A2(n_137),
.B(n_135),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_147),
.A2(n_129),
.B(n_128),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_148),
.B(n_134),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_151),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_SL g160 ( 
.A1(n_153),
.A2(n_132),
.B(n_136),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_149),
.A2(n_129),
.B(n_134),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_156),
.A2(n_147),
.B(n_143),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_SL g164 ( 
.A1(n_157),
.A2(n_159),
.B(n_160),
.C(n_161),
.Y(n_164)
);

OAI31xp33_ASAP7_75t_L g159 ( 
.A1(n_155),
.A2(n_152),
.A3(n_132),
.B(n_154),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_154),
.A2(n_138),
.B(n_9),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_L g162 ( 
.A1(n_158),
.A2(n_10),
.A3(n_40),
.B1(n_48),
.B2(n_7),
.C1(n_2),
.C2(n_5),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_162),
.B(n_8),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_160),
.A2(n_40),
.B1(n_5),
.B2(n_7),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_163),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_166),
.B(n_164),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_165),
.Y(n_168)
);


endmodule