module fake_jpeg_3197_n_62 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_62);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_62;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_18),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_6),
.B(n_13),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_20),
.B(n_2),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_20),
.Y(n_29)
);

NAND2xp33_ASAP7_75t_SL g27 ( 
.A(n_19),
.B(n_3),
.Y(n_27)
);

NAND3xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_20),
.C(n_19),
.Y(n_33)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_26),
.B(n_22),
.Y(n_30)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_3),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_31),
.A2(n_25),
.B1(n_28),
.B2(n_19),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_38),
.B1(n_34),
.B2(n_24),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_31),
.A2(n_25),
.B1(n_21),
.B2(n_24),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_SL g40 ( 
.A(n_32),
.B(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_39),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_21),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_42),
.B(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_34),
.C(n_24),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_46),
.A2(n_4),
.B1(n_5),
.B2(n_24),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_51),
.Y(n_52)
);

INVxp33_ASAP7_75t_SL g54 ( 
.A(n_50),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_4),
.B(n_5),
.C(n_7),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_41),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_55),
.B(n_52),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_48),
.A2(n_8),
.B1(n_10),
.B2(n_12),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_57),
.Y(n_58)
);

BUFx24_ASAP7_75t_SL g57 ( 
.A(n_55),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_54),
.C(n_49),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_15),
.C(n_16),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_61),
.B(n_17),
.Y(n_62)
);


endmodule