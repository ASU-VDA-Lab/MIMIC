module fake_aes_10648_n_673 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_673);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_673;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_73), .Y(n_90) );
BUFx8_ASAP7_75t_SL g91 ( .A(n_35), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_81), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_88), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_75), .Y(n_94) );
CKINVDCx20_ASAP7_75t_R g95 ( .A(n_61), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_22), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_68), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_3), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_6), .Y(n_99) );
INVx1_ASAP7_75t_SL g100 ( .A(n_79), .Y(n_100) );
INVxp67_ASAP7_75t_L g101 ( .A(n_16), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_8), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_13), .Y(n_103) );
INVxp67_ASAP7_75t_L g104 ( .A(n_43), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_34), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_27), .Y(n_106) );
HB1xp67_ASAP7_75t_L g107 ( .A(n_52), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_8), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_26), .Y(n_109) );
BUFx2_ASAP7_75t_L g110 ( .A(n_71), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_3), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_47), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_49), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_44), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_22), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_69), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_23), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_11), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_28), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_4), .Y(n_120) );
INVxp33_ASAP7_75t_L g121 ( .A(n_57), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_20), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_1), .Y(n_123) );
INVxp67_ASAP7_75t_SL g124 ( .A(n_6), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_0), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_37), .Y(n_126) );
INVxp67_ASAP7_75t_L g127 ( .A(n_18), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_83), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_0), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_77), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_99), .Y(n_131) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_92), .A2(n_41), .B(n_87), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_110), .B(n_1), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_110), .B(n_2), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_106), .Y(n_135) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_92), .A2(n_42), .B(n_86), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_99), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_106), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_107), .B(n_2), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_99), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_106), .Y(n_141) );
AND2x2_ASAP7_75t_L g142 ( .A(n_107), .B(n_4), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_112), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_119), .B(n_5), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g145 ( .A(n_119), .B(n_5), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_93), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_98), .B(n_7), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_98), .B(n_7), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_93), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_94), .Y(n_150) );
CKINVDCx8_ASAP7_75t_R g151 ( .A(n_116), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_112), .B(n_9), .Y(n_152) );
NOR2x1_ASAP7_75t_L g153 ( .A(n_94), .B(n_9), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_97), .Y(n_154) );
AND2x4_ASAP7_75t_L g155 ( .A(n_112), .B(n_10), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_97), .Y(n_156) );
OAI22xp5_ASAP7_75t_SL g157 ( .A1(n_108), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_157) );
OAI22xp5_ASAP7_75t_SL g158 ( .A1(n_124), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_138), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_135), .Y(n_160) );
INVx4_ASAP7_75t_L g161 ( .A(n_144), .Y(n_161) );
AND3x2_ASAP7_75t_L g162 ( .A(n_134), .B(n_124), .C(n_113), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_146), .B(n_104), .Y(n_163) );
OR2x2_ASAP7_75t_L g164 ( .A(n_134), .B(n_101), .Y(n_164) );
INVx2_ASAP7_75t_SL g165 ( .A(n_146), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_149), .B(n_104), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_138), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_134), .B(n_121), .Y(n_168) );
INVxp67_ASAP7_75t_SL g169 ( .A(n_139), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_138), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_152), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_142), .B(n_102), .Y(n_172) );
AND2x6_ASAP7_75t_L g173 ( .A(n_152), .B(n_105), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_149), .B(n_105), .Y(n_174) );
BUFx2_ASAP7_75t_L g175 ( .A(n_133), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_133), .A2(n_90), .B1(n_128), .B2(n_95), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_138), .Y(n_177) );
OR2x2_ASAP7_75t_L g178 ( .A(n_142), .B(n_101), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_150), .B(n_114), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_150), .B(n_114), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_133), .B(n_126), .Y(n_181) );
INVx2_ASAP7_75t_SL g182 ( .A(n_154), .Y(n_182) );
BUFx3_ASAP7_75t_L g183 ( .A(n_152), .Y(n_183) );
XNOR2xp5_ASAP7_75t_L g184 ( .A(n_157), .B(n_96), .Y(n_184) );
OR2x6_ASAP7_75t_L g185 ( .A(n_133), .B(n_102), .Y(n_185) );
BUFx3_ASAP7_75t_L g186 ( .A(n_152), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_151), .Y(n_187) );
AND2x6_ASAP7_75t_L g188 ( .A(n_152), .B(n_126), .Y(n_188) );
AO22x2_ASAP7_75t_L g189 ( .A1(n_144), .A2(n_113), .B1(n_130), .B2(n_126), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_154), .B(n_130), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_138), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g192 ( .A1(n_155), .A2(n_118), .B1(n_129), .B2(n_103), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_138), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_169), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_169), .Y(n_195) );
NOR3x1_ASAP7_75t_L g196 ( .A(n_164), .B(n_157), .C(n_139), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_189), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_185), .B(n_133), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_178), .B(n_151), .Y(n_199) );
OR2x6_ASAP7_75t_L g200 ( .A(n_185), .B(n_158), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_168), .B(n_142), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_185), .A2(n_144), .B1(n_155), .B2(n_147), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_189), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_160), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_189), .Y(n_205) );
INVx2_ASAP7_75t_SL g206 ( .A(n_161), .Y(n_206) );
INVxp67_ASAP7_75t_SL g207 ( .A(n_165), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g208 ( .A1(n_189), .A2(n_144), .B1(n_155), .B2(n_145), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_183), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_168), .B(n_144), .Y(n_210) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_189), .A2(n_155), .B1(n_145), .B2(n_156), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_161), .B(n_155), .Y(n_212) );
NOR2x2_ASAP7_75t_L g213 ( .A(n_185), .B(n_158), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_189), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_160), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_178), .B(n_151), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_161), .B(n_156), .Y(n_217) );
INVx2_ASAP7_75t_SL g218 ( .A(n_161), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_168), .B(n_147), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_163), .B(n_148), .Y(n_220) );
AND2x6_ASAP7_75t_L g221 ( .A(n_183), .B(n_153), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_178), .B(n_148), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g223 ( .A1(n_185), .A2(n_109), .B1(n_123), .B2(n_127), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_161), .Y(n_224) );
INVxp67_ASAP7_75t_L g225 ( .A(n_164), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_164), .B(n_127), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_188), .A2(n_153), .B1(n_129), .B2(n_125), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_163), .B(n_131), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_171), .A2(n_143), .B(n_141), .C(n_135), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_183), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_185), .A2(n_125), .B1(n_122), .B2(n_103), .Y(n_231) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_173), .A2(n_118), .B1(n_120), .B2(n_122), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_186), .Y(n_233) );
NAND2xp33_ASAP7_75t_L g234 ( .A(n_173), .B(n_138), .Y(n_234) );
INVxp67_ASAP7_75t_L g235 ( .A(n_166), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_166), .B(n_131), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_188), .A2(n_115), .B1(n_117), .B2(n_120), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_186), .Y(n_238) );
AND2x2_ASAP7_75t_SL g239 ( .A(n_175), .B(n_132), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_SL g240 ( .A1(n_199), .A2(n_180), .B(n_179), .C(n_174), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_216), .B(n_172), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_194), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_235), .B(n_172), .Y(n_243) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_222), .A2(n_171), .B(n_175), .C(n_186), .Y(n_244) );
NOR3xp33_ASAP7_75t_SL g245 ( .A(n_219), .B(n_187), .C(n_184), .Y(n_245) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_202), .A2(n_171), .B(n_174), .C(n_179), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_207), .A2(n_181), .B(n_165), .Y(n_247) );
NAND2x2_ASAP7_75t_L g248 ( .A(n_196), .B(n_184), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_217), .A2(n_165), .B(n_182), .Y(n_249) );
NAND2xp33_ASAP7_75t_R g250 ( .A(n_198), .B(n_162), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g251 ( .A(n_223), .Y(n_251) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_198), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_L g253 ( .A1(n_225), .A2(n_171), .B(n_172), .C(n_182), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_195), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_L g255 ( .A1(n_210), .A2(n_171), .B(n_182), .C(n_190), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_L g256 ( .A1(n_197), .A2(n_203), .B(n_205), .C(n_214), .Y(n_256) );
INVx3_ASAP7_75t_L g257 ( .A(n_209), .Y(n_257) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_229), .A2(n_180), .B(n_192), .C(n_190), .Y(n_258) );
INVx3_ASAP7_75t_L g259 ( .A(n_209), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_217), .A2(n_192), .B(n_132), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_201), .B(n_162), .Y(n_261) );
AOI33xp33_ASAP7_75t_L g262 ( .A1(n_226), .A2(n_140), .A3(n_137), .B1(n_111), .B2(n_115), .B3(n_117), .Y(n_262) );
AND2x4_ASAP7_75t_L g263 ( .A(n_198), .B(n_173), .Y(n_263) );
INVx3_ASAP7_75t_L g264 ( .A(n_209), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_212), .A2(n_132), .B(n_136), .Y(n_265) );
NAND2x1p5_ASAP7_75t_L g266 ( .A(n_224), .B(n_111), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_206), .B(n_138), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_L g268 ( .A1(n_229), .A2(n_143), .B(n_135), .C(n_141), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_220), .B(n_173), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_208), .A2(n_176), .B1(n_173), .B2(n_188), .Y(n_270) );
NAND2x1p5_ASAP7_75t_L g271 ( .A(n_224), .B(n_137), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_201), .B(n_176), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_211), .B(n_173), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_200), .B(n_173), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_231), .B(n_173), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_209), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_204), .Y(n_277) );
OAI22xp5_ASAP7_75t_L g278 ( .A1(n_232), .A2(n_173), .B1(n_188), .B2(n_100), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_206), .B(n_130), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_228), .B(n_188), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_212), .A2(n_136), .B(n_132), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_204), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_224), .Y(n_283) );
OAI22xp5_ASAP7_75t_L g284 ( .A1(n_215), .A2(n_188), .B1(n_100), .B2(n_143), .Y(n_284) );
A2O1A1Ixp33_ASAP7_75t_L g285 ( .A1(n_241), .A2(n_238), .B(n_230), .C(n_233), .Y(n_285) );
A2O1A1Ixp33_ASAP7_75t_L g286 ( .A1(n_241), .A2(n_227), .B(n_236), .C(n_237), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_243), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_242), .Y(n_288) );
O2A1O1Ixp33_ASAP7_75t_L g289 ( .A1(n_240), .A2(n_200), .B(n_234), .C(n_140), .Y(n_289) );
AO31x2_ASAP7_75t_L g290 ( .A1(n_265), .A2(n_143), .A3(n_135), .B(n_141), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_272), .B(n_200), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_272), .B(n_221), .Y(n_292) );
A2O1A1Ixp33_ASAP7_75t_L g293 ( .A1(n_255), .A2(n_239), .B(n_234), .C(n_218), .Y(n_293) );
A2O1A1Ixp33_ASAP7_75t_L g294 ( .A1(n_246), .A2(n_239), .B(n_218), .C(n_141), .Y(n_294) );
AOI221x1_ASAP7_75t_L g295 ( .A1(n_281), .A2(n_177), .B1(n_159), .B2(n_193), .C(n_191), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_267), .A2(n_132), .B(n_136), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_270), .A2(n_200), .B1(n_221), .B2(n_188), .Y(n_297) );
A2O1A1Ixp33_ASAP7_75t_L g298 ( .A1(n_253), .A2(n_221), .B(n_177), .C(n_193), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_251), .A2(n_221), .B1(n_188), .B2(n_213), .Y(n_299) );
INVxp67_ASAP7_75t_L g300 ( .A(n_250), .Y(n_300) );
OAI21xp5_ASAP7_75t_L g301 ( .A1(n_260), .A2(n_221), .B(n_188), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_261), .B(n_221), .Y(n_302) );
AO31x2_ASAP7_75t_L g303 ( .A1(n_258), .A2(n_170), .A3(n_193), .B(n_191), .Y(n_303) );
AOI22xp33_ASAP7_75t_SL g304 ( .A1(n_248), .A2(n_213), .B1(n_136), .B2(n_91), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_254), .Y(n_305) );
O2A1O1Ixp33_ASAP7_75t_SL g306 ( .A1(n_240), .A2(n_191), .B(n_177), .C(n_170), .Y(n_306) );
O2A1O1Ixp33_ASAP7_75t_L g307 ( .A1(n_244), .A2(n_170), .B(n_167), .C(n_159), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_261), .B(n_14), .Y(n_308) );
BUFx2_ASAP7_75t_L g309 ( .A(n_263), .Y(n_309) );
O2A1O1Ixp33_ASAP7_75t_L g310 ( .A1(n_269), .A2(n_167), .B(n_159), .C(n_136), .Y(n_310) );
OAI21xp5_ASAP7_75t_L g311 ( .A1(n_280), .A2(n_167), .B(n_51), .Y(n_311) );
AOI221xp5_ASAP7_75t_L g312 ( .A1(n_245), .A2(n_15), .B1(n_16), .B2(n_17), .C(n_18), .Y(n_312) );
CKINVDCx20_ASAP7_75t_R g313 ( .A(n_245), .Y(n_313) );
O2A1O1Ixp33_ASAP7_75t_L g314 ( .A1(n_273), .A2(n_15), .B(n_17), .C(n_19), .Y(n_314) );
A2O1A1Ixp33_ASAP7_75t_L g315 ( .A1(n_268), .A2(n_19), .B(n_20), .C(n_21), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_266), .Y(n_316) );
NAND2x1p5_ASAP7_75t_L g317 ( .A(n_263), .B(n_21), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_274), .B(n_23), .Y(n_318) );
AO32x2_ASAP7_75t_L g319 ( .A1(n_284), .A2(n_24), .A3(n_25), .B1(n_26), .B2(n_29), .Y(n_319) );
OAI21xp33_ASAP7_75t_SL g320 ( .A1(n_262), .A2(n_24), .B(n_25), .Y(n_320) );
OAI21xp5_ASAP7_75t_L g321 ( .A1(n_249), .A2(n_30), .B(n_31), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_287), .B(n_256), .Y(n_322) );
OA21x2_ASAP7_75t_L g323 ( .A1(n_295), .A2(n_279), .B(n_267), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_291), .A2(n_248), .B1(n_278), .B2(n_252), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_297), .A2(n_266), .B1(n_275), .B2(n_277), .Y(n_325) );
A2O1A1Ixp33_ASAP7_75t_L g326 ( .A1(n_320), .A2(n_247), .B(n_282), .C(n_283), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_288), .B(n_252), .Y(n_327) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_306), .A2(n_279), .B(n_276), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_292), .B(n_252), .Y(n_329) );
O2A1O1Ixp33_ASAP7_75t_L g330 ( .A1(n_286), .A2(n_271), .B(n_276), .C(n_264), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_310), .A2(n_264), .B(n_259), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_305), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_299), .B(n_252), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_301), .A2(n_259), .B(n_257), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_302), .B(n_271), .Y(n_335) );
INVxp67_ASAP7_75t_L g336 ( .A(n_318), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_301), .A2(n_257), .B(n_250), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_317), .Y(n_338) );
AOI21xp5_ASAP7_75t_L g339 ( .A1(n_294), .A2(n_32), .B(n_33), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_317), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_290), .Y(n_341) );
AOI222xp33_ASAP7_75t_L g342 ( .A1(n_300), .A2(n_36), .B1(n_38), .B2(n_39), .C1(n_40), .C2(n_45), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_290), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_290), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_303), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_303), .Y(n_346) );
INVx4_ASAP7_75t_SL g347 ( .A(n_318), .Y(n_347) );
O2A1O1Ixp33_ASAP7_75t_L g348 ( .A1(n_315), .A2(n_46), .B(n_48), .C(n_50), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_303), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_316), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_309), .B(n_53), .Y(n_351) );
OAI21x1_ASAP7_75t_L g352 ( .A1(n_345), .A2(n_311), .B(n_321), .Y(n_352) );
INVx3_ASAP7_75t_L g353 ( .A(n_343), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_347), .B(n_319), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_338), .A2(n_304), .B1(n_308), .B2(n_285), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_341), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_341), .B(n_298), .Y(n_357) );
OAI21xp5_ASAP7_75t_L g358 ( .A1(n_326), .A2(n_289), .B(n_293), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_343), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_347), .B(n_319), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_332), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_332), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_344), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_344), .Y(n_364) );
OAI21xp33_ASAP7_75t_L g365 ( .A1(n_342), .A2(n_312), .B(n_314), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_345), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_346), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_346), .Y(n_368) );
INVx1_ASAP7_75t_SL g369 ( .A(n_347), .Y(n_369) );
INVx5_ASAP7_75t_L g370 ( .A(n_347), .Y(n_370) );
INVx3_ASAP7_75t_L g371 ( .A(n_338), .Y(n_371) );
OA21x2_ASAP7_75t_L g372 ( .A1(n_349), .A2(n_296), .B(n_321), .Y(n_372) );
AOI221xp5_ASAP7_75t_L g373 ( .A1(n_324), .A2(n_313), .B1(n_307), .B2(n_319), .C(n_58), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_322), .B(n_54), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_349), .Y(n_375) );
OR2x6_ASAP7_75t_L g376 ( .A(n_337), .B(n_55), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_329), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_322), .B(n_56), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_323), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_323), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_359), .B(n_364), .Y(n_381) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_353), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_356), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_359), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_359), .B(n_340), .Y(n_385) );
INVx1_ASAP7_75t_SL g386 ( .A(n_371), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_359), .Y(n_387) );
BUFx2_ASAP7_75t_L g388 ( .A(n_353), .Y(n_388) );
AOI222xp33_ASAP7_75t_L g389 ( .A1(n_355), .A2(n_336), .B1(n_340), .B2(n_325), .C1(n_351), .C2(n_329), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_363), .B(n_350), .Y(n_390) );
OA21x2_ASAP7_75t_L g391 ( .A1(n_358), .A2(n_331), .B(n_328), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_356), .Y(n_392) );
INVxp67_ASAP7_75t_L g393 ( .A(n_354), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_363), .B(n_350), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_366), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_366), .Y(n_396) );
BUFx2_ASAP7_75t_L g397 ( .A(n_353), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_363), .B(n_323), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_368), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_368), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_363), .B(n_323), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_375), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_353), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_375), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_355), .A2(n_342), .B1(n_325), .B2(n_333), .Y(n_405) );
BUFx3_ASAP7_75t_L g406 ( .A(n_370), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_364), .B(n_335), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_377), .B(n_361), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_364), .B(n_334), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_353), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_361), .Y(n_411) );
CKINVDCx14_ASAP7_75t_R g412 ( .A(n_370), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_374), .A2(n_335), .B1(n_330), .B2(n_327), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_362), .Y(n_414) );
INVxp67_ASAP7_75t_SL g415 ( .A(n_364), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_367), .B(n_339), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_384), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_393), .B(n_357), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_393), .B(n_367), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_411), .B(n_362), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_407), .B(n_357), .Y(n_421) );
AO21x2_ASAP7_75t_L g422 ( .A1(n_413), .A2(n_358), .B(n_380), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_411), .B(n_377), .Y(n_423) );
INVx3_ASAP7_75t_L g424 ( .A(n_406), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_383), .Y(n_425) );
BUFx3_ASAP7_75t_L g426 ( .A(n_406), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_383), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_407), .B(n_357), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_390), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_381), .B(n_367), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_406), .B(n_370), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_381), .B(n_367), .Y(n_432) );
INVx3_ASAP7_75t_R g433 ( .A(n_412), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_392), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_381), .B(n_354), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_392), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_395), .Y(n_437) );
NOR2x1_ASAP7_75t_L g438 ( .A(n_406), .B(n_371), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_407), .B(n_371), .Y(n_439) );
AND2x4_ASAP7_75t_L g440 ( .A(n_385), .B(n_370), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_414), .B(n_371), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_385), .B(n_354), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_395), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_385), .B(n_360), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_389), .A2(n_365), .B1(n_405), .B2(n_373), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_384), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_414), .B(n_360), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_395), .B(n_371), .Y(n_448) );
AOI22xp33_ASAP7_75t_SL g449 ( .A1(n_412), .A2(n_370), .B1(n_360), .B2(n_369), .Y(n_449) );
INVx1_ASAP7_75t_SL g450 ( .A(n_390), .Y(n_450) );
INVx4_ASAP7_75t_L g451 ( .A(n_388), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_408), .B(n_374), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_408), .B(n_374), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_396), .B(n_380), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_396), .B(n_379), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_396), .B(n_379), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_399), .B(n_394), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_399), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_390), .B(n_365), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_399), .B(n_380), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_400), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_400), .Y(n_462) );
NOR2x1_ASAP7_75t_L g463 ( .A(n_402), .B(n_369), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_394), .B(n_380), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_402), .B(n_379), .Y(n_465) );
NOR2xp33_ASAP7_75t_R g466 ( .A(n_394), .B(n_370), .Y(n_466) );
AND2x4_ASAP7_75t_SL g467 ( .A(n_382), .B(n_376), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_459), .B(n_389), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_425), .Y(n_469) );
OR2x6_ASAP7_75t_L g470 ( .A(n_451), .B(n_431), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_435), .B(n_397), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_417), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_425), .Y(n_473) );
NAND3xp33_ASAP7_75t_SL g474 ( .A(n_445), .B(n_373), .C(n_405), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_427), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_457), .B(n_404), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_435), .B(n_397), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_457), .B(n_404), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_417), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_442), .B(n_397), .Y(n_480) );
NOR2x1p5_ASAP7_75t_L g481 ( .A(n_426), .B(n_415), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_427), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_442), .B(n_388), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_444), .B(n_388), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_434), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_450), .B(n_415), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_434), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_446), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_436), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_444), .B(n_382), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_436), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_446), .Y(n_492) );
INVx3_ASAP7_75t_L g493 ( .A(n_431), .Y(n_493) );
AND2x4_ASAP7_75t_L g494 ( .A(n_430), .B(n_409), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_429), .B(n_387), .Y(n_495) );
INVx3_ASAP7_75t_L g496 ( .A(n_431), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_437), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_466), .B(n_370), .Y(n_498) );
INVxp67_ASAP7_75t_L g499 ( .A(n_438), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_455), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_447), .B(n_403), .Y(n_501) );
INVx1_ASAP7_75t_SL g502 ( .A(n_426), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_447), .B(n_387), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_437), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_443), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_433), .B(n_370), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_443), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_461), .B(n_387), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_464), .B(n_403), .Y(n_509) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_463), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_461), .B(n_387), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_462), .B(n_384), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_458), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_464), .B(n_410), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_458), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_418), .B(n_384), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_462), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_454), .Y(n_518) );
AND3x2_ASAP7_75t_L g519 ( .A(n_433), .B(n_410), .C(n_370), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_454), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_455), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_418), .B(n_386), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_452), .B(n_413), .Y(n_523) );
INVx2_ASAP7_75t_SL g524 ( .A(n_451), .Y(n_524) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_451), .Y(n_525) );
INVx1_ASAP7_75t_SL g526 ( .A(n_440), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_430), .B(n_409), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_432), .B(n_409), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_490), .B(n_440), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_468), .B(n_419), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_469), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_518), .B(n_428), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_490), .B(n_440), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_524), .B(n_449), .Y(n_534) );
AND2x4_ASAP7_75t_L g535 ( .A(n_481), .B(n_424), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_480), .B(n_467), .Y(n_536) );
NAND2xp5_ASAP7_75t_R g537 ( .A(n_506), .B(n_419), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_469), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_523), .B(n_421), .Y(n_539) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_486), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_521), .B(n_421), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_474), .B(n_420), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_473), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_521), .B(n_428), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_518), .B(n_439), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_476), .B(n_422), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_478), .B(n_422), .Y(n_547) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_481), .A2(n_467), .B(n_424), .C(n_439), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_473), .Y(n_549) );
AOI21xp33_ASAP7_75t_SL g550 ( .A1(n_498), .A2(n_470), .B(n_524), .Y(n_550) );
OAI222xp33_ASAP7_75t_L g551 ( .A1(n_470), .A2(n_424), .B1(n_448), .B2(n_453), .C1(n_386), .C2(n_376), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_470), .A2(n_422), .B1(n_423), .B2(n_432), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_494), .B(n_460), .Y(n_553) );
INVxp67_ASAP7_75t_L g554 ( .A(n_525), .Y(n_554) );
INVxp67_ASAP7_75t_L g555 ( .A(n_510), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_494), .B(n_460), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_475), .Y(n_557) );
INVx2_ASAP7_75t_SL g558 ( .A(n_519), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_475), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_482), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_482), .Y(n_561) );
XNOR2x1_ASAP7_75t_L g562 ( .A(n_502), .B(n_448), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_485), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_499), .B(n_441), .Y(n_564) );
NAND2x1_ASAP7_75t_L g565 ( .A(n_470), .B(n_376), .Y(n_565) );
NOR2x1_ASAP7_75t_L g566 ( .A(n_470), .B(n_376), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_493), .B(n_456), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_493), .A2(n_376), .B1(n_456), .B2(n_465), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_480), .B(n_465), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_485), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_494), .B(n_401), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_494), .B(n_401), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_483), .B(n_401), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_487), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_493), .A2(n_376), .B1(n_378), .B2(n_398), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_487), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_518), .B(n_398), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_483), .B(n_398), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_489), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_527), .B(n_416), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_489), .Y(n_581) );
OAI22xp33_ASAP7_75t_L g582 ( .A1(n_565), .A2(n_496), .B1(n_493), .B2(n_526), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_569), .B(n_496), .Y(n_583) );
AOI21xp33_ASAP7_75t_SL g584 ( .A1(n_534), .A2(n_496), .B(n_486), .Y(n_584) );
XNOR2xp5_ASAP7_75t_L g585 ( .A(n_562), .B(n_528), .Y(n_585) );
INVx1_ASAP7_75t_SL g586 ( .A(n_540), .Y(n_586) );
INVx2_ASAP7_75t_SL g587 ( .A(n_529), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_541), .Y(n_588) );
OAI211xp5_ASAP7_75t_SL g589 ( .A1(n_542), .A2(n_496), .B(n_522), .C(n_495), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_544), .Y(n_590) );
NOR3xp33_ASAP7_75t_SL g591 ( .A(n_534), .B(n_503), .C(n_491), .Y(n_591) );
INVx2_ASAP7_75t_SL g592 ( .A(n_533), .Y(n_592) );
NOR2xp67_ASAP7_75t_L g593 ( .A(n_550), .B(n_520), .Y(n_593) );
INVx1_ASAP7_75t_SL g594 ( .A(n_540), .Y(n_594) );
AOI31xp33_ASAP7_75t_L g595 ( .A1(n_566), .A2(n_471), .A3(n_477), .B(n_484), .Y(n_595) );
INVx2_ASAP7_75t_SL g596 ( .A(n_535), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_546), .B(n_528), .Y(n_597) );
AOI222xp33_ASAP7_75t_L g598 ( .A1(n_542), .A2(n_484), .B1(n_471), .B2(n_477), .C1(n_501), .C2(n_514), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_548), .A2(n_501), .B1(n_509), .B2(n_514), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_531), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_532), .B(n_545), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_530), .B(n_500), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_567), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_555), .B(n_500), .Y(n_604) );
AOI322xp5_ASAP7_75t_L g605 ( .A1(n_539), .A2(n_527), .A3(n_509), .B1(n_520), .B2(n_517), .C1(n_491), .C2(n_505), .Y(n_605) );
OAI21xp5_ASAP7_75t_L g606 ( .A1(n_567), .A2(n_376), .B(n_517), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_548), .A2(n_522), .B1(n_516), .B2(n_520), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_580), .B(n_516), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_554), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_564), .A2(n_515), .B1(n_513), .B2(n_497), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g611 ( .A1(n_547), .A2(n_515), .B1(n_513), .B2(n_497), .C(n_504), .Y(n_611) );
NAND3xp33_ASAP7_75t_L g612 ( .A(n_555), .B(n_507), .C(n_505), .Y(n_612) );
OA21x2_ASAP7_75t_SL g613 ( .A1(n_535), .A2(n_512), .B(n_511), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_558), .B(n_472), .Y(n_614) );
NAND3x2_ASAP7_75t_L g615 ( .A(n_536), .B(n_507), .C(n_504), .Y(n_615) );
O2A1O1Ixp5_ASAP7_75t_L g616 ( .A1(n_551), .A2(n_508), .B(n_472), .C(n_488), .Y(n_616) );
AOI222xp33_ASAP7_75t_L g617 ( .A1(n_551), .A2(n_492), .B1(n_488), .B2(n_479), .C1(n_378), .C2(n_416), .Y(n_617) );
AOI322xp5_ASAP7_75t_L g618 ( .A1(n_591), .A2(n_578), .A3(n_573), .B1(n_556), .B2(n_553), .C1(n_554), .C2(n_552), .Y(n_618) );
A2O1A1Ixp33_ASAP7_75t_L g619 ( .A1(n_584), .A2(n_564), .B(n_568), .C(n_571), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g620 ( .A1(n_606), .A2(n_575), .B(n_572), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_605), .B(n_581), .Y(n_621) );
OAI221xp5_ASAP7_75t_L g622 ( .A1(n_616), .A2(n_579), .B1(n_549), .B2(n_576), .C(n_574), .Y(n_622) );
OAI21xp33_ASAP7_75t_L g623 ( .A1(n_589), .A2(n_537), .B(n_570), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_600), .Y(n_624) );
OAI211xp5_ASAP7_75t_L g625 ( .A1(n_615), .A2(n_559), .B(n_563), .C(n_561), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_608), .Y(n_626) );
OAI31xp33_ASAP7_75t_L g627 ( .A1(n_582), .A2(n_560), .A3(n_557), .B(n_543), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_599), .A2(n_538), .B1(n_577), .B2(n_492), .Y(n_628) );
O2A1O1Ixp33_ASAP7_75t_L g629 ( .A1(n_595), .A2(n_348), .B(n_488), .C(n_479), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_612), .Y(n_630) );
AOI222xp33_ASAP7_75t_L g631 ( .A1(n_607), .A2(n_492), .B1(n_479), .B2(n_416), .C1(n_379), .C2(n_352), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_601), .Y(n_632) );
OAI322xp33_ASAP7_75t_SL g633 ( .A1(n_597), .A2(n_391), .A3(n_372), .B1(n_352), .B2(n_63), .C1(n_64), .C2(n_65), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_598), .B(n_391), .Y(n_634) );
INVx1_ASAP7_75t_SL g635 ( .A(n_586), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_606), .A2(n_391), .B(n_352), .Y(n_636) );
AND2x2_ASAP7_75t_SL g637 ( .A(n_613), .B(n_391), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_609), .Y(n_638) );
AOI222xp33_ASAP7_75t_L g639 ( .A1(n_607), .A2(n_391), .B1(n_372), .B2(n_62), .C1(n_66), .C2(n_67), .Y(n_639) );
NOR3xp33_ASAP7_75t_L g640 ( .A(n_630), .B(n_599), .C(n_614), .Y(n_640) );
OAI222xp33_ASAP7_75t_L g641 ( .A1(n_634), .A2(n_585), .B1(n_596), .B2(n_594), .C1(n_603), .C2(n_590), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_635), .B(n_588), .Y(n_642) );
OAI221xp5_ASAP7_75t_SL g643 ( .A1(n_618), .A2(n_617), .B1(n_610), .B2(n_611), .C(n_597), .Y(n_643) );
A2O1A1Ixp33_ASAP7_75t_L g644 ( .A1(n_619), .A2(n_593), .B(n_604), .C(n_602), .Y(n_644) );
NOR2x1_ASAP7_75t_L g645 ( .A(n_625), .B(n_583), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_632), .Y(n_646) );
NAND4xp25_ASAP7_75t_L g647 ( .A(n_639), .B(n_611), .C(n_592), .D(n_587), .Y(n_647) );
NOR3xp33_ASAP7_75t_L g648 ( .A(n_623), .B(n_59), .C(n_60), .Y(n_648) );
NOR4xp25_ASAP7_75t_SL g649 ( .A(n_622), .B(n_391), .C(n_372), .D(n_74), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_621), .B(n_372), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_626), .Y(n_651) );
OAI21xp5_ASAP7_75t_L g652 ( .A1(n_627), .A2(n_372), .B(n_72), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_646), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_640), .A2(n_637), .B1(n_628), .B2(n_631), .Y(n_654) );
OAI321xp33_ASAP7_75t_L g655 ( .A1(n_643), .A2(n_620), .A3(n_638), .B1(n_636), .B2(n_629), .C(n_624), .Y(n_655) );
OAI22xp33_ASAP7_75t_L g656 ( .A1(n_647), .A2(n_620), .B1(n_636), .B2(n_633), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_642), .Y(n_657) );
NOR4xp25_ASAP7_75t_L g658 ( .A(n_641), .B(n_372), .C(n_76), .D(n_78), .Y(n_658) );
NAND4xp25_ASAP7_75t_L g659 ( .A(n_648), .B(n_70), .C(n_80), .D(n_82), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_657), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_654), .A2(n_644), .B1(n_645), .B2(n_650), .Y(n_661) );
NAND4xp25_ASAP7_75t_L g662 ( .A(n_659), .B(n_652), .C(n_642), .D(n_651), .Y(n_662) );
OR2x2_ASAP7_75t_L g663 ( .A(n_653), .B(n_656), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_660), .Y(n_664) );
OAI22x1_ASAP7_75t_L g665 ( .A1(n_663), .A2(n_655), .B1(n_658), .B2(n_649), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_661), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_664), .Y(n_667) );
INVx3_ASAP7_75t_L g668 ( .A(n_666), .Y(n_668) );
AOI22x1_ASAP7_75t_L g669 ( .A1(n_668), .A2(n_666), .B1(n_665), .B2(n_662), .Y(n_669) );
AOI221xp5_ASAP7_75t_L g670 ( .A1(n_669), .A2(n_668), .B1(n_667), .B2(n_89), .C(n_85), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_670), .B(n_668), .Y(n_671) );
OA21x2_ASAP7_75t_L g672 ( .A1(n_671), .A2(n_667), .B(n_668), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_672), .A2(n_668), .B1(n_667), .B2(n_84), .Y(n_673) );
endmodule