module fake_jpeg_1948_n_618 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_618);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_618;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_12),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_17),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_58),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_59),
.Y(n_146)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_60),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_21),
.B(n_19),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_61),
.B(n_62),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_18),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_63),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_64),
.Y(n_174)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_66),
.B(n_89),
.Y(n_136)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_67),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_68),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_69),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_18),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_70),
.B(n_71),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_37),
.B(n_0),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_72),
.Y(n_182)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_73),
.Y(n_144)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g156 ( 
.A(n_74),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_75),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_76),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_77),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_78),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_41),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_79),
.A2(n_14),
.B1(n_15),
.B2(n_121),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_80),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_0),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_81),
.B(n_93),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_82),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_83),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_84),
.Y(n_209)
);

INVx3_ASAP7_75t_SL g85 ( 
.A(n_38),
.Y(n_85)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

INVx2_ASAP7_75t_R g86 ( 
.A(n_38),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_86),
.B(n_105),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_88),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_48),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_90),
.Y(n_178)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_91),
.Y(n_185)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_0),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_95),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

AOI21xp33_ASAP7_75t_L g97 ( 
.A1(n_56),
.A2(n_1),
.B(n_2),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_97),
.B(n_106),
.Y(n_145)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

BUFx12_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_99),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_2),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_100),
.B(n_101),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_54),
.B(n_28),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_103),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_27),
.Y(n_104)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_104),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_22),
.B(n_2),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_54),
.B(n_5),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_35),
.Y(n_107)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_107),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_28),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_108),
.B(n_113),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_31),
.Y(n_109)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_109),
.Y(n_152)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_110),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_27),
.Y(n_111)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_111),
.Y(n_197)
);

BUFx12_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

BUFx4f_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_27),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_32),
.B(n_36),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_114),
.B(n_116),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_30),
.Y(n_115)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_115),
.Y(n_200)
);

BUFx12_ASAP7_75t_L g116 ( 
.A(n_29),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_35),
.Y(n_117)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_117),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_42),
.Y(n_118)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_118),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_30),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_129),
.Y(n_155)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_120),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_44),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_128),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_30),
.Y(n_122)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_46),
.Y(n_123)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_123),
.Y(n_164)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_42),
.Y(n_124)
);

NAND2xp33_ASAP7_75t_SL g140 ( 
.A(n_124),
.B(n_125),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_29),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_46),
.Y(n_126)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_126),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_46),
.Y(n_127)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_127),
.Y(n_186)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_42),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_44),
.Y(n_129)
);

AO22x1_ASAP7_75t_SL g135 ( 
.A1(n_67),
.A2(n_51),
.B1(n_52),
.B2(n_24),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_135),
.B(n_216),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_68),
.A2(n_24),
.B1(n_52),
.B2(n_51),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_139),
.A2(n_148),
.B1(n_157),
.B2(n_165),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_79),
.A2(n_123),
.B1(n_104),
.B2(n_127),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_85),
.A2(n_51),
.B1(n_52),
.B2(n_24),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_150),
.B(n_176),
.Y(n_282)
);

NAND2xp33_ASAP7_75t_SL g153 ( 
.A(n_86),
.B(n_75),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_L g290 ( 
.A1(n_153),
.A2(n_180),
.B(n_179),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_111),
.A2(n_22),
.B1(n_40),
.B2(n_34),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_115),
.A2(n_23),
.B1(n_40),
.B2(n_34),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_162),
.A2(n_189),
.B1(n_196),
.B2(n_215),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_122),
.A2(n_45),
.B1(n_32),
.B2(n_39),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_108),
.B(n_26),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_166),
.B(n_171),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_126),
.A2(n_26),
.B1(n_25),
.B2(n_23),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_179),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_76),
.A2(n_45),
.B1(n_39),
.B2(n_36),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_59),
.A2(n_25),
.B1(n_44),
.B2(n_8),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_64),
.B(n_6),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_64),
.B(n_6),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_175),
.B(n_177),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_94),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_63),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_92),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_98),
.A2(n_124),
.B1(n_118),
.B2(n_96),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_180),
.A2(n_184),
.B1(n_217),
.B2(n_219),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_72),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_181),
.A2(n_193),
.B1(n_169),
.B2(n_184),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_109),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_77),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_69),
.B(n_13),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_194),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_78),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_95),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_80),
.A2(n_90),
.B1(n_87),
.B2(n_82),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_120),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_202),
.Y(n_231)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_83),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_84),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_203),
.B(n_204),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_69),
.B(n_14),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_128),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_206),
.B(n_212),
.Y(n_251)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_110),
.Y(n_212)
);

OA22x2_ASAP7_75t_L g216 ( 
.A1(n_116),
.A2(n_73),
.B1(n_99),
.B2(n_112),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_140),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_121),
.A2(n_129),
.B1(n_116),
.B2(n_73),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_99),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_220),
.B(n_221),
.Y(n_270)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_112),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_129),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_223),
.B(n_188),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_61),
.A2(n_70),
.B1(n_106),
.B2(n_105),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_224),
.A2(n_183),
.B1(n_162),
.B2(n_149),
.Y(n_245)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_164),
.Y(n_228)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_228),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_230),
.B(n_262),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_130),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_232),
.Y(n_340)
);

INVx13_ASAP7_75t_L g233 ( 
.A(n_219),
.Y(n_233)
);

BUFx24_ASAP7_75t_L g317 ( 
.A(n_233),
.Y(n_317)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_135),
.Y(n_234)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_234),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_235),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_158),
.B(n_170),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_236),
.B(n_238),
.Y(n_313)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_237),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_136),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_239),
.Y(n_353)
);

FAx1_ASAP7_75t_SL g240 ( 
.A(n_145),
.B(n_137),
.CI(n_195),
.CON(n_240),
.SN(n_240)
);

FAx1_ASAP7_75t_SL g339 ( 
.A(n_240),
.B(n_227),
.CI(n_238),
.CON(n_339),
.SN(n_339)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_207),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_242),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_154),
.B(n_134),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_243),
.B(n_267),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_244),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_245),
.A2(n_248),
.B1(n_249),
.B2(n_240),
.Y(n_334)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_142),
.Y(n_246)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_246),
.Y(n_367)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_197),
.Y(n_247)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_247),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_155),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_249),
.B(n_254),
.Y(n_320)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_135),
.Y(n_250)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_250),
.Y(n_338)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_200),
.Y(n_252)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_252),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_137),
.A2(n_211),
.B1(n_130),
.B2(n_210),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_253),
.A2(n_279),
.B1(n_288),
.B2(n_295),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_211),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_216),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_256),
.B(n_261),
.Y(n_332)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_147),
.Y(n_257)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_257),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_146),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_258),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_173),
.B(n_190),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_259),
.Y(n_342)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_172),
.Y(n_260)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_260),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_163),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_185),
.B(n_163),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_186),
.Y(n_263)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_263),
.Y(n_351)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_208),
.Y(n_264)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_264),
.Y(n_358)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_208),
.Y(n_265)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_265),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_159),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_266),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_131),
.B(n_189),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_192),
.B(n_201),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_268),
.B(n_274),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_139),
.A2(n_168),
.B(n_217),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_269),
.A2(n_290),
.B(n_244),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_146),
.Y(n_271)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_271),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_272),
.B(n_273),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_161),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_218),
.Y(n_274)
);

INVx13_ASAP7_75t_L g275 ( 
.A(n_188),
.Y(n_275)
);

INVx11_ASAP7_75t_L g315 ( 
.A(n_275),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_276),
.A2(n_301),
.B1(n_302),
.B2(n_229),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_141),
.B(n_214),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_277),
.B(n_280),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_165),
.B(n_181),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_278),
.B(n_283),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_222),
.A2(n_152),
.B1(n_138),
.B2(n_132),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_161),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_178),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_281),
.Y(n_356)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_144),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_138),
.B(n_152),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_284),
.B(n_285),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_187),
.B(n_205),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_144),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_286),
.B(n_287),
.Y(n_362)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_133),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_222),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_159),
.Y(n_289)
);

BUFx5_ASAP7_75t_L g324 ( 
.A(n_289),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_156),
.B(n_188),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_291),
.B(n_292),
.Y(n_363)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_133),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_156),
.B(n_160),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_293),
.B(n_294),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_187),
.B(n_209),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_143),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_226),
.A2(n_160),
.B1(n_143),
.B2(n_178),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_296),
.A2(n_300),
.B1(n_303),
.B2(n_305),
.Y(n_346)
);

HAxp5_ASAP7_75t_SL g297 ( 
.A(n_174),
.B(n_226),
.CON(n_297),
.SN(n_297)
);

FAx1_ASAP7_75t_L g336 ( 
.A(n_297),
.B(n_309),
.CI(n_282),
.CON(n_336),
.SN(n_336)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_205),
.B(n_209),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_298),
.B(n_304),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_174),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_151),
.A2(n_182),
.B1(n_198),
.B2(n_213),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_151),
.A2(n_182),
.B1(n_198),
.B2(n_213),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_225),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_225),
.B(n_145),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_154),
.B(n_195),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_164),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_306),
.A2(n_308),
.B1(n_280),
.B2(n_281),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_154),
.B(n_195),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_309),
.C(n_243),
.Y(n_321)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_207),
.Y(n_308)
);

A2O1A1Ixp33_ASAP7_75t_L g309 ( 
.A1(n_145),
.A2(n_137),
.B(n_195),
.C(n_170),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_234),
.A2(n_250),
.B1(n_255),
.B2(n_267),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_311),
.A2(n_314),
.B1(n_330),
.B2(n_350),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_255),
.A2(n_276),
.B1(n_278),
.B2(n_230),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_316),
.A2(n_325),
.B1(n_341),
.B2(n_345),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_318),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_321),
.B(n_246),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_310),
.A2(n_261),
.B1(n_269),
.B2(n_304),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_282),
.A2(n_244),
.B1(n_294),
.B2(n_298),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_333),
.A2(n_358),
.B(n_353),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_334),
.B(n_319),
.Y(n_395)
);

MAJx2_ASAP7_75t_L g335 ( 
.A(n_240),
.B(n_299),
.C(n_262),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_335),
.B(n_274),
.C(n_306),
.Y(n_378)
);

CKINVDCx14_ASAP7_75t_R g397 ( 
.A(n_336),
.Y(n_397)
);

BUFx24_ASAP7_75t_SL g371 ( 
.A(n_339),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_285),
.A2(n_268),
.B1(n_302),
.B2(n_301),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_241),
.A2(n_262),
.B1(n_284),
.B2(n_259),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_259),
.A2(n_257),
.B1(n_303),
.B2(n_273),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_228),
.A2(n_265),
.B1(n_264),
.B2(n_252),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_359),
.A2(n_369),
.B1(n_286),
.B2(n_283),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_297),
.A2(n_251),
.B(n_231),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_368),
.A2(n_346),
.B(n_329),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_247),
.A2(n_263),
.B1(n_260),
.B2(n_271),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_362),
.Y(n_370)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_370),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_321),
.B(n_270),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_373),
.B(n_388),
.Y(n_427)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_362),
.Y(n_374)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_374),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_363),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_375),
.B(n_376),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_359),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_343),
.A2(n_288),
.B1(n_239),
.B2(n_237),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_377),
.A2(n_409),
.B(n_413),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_378),
.B(n_380),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_340),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_379),
.B(n_386),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_352),
.B(n_295),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_381),
.B(n_393),
.C(n_344),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_316),
.A2(n_258),
.B1(n_242),
.B2(n_308),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_383),
.A2(n_385),
.B1(n_390),
.B2(n_400),
.Y(n_449)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_384),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_314),
.A2(n_287),
.B1(n_292),
.B2(n_289),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_340),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_313),
.B(n_266),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_R g389 ( 
.A(n_332),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_389),
.B(n_394),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_323),
.A2(n_233),
.B1(n_275),
.B2(n_338),
.Y(n_390)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_315),
.Y(n_391)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_391),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_368),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_392),
.B(n_395),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_352),
.B(n_357),
.C(n_335),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_320),
.B(n_337),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_327),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_396),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_311),
.A2(n_330),
.B1(n_323),
.B2(n_338),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_398),
.A2(n_404),
.B1(n_405),
.B2(n_408),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_333),
.B(n_342),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_399),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_357),
.A2(n_319),
.B1(n_355),
.B2(n_349),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_347),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_401),
.B(n_406),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_363),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_402),
.B(n_403),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_361),
.B(n_345),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_357),
.A2(n_349),
.B1(n_341),
.B2(n_355),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_365),
.A2(n_336),
.B1(n_366),
.B2(n_331),
.Y(n_405)
);

AO22x1_ASAP7_75t_L g406 ( 
.A1(n_336),
.A2(n_350),
.B1(n_347),
.B2(n_369),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_331),
.B(n_365),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_407),
.B(n_348),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_366),
.A2(n_356),
.B1(n_312),
.B2(n_360),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_317),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_410),
.Y(n_426)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_312),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_411),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_358),
.B(n_360),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_412),
.Y(n_450)
);

INVx8_ASAP7_75t_L g414 ( 
.A(n_354),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_414),
.A2(n_415),
.B(n_410),
.Y(n_422)
);

CKINVDCx14_ASAP7_75t_R g415 ( 
.A(n_317),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_393),
.B(n_339),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_419),
.B(n_423),
.C(n_437),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_422),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_372),
.A2(n_339),
.B1(n_364),
.B2(n_353),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_430),
.A2(n_431),
.B1(n_432),
.B2(n_452),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_372),
.A2(n_364),
.B1(n_354),
.B2(n_351),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_404),
.A2(n_351),
.B1(n_348),
.B2(n_328),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_434),
.B(n_401),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_382),
.A2(n_326),
.B1(n_322),
.B2(n_367),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_436),
.A2(n_442),
.B1(n_449),
.B2(n_421),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_381),
.B(n_367),
.C(n_326),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_413),
.A2(n_315),
.B(n_317),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_438),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_397),
.A2(n_324),
.B(n_327),
.Y(n_439)
);

OA21x2_ASAP7_75t_L g484 ( 
.A1(n_439),
.A2(n_454),
.B(n_391),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_378),
.B(n_322),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_440),
.B(n_441),
.C(n_444),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_407),
.B(n_400),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_382),
.A2(n_324),
.B1(n_398),
.B2(n_405),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_380),
.B(n_399),
.C(n_395),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_399),
.B(n_395),
.C(n_403),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_447),
.B(n_453),
.C(n_414),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_370),
.A2(n_374),
.B1(n_376),
.B2(n_389),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_373),
.B(n_375),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_409),
.A2(n_392),
.B(n_406),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_443),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_455),
.Y(n_499)
);

OAI32xp33_ASAP7_75t_L g456 ( 
.A1(n_424),
.A2(n_406),
.A3(n_402),
.B1(n_394),
.B2(n_387),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_456),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_424),
.B(n_408),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_457),
.A2(n_459),
.B1(n_469),
.B2(n_475),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_433),
.A2(n_385),
.B1(n_383),
.B2(n_388),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_458),
.A2(n_484),
.B(n_418),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_SL g459 ( 
.A1(n_421),
.A2(n_390),
.B1(n_379),
.B2(n_386),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_450),
.B(n_412),
.Y(n_461)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_461),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_448),
.B(n_371),
.Y(n_462)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_462),
.Y(n_492)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_443),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_SL g510 ( 
.A(n_465),
.B(n_471),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_450),
.B(n_411),
.Y(n_466)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_466),
.Y(n_505)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_432),
.Y(n_467)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_467),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_448),
.B(n_377),
.Y(n_468)
);

OR2x2_ASAP7_75t_L g518 ( 
.A(n_468),
.B(n_470),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_427),
.B(n_396),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_428),
.B(n_384),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_452),
.B(n_415),
.Y(n_472)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_472),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_428),
.B(n_396),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_473),
.B(n_487),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_422),
.Y(n_474)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_474),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_442),
.A2(n_391),
.B1(n_414),
.B2(n_417),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_417),
.Y(n_476)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_425),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g517 ( 
.A(n_479),
.Y(n_517)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_420),
.Y(n_480)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_480),
.Y(n_508)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_420),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_482),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_434),
.B(n_441),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_483),
.Y(n_507)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_446),
.Y(n_485)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_485),
.Y(n_504)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_431),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_486),
.A2(n_488),
.B1(n_490),
.B2(n_449),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_427),
.B(n_451),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_423),
.B(n_440),
.C(n_444),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_489),
.B(n_437),
.C(n_419),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_451),
.B(n_447),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_467),
.A2(n_429),
.B1(n_446),
.B2(n_430),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_493),
.A2(n_495),
.B1(n_509),
.B2(n_512),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_481),
.B(n_453),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_494),
.B(n_497),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_486),
.A2(n_429),
.B1(n_464),
.B2(n_475),
.Y(n_495)
);

XNOR2x1_ASAP7_75t_L g497 ( 
.A(n_471),
.B(n_454),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_502),
.B(n_477),
.C(n_489),
.Y(n_522)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_506),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_464),
.A2(n_435),
.B1(n_436),
.B2(n_439),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_463),
.A2(n_435),
.B1(n_441),
.B2(n_445),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_478),
.A2(n_418),
.B1(n_426),
.B2(n_445),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_513),
.B(n_514),
.Y(n_526)
);

XNOR2x1_ASAP7_75t_L g514 ( 
.A(n_473),
.B(n_419),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_515),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_478),
.A2(n_438),
.B(n_426),
.Y(n_516)
);

CKINVDCx14_ASAP7_75t_R g536 ( 
.A(n_516),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_455),
.A2(n_457),
.B1(n_484),
.B2(n_472),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_519),
.A2(n_520),
.B1(n_479),
.B2(n_425),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_458),
.A2(n_460),
.B1(n_456),
.B2(n_466),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_522),
.B(n_537),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_491),
.B(n_481),
.C(n_477),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_523),
.B(n_527),
.C(n_531),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_499),
.B(n_461),
.Y(n_525)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_525),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_491),
.B(n_487),
.C(n_483),
.Y(n_527)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_503),
.Y(n_529)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_529),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_492),
.B(n_488),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_530),
.B(n_535),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_502),
.B(n_465),
.C(n_460),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_507),
.B(n_490),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_SL g562 ( 
.A(n_533),
.B(n_534),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_518),
.B(n_416),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_518),
.B(n_476),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_494),
.B(n_484),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_508),
.Y(n_538)
);

BUFx4f_ASAP7_75t_SL g552 ( 
.A(n_538),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_514),
.B(n_480),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_510),
.B(n_482),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g564 ( 
.A1(n_541),
.A2(n_519),
.B(n_509),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_496),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_542),
.Y(n_547)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_508),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_543),
.B(n_544),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_496),
.B(n_504),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_497),
.B(n_510),
.C(n_501),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_546),
.B(n_512),
.C(n_505),
.Y(n_556)
);

INVxp33_ASAP7_75t_SL g548 ( 
.A(n_528),
.Y(n_548)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_548),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_524),
.B(n_520),
.Y(n_551)
);

MAJx2_ASAP7_75t_L g566 ( 
.A(n_551),
.B(n_556),
.C(n_559),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_527),
.B(n_516),
.C(n_513),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_558),
.B(n_563),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_522),
.B(n_531),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_524),
.B(n_515),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_560),
.B(n_546),
.C(n_545),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_545),
.B(n_511),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_SL g577 ( 
.A(n_561),
.B(n_504),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_523),
.B(n_537),
.C(n_539),
.Y(n_563)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_564),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_565),
.B(n_563),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_559),
.B(n_536),
.C(n_526),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_568),
.B(n_571),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_564),
.A2(n_532),
.B1(n_500),
.B2(n_511),
.Y(n_570)
);

INVxp33_ASAP7_75t_L g588 ( 
.A(n_570),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_562),
.B(n_532),
.Y(n_571)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_558),
.A2(n_526),
.B(n_521),
.Y(n_572)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_572),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_554),
.B(n_526),
.C(n_540),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_573),
.B(n_574),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_554),
.B(n_498),
.C(n_495),
.Y(n_574)
);

NOR2x1_ASAP7_75t_SL g576 ( 
.A(n_556),
.B(n_521),
.Y(n_576)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_576),
.Y(n_587)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_577),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_549),
.B(n_493),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_SL g593 ( 
.A(n_578),
.B(n_569),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_553),
.A2(n_505),
.B1(n_508),
.B2(n_517),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_579),
.B(n_580),
.Y(n_581)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_547),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_582),
.B(n_573),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_574),
.B(n_550),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_586),
.B(n_589),
.Y(n_598)
);

FAx1_ASAP7_75t_SL g589 ( 
.A(n_568),
.B(n_560),
.CI(n_551),
.CON(n_589),
.SN(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_567),
.B(n_555),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_590),
.B(n_593),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_580),
.B(n_547),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_L g597 ( 
.A1(n_592),
.A2(n_576),
.B(n_567),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_SL g594 ( 
.A(n_582),
.B(n_575),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_594),
.B(n_596),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g603 ( 
.A1(n_595),
.A2(n_599),
.B(n_572),
.Y(n_603)
);

XNOR2xp5_ASAP7_75t_L g596 ( 
.A(n_584),
.B(n_566),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_SL g607 ( 
.A1(n_597),
.A2(n_601),
.B(n_592),
.Y(n_607)
);

NOR2xp67_ASAP7_75t_SL g599 ( 
.A(n_583),
.B(n_565),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_591),
.B(n_552),
.Y(n_601)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_585),
.B(n_557),
.Y(n_602)
);

XOR2xp5_ASAP7_75t_L g604 ( 
.A(n_602),
.B(n_566),
.Y(n_604)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_603),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_604),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_598),
.B(n_587),
.Y(n_605)
);

BUFx24_ASAP7_75t_SL g611 ( 
.A(n_605),
.Y(n_611)
);

FAx1_ASAP7_75t_SL g612 ( 
.A(n_607),
.B(n_608),
.CI(n_601),
.CON(n_612),
.SN(n_612)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_595),
.A2(n_581),
.B(n_588),
.Y(n_608)
);

OAI21xp5_ASAP7_75t_L g613 ( 
.A1(n_612),
.A2(n_606),
.B(n_609),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_613),
.A2(n_614),
.B(n_611),
.Y(n_615)
);

OAI21xp5_ASAP7_75t_L g614 ( 
.A1(n_610),
.A2(n_600),
.B(n_581),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_615),
.Y(n_616)
);

XOR2xp5_ASAP7_75t_L g617 ( 
.A(n_616),
.B(n_588),
.Y(n_617)
);

XOR2xp5_ASAP7_75t_L g618 ( 
.A(n_617),
.B(n_570),
.Y(n_618)
);


endmodule