module fake_netlist_1_10004_n_642 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_642);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_642;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_624;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_295;
wire n_143;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_54), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_15), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_33), .Y(n_79) );
INVx2_ASAP7_75t_L g80 ( .A(n_30), .Y(n_80) );
BUFx6f_ASAP7_75t_L g81 ( .A(n_64), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_32), .Y(n_82) );
INVxp67_ASAP7_75t_SL g83 ( .A(n_8), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_15), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_51), .Y(n_85) );
INVxp33_ASAP7_75t_SL g86 ( .A(n_66), .Y(n_86) );
NOR2xp67_ASAP7_75t_L g87 ( .A(n_35), .B(n_39), .Y(n_87) );
BUFx3_ASAP7_75t_L g88 ( .A(n_69), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_42), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_45), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_27), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_34), .Y(n_92) );
NOR2xp67_ASAP7_75t_L g93 ( .A(n_4), .B(n_58), .Y(n_93) );
INVxp67_ASAP7_75t_L g94 ( .A(n_25), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_14), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_14), .Y(n_96) );
BUFx2_ASAP7_75t_L g97 ( .A(n_65), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_55), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_37), .Y(n_99) );
CKINVDCx14_ASAP7_75t_R g100 ( .A(n_72), .Y(n_100) );
BUFx6f_ASAP7_75t_L g101 ( .A(n_44), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_60), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_17), .Y(n_103) );
BUFx3_ASAP7_75t_L g104 ( .A(n_21), .Y(n_104) );
BUFx6f_ASAP7_75t_L g105 ( .A(n_36), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_43), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_20), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_28), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_56), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_46), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_12), .Y(n_111) );
INVx3_ASAP7_75t_L g112 ( .A(n_75), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_47), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_5), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_40), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_8), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_2), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_5), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_73), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_117), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_97), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_112), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_97), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_100), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_77), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_117), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_112), .B(n_0), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_81), .Y(n_128) );
AOI22xp5_ASAP7_75t_L g129 ( .A1(n_78), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_77), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_112), .B(n_1), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_79), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_81), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_112), .B(n_3), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_80), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_80), .B(n_3), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_110), .B(n_4), .Y(n_137) );
AND2x2_ASAP7_75t_SL g138 ( .A(n_79), .B(n_76), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_85), .Y(n_139) );
INVxp67_ASAP7_75t_SL g140 ( .A(n_95), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_110), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_85), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_81), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_89), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_89), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_90), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_90), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_81), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_92), .Y(n_149) );
AND2x4_ASAP7_75t_L g150 ( .A(n_95), .B(n_6), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_96), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_103), .Y(n_152) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_116), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_103), .B(n_6), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_92), .Y(n_155) );
BUFx10_ASAP7_75t_L g156 ( .A(n_124), .Y(n_156) );
INVx4_ASAP7_75t_L g157 ( .A(n_150), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_128), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_128), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_150), .Y(n_160) );
INVx3_ASAP7_75t_L g161 ( .A(n_150), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_122), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_120), .B(n_78), .Y(n_163) );
NAND2x1p5_ASAP7_75t_L g164 ( .A(n_138), .B(n_119), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_122), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_120), .B(n_118), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_128), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_121), .B(n_118), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_128), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_124), .B(n_94), .Y(n_170) );
BUFx2_ASAP7_75t_L g171 ( .A(n_126), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_150), .Y(n_172) );
OR2x2_ASAP7_75t_SL g173 ( .A(n_123), .B(n_114), .Y(n_173) );
INVx2_ASAP7_75t_SL g174 ( .A(n_125), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_153), .B(n_86), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_128), .Y(n_176) );
BUFx3_ASAP7_75t_L g177 ( .A(n_135), .Y(n_177) );
AND2x2_ASAP7_75t_L g178 ( .A(n_140), .B(n_114), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_126), .B(n_104), .Y(n_179) );
AND2x4_ASAP7_75t_L g180 ( .A(n_125), .B(n_84), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_135), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_141), .Y(n_182) );
INVx4_ASAP7_75t_L g183 ( .A(n_138), .Y(n_183) );
NOR2xp33_ASAP7_75t_R g184 ( .A(n_151), .B(n_138), .Y(n_184) );
HB1xp67_ASAP7_75t_L g185 ( .A(n_151), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_141), .Y(n_186) );
BUFx10_ASAP7_75t_L g187 ( .A(n_127), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_133), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_144), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_144), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_130), .B(n_107), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_130), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_132), .B(n_139), .Y(n_193) );
INVx1_ASAP7_75t_SL g194 ( .A(n_154), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_132), .Y(n_195) );
INVx2_ASAP7_75t_SL g196 ( .A(n_139), .Y(n_196) );
AO22x2_ASAP7_75t_L g197 ( .A1(n_142), .A2(n_119), .B1(n_113), .B2(n_98), .Y(n_197) );
AO21x1_ASAP7_75t_L g198 ( .A1(n_164), .A2(n_131), .B(n_134), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g199 ( .A1(n_183), .A2(n_154), .B1(n_155), .B2(n_142), .Y(n_199) );
INVx2_ASAP7_75t_SL g200 ( .A(n_194), .Y(n_200) );
AND2x4_ASAP7_75t_L g201 ( .A(n_194), .B(n_129), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_178), .B(n_145), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_183), .A2(n_155), .B1(n_145), .B2(n_149), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_178), .B(n_149), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_189), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_189), .Y(n_206) );
NAND3xp33_ASAP7_75t_SL g207 ( .A(n_184), .B(n_111), .C(n_115), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_162), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_157), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_162), .Y(n_210) );
O2A1O1Ixp5_ASAP7_75t_L g211 ( .A1(n_157), .A2(n_136), .B(n_137), .C(n_147), .Y(n_211) );
NOR2x1_ASAP7_75t_R g212 ( .A(n_171), .B(n_83), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_174), .B(n_147), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_165), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_190), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_183), .A2(n_146), .B1(n_84), .B2(n_99), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_178), .B(n_146), .Y(n_217) );
NOR2xp33_ASAP7_75t_R g218 ( .A(n_156), .B(n_108), .Y(n_218) );
AOI21x1_ASAP7_75t_L g219 ( .A1(n_193), .A2(n_106), .B(n_98), .Y(n_219) );
NAND2x1p5_ASAP7_75t_L g220 ( .A(n_157), .B(n_93), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_175), .B(n_152), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_190), .Y(n_222) );
INVx2_ASAP7_75t_SL g223 ( .A(n_180), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_174), .B(n_102), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_168), .B(n_109), .Y(n_225) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_183), .A2(n_113), .B1(n_109), .B2(n_106), .Y(n_226) );
BUFx3_ASAP7_75t_L g227 ( .A(n_177), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_180), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_174), .B(n_82), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_180), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_177), .Y(n_231) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_171), .Y(n_232) );
NOR2x2_ASAP7_75t_L g233 ( .A(n_164), .B(n_7), .Y(n_233) );
INVx3_ASAP7_75t_L g234 ( .A(n_157), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_165), .Y(n_235) );
OR2x2_ASAP7_75t_L g236 ( .A(n_185), .B(n_7), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_192), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_196), .B(n_180), .Y(n_238) );
AOI22xp5_ASAP7_75t_L g239 ( .A1(n_164), .A2(n_91), .B1(n_88), .B2(n_104), .Y(n_239) );
BUFx2_ASAP7_75t_L g240 ( .A(n_185), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_181), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_196), .B(n_101), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_170), .B(n_88), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_179), .B(n_81), .Y(n_244) );
BUFx8_ASAP7_75t_SL g245 ( .A(n_163), .Y(n_245) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_163), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_196), .B(n_87), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_192), .B(n_87), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_209), .Y(n_249) );
AO22x1_ASAP7_75t_L g250 ( .A1(n_232), .A2(n_166), .B1(n_163), .B2(n_164), .Y(n_250) );
BUFx3_ASAP7_75t_L g251 ( .A(n_245), .Y(n_251) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_231), .Y(n_252) );
INVx3_ASAP7_75t_L g253 ( .A(n_209), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_211), .A2(n_160), .B(n_161), .C(n_172), .Y(n_254) );
INVx1_ASAP7_75t_SL g255 ( .A(n_240), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_238), .A2(n_172), .B(n_160), .Y(n_256) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_231), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_198), .B(n_187), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_213), .A2(n_160), .B(n_161), .Y(n_259) );
BUFx8_ASAP7_75t_L g260 ( .A(n_236), .Y(n_260) );
INVx1_ASAP7_75t_SL g261 ( .A(n_245), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_209), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_200), .Y(n_263) );
INVx2_ASAP7_75t_SL g264 ( .A(n_200), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g265 ( .A(n_218), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_234), .Y(n_266) );
BUFx2_ASAP7_75t_R g267 ( .A(n_236), .Y(n_267) );
AND2x4_ASAP7_75t_L g268 ( .A(n_204), .B(n_168), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_198), .B(n_187), .Y(n_269) );
A2O1A1Ixp33_ASAP7_75t_L g270 ( .A1(n_237), .A2(n_160), .B(n_161), .C(n_195), .Y(n_270) );
AOI21x1_ASAP7_75t_L g271 ( .A1(n_213), .A2(n_195), .B(n_197), .Y(n_271) );
BUFx2_ASAP7_75t_L g272 ( .A(n_218), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_234), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_228), .Y(n_274) );
A2O1A1Ixp33_ASAP7_75t_L g275 ( .A1(n_237), .A2(n_161), .B(n_182), .C(n_186), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_223), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_204), .B(n_166), .Y(n_277) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_223), .B(n_187), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_231), .Y(n_279) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_202), .A2(n_191), .B(n_197), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_204), .B(n_173), .Y(n_281) );
NOR2x1_ASAP7_75t_L g282 ( .A(n_207), .B(n_166), .Y(n_282) );
OR2x2_ASAP7_75t_L g283 ( .A(n_246), .B(n_173), .Y(n_283) );
OAI22xp5_ASAP7_75t_L g284 ( .A1(n_199), .A2(n_197), .B1(n_168), .B2(n_177), .Y(n_284) );
OR2x6_ASAP7_75t_L g285 ( .A(n_201), .B(n_197), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g286 ( .A1(n_217), .A2(n_197), .B(n_181), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_225), .B(n_187), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_230), .Y(n_288) );
NAND3xp33_ASAP7_75t_L g289 ( .A(n_226), .B(n_182), .C(n_186), .Y(n_289) );
AOI22xp33_ASAP7_75t_SL g290 ( .A1(n_225), .A2(n_156), .B1(n_81), .B2(n_101), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_234), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_208), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_203), .B(n_156), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_231), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_292), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_268), .B(n_201), .Y(n_296) );
AO21x1_ASAP7_75t_L g297 ( .A1(n_258), .A2(n_248), .B(n_247), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_252), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_274), .Y(n_299) );
OAI21x1_ASAP7_75t_L g300 ( .A1(n_258), .A2(n_219), .B(n_242), .Y(n_300) );
OAI21x1_ASAP7_75t_L g301 ( .A1(n_269), .A2(n_242), .B(n_220), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_252), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_255), .B(n_201), .Y(n_303) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_285), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_268), .B(n_225), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_288), .Y(n_306) );
AOI22xp5_ASAP7_75t_L g307 ( .A1(n_285), .A2(n_221), .B1(n_216), .B2(n_239), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_252), .Y(n_308) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_252), .Y(n_309) );
OAI21x1_ASAP7_75t_L g310 ( .A1(n_269), .A2(n_220), .B(n_244), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_257), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_285), .B(n_214), .Y(n_312) );
NAND2x1p5_ASAP7_75t_L g313 ( .A(n_257), .B(n_227), .Y(n_313) );
OAI21x1_ASAP7_75t_L g314 ( .A1(n_286), .A2(n_208), .B(n_210), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_270), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_257), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_277), .B(n_214), .Y(n_317) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_257), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g319 ( .A1(n_254), .A2(n_205), .B(n_222), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_279), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_281), .A2(n_206), .B1(n_215), .B2(n_241), .Y(n_321) );
AOI21x1_ASAP7_75t_L g322 ( .A1(n_271), .A2(n_169), .B(n_159), .Y(n_322) );
OA21x2_ASAP7_75t_L g323 ( .A1(n_275), .A2(n_210), .B(n_235), .Y(n_323) );
OAI21x1_ASAP7_75t_SL g324 ( .A1(n_280), .A2(n_284), .B(n_287), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_264), .B(n_235), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_290), .A2(n_227), .B1(n_233), .B2(n_243), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_319), .A2(n_278), .B(n_275), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_326), .A2(n_281), .B1(n_282), .B2(n_260), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_309), .Y(n_329) );
OAI22xp5_ASAP7_75t_SL g330 ( .A1(n_326), .A2(n_265), .B1(n_261), .B2(n_251), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_317), .B(n_263), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_295), .Y(n_332) );
OAI21xp5_ASAP7_75t_L g333 ( .A1(n_307), .A2(n_270), .B(n_289), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_296), .A2(n_260), .B1(n_290), .B2(n_283), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_319), .A2(n_297), .B(n_314), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g336 ( .A1(n_307), .A2(n_250), .B1(n_293), .B2(n_272), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_304), .A2(n_267), .B1(n_276), .B2(n_293), .Y(n_337) );
AO21x2_ASAP7_75t_L g338 ( .A1(n_324), .A2(n_278), .B(n_256), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_303), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_297), .A2(n_259), .B(n_276), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_303), .Y(n_341) );
BUFx4f_ASAP7_75t_SL g342 ( .A(n_325), .Y(n_342) );
BUFx2_ASAP7_75t_L g343 ( .A(n_304), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_314), .A2(n_294), .B(n_279), .Y(n_344) );
A2O1A1Ixp33_ASAP7_75t_L g345 ( .A1(n_315), .A2(n_253), .B(n_291), .C(n_273), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_296), .A2(n_233), .B1(n_253), .B2(n_262), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g347 ( .A1(n_321), .A2(n_229), .B1(n_224), .B2(n_249), .C(n_266), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_324), .A2(n_279), .B1(n_156), .B2(n_101), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_315), .A2(n_279), .B1(n_101), .B2(n_105), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_299), .Y(n_350) );
OR2x6_ASAP7_75t_L g351 ( .A(n_312), .B(n_212), .Y(n_351) );
OAI221xp5_ASAP7_75t_L g352 ( .A1(n_305), .A2(n_101), .B1(n_105), .B2(n_133), .C(n_143), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_305), .B(n_9), .Y(n_353) );
INVxp67_ASAP7_75t_L g354 ( .A(n_332), .Y(n_354) );
OAI221xp5_ASAP7_75t_L g355 ( .A1(n_328), .A2(n_299), .B1(n_306), .B2(n_295), .C(n_312), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_350), .B(n_295), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_333), .B(n_306), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_329), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_339), .B(n_317), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_328), .B(n_314), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_329), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_329), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_331), .B(n_323), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_331), .B(n_323), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_338), .B(n_323), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_341), .B(n_323), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_338), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_345), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_329), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_343), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_340), .Y(n_371) );
INVx5_ASAP7_75t_L g372 ( .A(n_342), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_336), .B(n_327), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_348), .B(n_323), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_348), .B(n_310), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_346), .B(n_325), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_342), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_346), .B(n_325), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_335), .B(n_310), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_334), .B(n_325), .Y(n_380) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_344), .Y(n_381) );
AO21x2_ASAP7_75t_L g382 ( .A1(n_352), .A2(n_322), .B(n_310), .Y(n_382) );
INVx3_ASAP7_75t_L g383 ( .A(n_353), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_370), .B(n_334), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_367), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_367), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_363), .B(n_301), .Y(n_387) );
A2O1A1Ixp33_ASAP7_75t_SL g388 ( .A1(n_371), .A2(n_337), .B(n_349), .C(n_158), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_366), .Y(n_389) );
NOR3xp33_ASAP7_75t_SL g390 ( .A(n_355), .B(n_330), .C(n_347), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_363), .B(n_301), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_355), .A2(n_351), .B1(n_349), .B2(n_301), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_370), .B(n_351), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_354), .Y(n_394) );
OAI221xp5_ASAP7_75t_L g395 ( .A1(n_380), .A2(n_351), .B1(n_101), .B2(n_105), .C(n_313), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_365), .Y(n_396) );
INVx1_ASAP7_75t_SL g397 ( .A(n_370), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_366), .Y(n_398) );
NAND2xp33_ASAP7_75t_R g399 ( .A(n_383), .B(n_9), .Y(n_399) );
INVxp67_ASAP7_75t_SL g400 ( .A(n_383), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_364), .B(n_105), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_359), .B(n_316), .Y(n_402) );
AND2x4_ASAP7_75t_L g403 ( .A(n_360), .B(n_311), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_365), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_357), .Y(n_405) );
OAI33xp33_ASAP7_75t_L g406 ( .A1(n_357), .A2(n_10), .A3(n_11), .B1(n_12), .B2(n_13), .B3(n_16), .Y(n_406) );
NAND3x1_ASAP7_75t_L g407 ( .A(n_364), .B(n_322), .C(n_11), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_365), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_360), .B(n_105), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_356), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_360), .B(n_105), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_359), .B(n_320), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_371), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_380), .A2(n_320), .B1(n_298), .B2(n_316), .Y(n_414) );
INVx3_ASAP7_75t_L g415 ( .A(n_358), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_356), .B(n_320), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_379), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_354), .B(n_298), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_376), .B(n_298), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_383), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_381), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_383), .B(n_313), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_376), .B(n_316), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_378), .A2(n_311), .B1(n_308), .B2(n_302), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_379), .Y(n_425) );
INVx1_ASAP7_75t_SL g426 ( .A(n_394), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_396), .B(n_373), .Y(n_427) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_401), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_396), .B(n_381), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_410), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_385), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_396), .B(n_373), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_401), .Y(n_433) );
INVx4_ASAP7_75t_L g434 ( .A(n_422), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_404), .B(n_374), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_410), .B(n_378), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_393), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_404), .B(n_374), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_404), .B(n_375), .Y(n_439) );
INVx2_ASAP7_75t_SL g440 ( .A(n_397), .Y(n_440) );
INVx3_ASAP7_75t_L g441 ( .A(n_421), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_399), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_390), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_385), .Y(n_444) );
OAI221xp5_ASAP7_75t_L g445 ( .A1(n_392), .A2(n_377), .B1(n_368), .B2(n_375), .C(n_372), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_408), .B(n_361), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_386), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_408), .B(n_361), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_389), .B(n_377), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_386), .Y(n_450) );
AOI21xp33_ASAP7_75t_L g451 ( .A1(n_393), .A2(n_377), .B(n_368), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_389), .B(n_358), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_408), .B(n_358), .Y(n_453) );
INVxp67_ASAP7_75t_L g454 ( .A(n_420), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_409), .B(n_369), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_384), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_395), .A2(n_372), .B1(n_382), .B2(n_369), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_398), .B(n_369), .Y(n_458) );
NOR3xp33_ASAP7_75t_SL g459 ( .A(n_406), .B(n_372), .C(n_13), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_384), .Y(n_460) );
INVx1_ASAP7_75t_SL g461 ( .A(n_397), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_409), .B(n_362), .Y(n_462) );
NAND3xp33_ASAP7_75t_L g463 ( .A(n_411), .B(n_133), .C(n_143), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_411), .B(n_362), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_413), .Y(n_465) );
NAND4xp25_ASAP7_75t_L g466 ( .A(n_424), .B(n_361), .C(n_362), .D(n_17), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_402), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_398), .B(n_382), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_387), .B(n_391), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_400), .A2(n_372), .B1(n_382), .B2(n_311), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_405), .B(n_372), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_387), .B(n_382), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_412), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_405), .B(n_372), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_391), .B(n_148), .Y(n_475) );
AND2x4_ASAP7_75t_L g476 ( .A(n_403), .B(n_372), .Y(n_476) );
INVx2_ASAP7_75t_SL g477 ( .A(n_422), .Y(n_477) );
NOR2xp33_ASAP7_75t_R g478 ( .A(n_416), .B(n_10), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_423), .B(n_133), .Y(n_479) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_418), .Y(n_480) );
AND2x2_ASAP7_75t_SL g481 ( .A(n_421), .B(n_318), .Y(n_481) );
INVxp67_ASAP7_75t_L g482 ( .A(n_468), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_444), .Y(n_483) );
OR2x6_ASAP7_75t_L g484 ( .A(n_434), .B(n_421), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_426), .B(n_425), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_480), .B(n_419), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_444), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_456), .B(n_423), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_431), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_460), .B(n_425), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_431), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_447), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_465), .Y(n_493) );
AND3x2_ASAP7_75t_L g494 ( .A(n_428), .B(n_418), .C(n_417), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_447), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_469), .B(n_403), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_469), .B(n_403), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_467), .B(n_417), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_465), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_434), .B(n_403), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_434), .B(n_413), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_473), .B(n_413), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_433), .B(n_415), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_461), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_477), .B(n_415), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_430), .B(n_414), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_450), .Y(n_507) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_459), .A2(n_407), .B(n_388), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_472), .B(n_415), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_443), .A2(n_415), .B1(n_308), .B2(n_302), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_477), .B(n_16), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_437), .B(n_407), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_450), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_436), .B(n_133), .Y(n_514) );
NAND2x1_ASAP7_75t_L g515 ( .A(n_476), .B(n_318), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_449), .Y(n_516) );
INVx2_ASAP7_75t_SL g517 ( .A(n_440), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_452), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_427), .B(n_143), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_458), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_429), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_427), .B(n_435), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_432), .B(n_143), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_432), .B(n_143), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_466), .A2(n_300), .B(n_308), .C(n_302), .Y(n_525) );
AND2x2_ASAP7_75t_SL g526 ( .A(n_481), .B(n_318), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_472), .B(n_148), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_443), .A2(n_313), .B1(n_300), .B2(n_148), .Y(n_528) );
OAI21xp5_ASAP7_75t_SL g529 ( .A1(n_476), .A2(n_313), .B(n_148), .Y(n_529) );
BUFx4_ASAP7_75t_SL g530 ( .A(n_442), .Y(n_530) );
NAND4xp25_ASAP7_75t_L g531 ( .A(n_457), .B(n_188), .C(n_176), .D(n_169), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_455), .B(n_148), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_458), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_429), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_435), .B(n_318), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_438), .B(n_318), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_441), .Y(n_537) );
NOR4xp25_ASAP7_75t_L g538 ( .A(n_525), .B(n_445), .C(n_471), .D(n_474), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_516), .B(n_468), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_518), .B(n_475), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_485), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_530), .Y(n_542) );
OAI22xp33_ASAP7_75t_L g543 ( .A1(n_484), .A2(n_442), .B1(n_470), .B2(n_463), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_512), .A2(n_475), .B1(n_439), .B2(n_454), .Y(n_544) );
NAND3xp33_ASAP7_75t_SL g545 ( .A(n_529), .B(n_478), .C(n_479), .Y(n_545) );
AND2x4_ASAP7_75t_SL g546 ( .A(n_484), .B(n_476), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_530), .Y(n_547) );
INVx1_ASAP7_75t_SL g548 ( .A(n_504), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_522), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_483), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_487), .Y(n_551) );
OA21x2_ASAP7_75t_SL g552 ( .A1(n_494), .A2(n_481), .B(n_451), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_492), .Y(n_553) );
O2A1O1Ixp33_ASAP7_75t_L g554 ( .A1(n_508), .A2(n_479), .B(n_440), .C(n_441), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_495), .Y(n_555) );
OAI221xp5_ASAP7_75t_L g556 ( .A1(n_525), .A2(n_438), .B1(n_441), .B2(n_446), .C(n_453), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_484), .A2(n_439), .B1(n_462), .B2(n_455), .Y(n_557) );
AOI31xp33_ASAP7_75t_L g558 ( .A1(n_511), .A2(n_464), .A3(n_462), .B(n_453), .Y(n_558) );
OAI21xp5_ASAP7_75t_SL g559 ( .A1(n_494), .A2(n_464), .B(n_448), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_482), .B(n_448), .Y(n_560) );
NAND3xp33_ASAP7_75t_L g561 ( .A(n_504), .B(n_527), .C(n_514), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_482), .B(n_446), .Y(n_562) );
OAI21xp33_ASAP7_75t_SL g563 ( .A1(n_526), .A2(n_300), .B(n_19), .Y(n_563) );
OAI32xp33_ASAP7_75t_L g564 ( .A1(n_501), .A2(n_188), .A3(n_176), .B1(n_169), .B2(n_167), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_507), .Y(n_565) );
NOR2xp33_ASAP7_75t_SL g566 ( .A(n_526), .B(n_318), .Y(n_566) );
OAI221xp5_ASAP7_75t_L g567 ( .A1(n_506), .A2(n_188), .B1(n_176), .B2(n_167), .C(n_159), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_520), .B(n_318), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_500), .A2(n_515), .B1(n_510), .B2(n_486), .Y(n_569) );
NOR4xp25_ASAP7_75t_L g570 ( .A(n_527), .B(n_167), .C(n_159), .D(n_158), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_531), .A2(n_309), .B(n_158), .Y(n_571) );
A2O1A1Ixp33_ASAP7_75t_L g572 ( .A1(n_517), .A2(n_309), .B(n_22), .C(n_23), .Y(n_572) );
AOI222xp33_ASAP7_75t_L g573 ( .A1(n_533), .A2(n_309), .B1(n_24), .B2(n_26), .C1(n_29), .C2(n_31), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_490), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_503), .A2(n_309), .B1(n_38), .B2(n_41), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_509), .A2(n_309), .B1(n_48), .B2(n_49), .Y(n_576) );
NAND3xp33_ASAP7_75t_L g577 ( .A(n_517), .B(n_309), .C(n_50), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_497), .B(n_18), .Y(n_578) );
INVx1_ASAP7_75t_SL g579 ( .A(n_542), .Y(n_579) );
OAI22xp33_ASAP7_75t_SL g580 ( .A1(n_569), .A2(n_498), .B1(n_502), .B2(n_519), .Y(n_580) );
INVx1_ASAP7_75t_SL g581 ( .A(n_547), .Y(n_581) );
O2A1O1Ixp5_ASAP7_75t_SL g582 ( .A1(n_541), .A2(n_523), .B(n_524), .C(n_532), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_548), .B(n_534), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_550), .Y(n_584) );
O2A1O1Ixp33_ASAP7_75t_L g585 ( .A1(n_543), .A2(n_537), .B(n_513), .C(n_497), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_574), .B(n_549), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_544), .B(n_496), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_551), .Y(n_588) );
CKINVDCx14_ASAP7_75t_R g589 ( .A(n_545), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_562), .Y(n_590) );
OAI22xp33_ASAP7_75t_L g591 ( .A1(n_559), .A2(n_521), .B1(n_534), .B2(n_528), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_553), .Y(n_592) );
INVxp67_ASAP7_75t_L g593 ( .A(n_561), .Y(n_593) );
AOI222xp33_ASAP7_75t_L g594 ( .A1(n_559), .A2(n_509), .B1(n_521), .B2(n_505), .C1(n_513), .C2(n_489), .Y(n_594) );
INVxp67_ASAP7_75t_L g595 ( .A(n_558), .Y(n_595) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_554), .B(n_537), .Y(n_596) );
NAND3xp33_ASAP7_75t_L g597 ( .A(n_563), .B(n_510), .C(n_489), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_555), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_565), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_560), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_539), .Y(n_601) );
NOR2x1_ASAP7_75t_L g602 ( .A(n_577), .B(n_491), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_568), .Y(n_603) );
AOI322xp5_ASAP7_75t_L g604 ( .A1(n_589), .A2(n_557), .A3(n_552), .B1(n_540), .B2(n_578), .C1(n_566), .C2(n_491), .Y(n_604) );
OAI21xp33_ASAP7_75t_L g605 ( .A1(n_589), .A2(n_538), .B(n_556), .Y(n_605) );
AOI311xp33_ASAP7_75t_L g606 ( .A1(n_580), .A2(n_567), .A3(n_572), .B(n_571), .C(n_546), .Y(n_606) );
INVxp67_ASAP7_75t_L g607 ( .A(n_579), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_593), .B(n_493), .Y(n_608) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_584), .Y(n_609) );
OAI21xp33_ASAP7_75t_L g610 ( .A1(n_595), .A2(n_573), .B(n_570), .Y(n_610) );
INVx2_ASAP7_75t_SL g611 ( .A(n_581), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_590), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_584), .Y(n_613) );
INVxp67_ASAP7_75t_L g614 ( .A(n_588), .Y(n_614) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_591), .A2(n_585), .B(n_596), .Y(n_615) );
AOI22xp33_ASAP7_75t_SL g616 ( .A1(n_597), .A2(n_488), .B1(n_493), .B2(n_499), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_L g617 ( .A1(n_596), .A2(n_570), .B(n_564), .C(n_499), .Y(n_617) );
AO21x1_ASAP7_75t_L g618 ( .A1(n_586), .A2(n_575), .B(n_576), .Y(n_618) );
OAI21xp5_ASAP7_75t_L g619 ( .A1(n_615), .A2(n_602), .B(n_594), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_605), .A2(n_601), .B1(n_592), .B2(n_599), .C(n_598), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_616), .A2(n_587), .B1(n_600), .B2(n_583), .Y(n_621) );
OA22x2_ASAP7_75t_L g622 ( .A1(n_611), .A2(n_587), .B1(n_600), .B2(n_603), .Y(n_622) );
INVx1_ASAP7_75t_SL g623 ( .A(n_612), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_607), .B(n_603), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_610), .A2(n_536), .B1(n_535), .B2(n_582), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_618), .A2(n_582), .B1(n_53), .B2(n_57), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_617), .A2(n_52), .B(n_59), .Y(n_627) );
NAND4xp75_ASAP7_75t_L g628 ( .A(n_619), .B(n_606), .C(n_608), .D(n_604), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_623), .B(n_608), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_625), .B(n_614), .Y(n_630) );
NOR2xp33_ASAP7_75t_R g631 ( .A(n_624), .B(n_626), .Y(n_631) );
NAND3xp33_ASAP7_75t_SL g632 ( .A(n_620), .B(n_609), .C(n_613), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_629), .Y(n_633) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_630), .Y(n_634) );
OAI31xp33_ASAP7_75t_L g635 ( .A1(n_628), .A2(n_621), .A3(n_627), .B(n_622), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_633), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_633), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_636), .Y(n_638) );
OAI321xp33_ASAP7_75t_L g639 ( .A1(n_638), .A2(n_637), .A3(n_636), .B1(n_632), .B2(n_635), .C(n_634), .Y(n_639) );
OAI33xp33_ASAP7_75t_R g640 ( .A1(n_639), .A2(n_631), .A3(n_62), .B1(n_63), .B2(n_67), .B3(n_61), .Y(n_640) );
OA21x2_ASAP7_75t_L g641 ( .A1(n_640), .A2(n_68), .B(n_70), .Y(n_641) );
AOI21xp5_ASAP7_75t_L g642 ( .A1(n_641), .A2(n_71), .B(n_74), .Y(n_642) );
endmodule