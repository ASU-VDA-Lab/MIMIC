module fake_jpeg_10533_n_283 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_283);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_283;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_30),
.B1(n_19),
.B2(n_33),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_44),
.A2(n_51),
.B(n_16),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_46),
.B(n_49),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

NAND3xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_12),
.C(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_31),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_30),
.B1(n_19),
.B2(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_30),
.B1(n_26),
.B2(n_24),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_54),
.A2(n_57),
.B1(n_59),
.B2(n_16),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_30),
.B1(n_33),
.B2(n_22),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_36),
.A2(n_33),
.B1(n_22),
.B2(n_23),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_37),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_64),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_72),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_70),
.B(n_77),
.Y(n_112)
);

AO22x1_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_54),
.B1(n_57),
.B2(n_66),
.Y(n_71)
);

AND2x4_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_89),
.Y(n_110)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_19),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_59),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_56),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_16),
.B1(n_61),
.B2(n_20),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_27),
.C(n_22),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_29),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_58),
.A2(n_26),
.B1(n_24),
.B2(n_20),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_84),
.Y(n_109)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_26),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_52),
.Y(n_113)
);

AND2x4_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_29),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_R g104 ( 
.A(n_89),
.B(n_52),
.Y(n_104)
);

OAI22x1_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_27),
.B1(n_17),
.B2(n_31),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_93),
.B(n_94),
.Y(n_139)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_98),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_61),
.B1(n_58),
.B2(n_50),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_99),
.B1(n_113),
.B2(n_82),
.Y(n_117)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_45),
.Y(n_131)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

AOI32xp33_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_71),
.A3(n_88),
.B1(n_79),
.B2(n_70),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_103),
.A2(n_104),
.B(n_110),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_86),
.B(n_24),
.Y(n_129)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_29),
.Y(n_140)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_108),
.A2(n_111),
.B1(n_84),
.B2(n_83),
.Y(n_141)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_71),
.A2(n_73),
.B1(n_77),
.B2(n_89),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_114),
.A2(n_78),
.B1(n_67),
.B2(n_27),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_117),
.B(n_119),
.Y(n_168)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

AOI22x1_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_52),
.B1(n_64),
.B2(n_62),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_126),
.B1(n_134),
.B2(n_137),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_86),
.C(n_73),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_130),
.C(n_115),
.Y(n_147)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_125),
.Y(n_164)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

AOI22x1_ASAP7_75t_L g126 ( 
.A1(n_110),
.A2(n_64),
.B1(n_68),
.B2(n_47),
.Y(n_126)
);

NOR2xp67_ASAP7_75t_SL g127 ( 
.A(n_110),
.B(n_87),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_127),
.A2(n_104),
.B(n_114),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_129),
.A2(n_135),
.B1(n_141),
.B2(n_105),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_68),
.C(n_75),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_132),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_92),
.B(n_25),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_94),
.A2(n_97),
.B1(n_99),
.B2(n_101),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_92),
.B(n_93),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_138),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_97),
.A2(n_67),
.B1(n_78),
.B2(n_47),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_25),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_31),
.Y(n_159)
);

INVxp33_ASAP7_75t_SL g142 ( 
.A(n_126),
.Y(n_142)
);

INVxp67_ASAP7_75t_SL g177 ( 
.A(n_142),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_143),
.B(n_146),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_144),
.B(n_17),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_126),
.B1(n_120),
.B2(n_139),
.Y(n_145)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_118),
.C(n_133),
.Y(n_171)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_150),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_120),
.A2(n_108),
.B1(n_102),
.B2(n_106),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_149),
.A2(n_153),
.B1(n_161),
.B2(n_28),
.Y(n_175)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

OR2x2_ASAP7_75t_SL g151 ( 
.A(n_127),
.B(n_29),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_151),
.A2(n_154),
.B(n_159),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_131),
.A2(n_65),
.B1(n_53),
.B2(n_21),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_130),
.B(n_136),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_138),
.Y(n_157)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_0),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_158),
.A2(n_167),
.B(n_1),
.Y(n_186)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_160),
.A2(n_165),
.B(n_1),
.Y(n_191)
);

AO22x2_ASAP7_75t_L g161 ( 
.A1(n_134),
.A2(n_53),
.B1(n_29),
.B2(n_75),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_122),
.A2(n_123),
.B1(n_119),
.B2(n_125),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_162),
.A2(n_166),
.B1(n_28),
.B2(n_23),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_95),
.Y(n_163)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_163),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_123),
.A2(n_28),
.B1(n_23),
.B2(n_21),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_124),
.B(n_0),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_17),
.Y(n_169)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_169),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_180),
.C(n_183),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_159),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_181),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_175),
.A2(n_187),
.B1(n_184),
.B2(n_161),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_152),
.A2(n_21),
.B1(n_18),
.B2(n_91),
.Y(n_176)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_152),
.A2(n_18),
.B1(n_116),
.B2(n_31),
.Y(n_178)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_116),
.Y(n_180)
);

NAND3xp33_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_9),
.C(n_15),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_116),
.C(n_18),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_160),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_184),
.A2(n_186),
.B(n_151),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_8),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_188),
.C(n_156),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_149),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_169),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

AO21x1_ASAP7_75t_L g204 ( 
.A1(n_191),
.A2(n_161),
.B(n_166),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_192),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_197),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_196),
.B(n_204),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_191),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_199),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_189),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_193),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_203),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_201),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_178),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_215),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_174),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_214),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_170),
.A2(n_168),
.B1(n_156),
.B2(n_161),
.Y(n_208)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_172),
.A2(n_175),
.B1(n_187),
.B2(n_177),
.Y(n_209)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_209),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_171),
.B(n_155),
.C(n_150),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_212),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_155),
.C(n_146),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_176),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_189),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_202),
.A2(n_172),
.B1(n_182),
.B2(n_179),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_218),
.A2(n_214),
.B1(n_195),
.B2(n_182),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_185),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_224),
.C(n_227),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_183),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_186),
.Y(n_227)
);

XNOR2x1_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_158),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_198),
.Y(n_238)
);

AOI21xp33_ASAP7_75t_L g229 ( 
.A1(n_211),
.A2(n_158),
.B(n_167),
.Y(n_229)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_229),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_209),
.Y(n_232)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_232),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_223),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_237),
.Y(n_251)
);

INVxp67_ASAP7_75t_SL g235 ( 
.A(n_231),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_213),
.Y(n_248)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_218),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_236),
.A2(n_239),
.B(n_196),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_194),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_219),
.Y(n_249)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

O2A1O1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_226),
.A2(n_208),
.B(n_201),
.C(n_202),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_241),
.A2(n_242),
.B1(n_220),
.B2(n_228),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_210),
.C(n_212),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_245),
.C(n_224),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_206),
.C(n_213),
.Y(n_245)
);

OAI321xp33_ASAP7_75t_L g246 ( 
.A1(n_241),
.A2(n_204),
.A3(n_195),
.B1(n_161),
.B2(n_216),
.C(n_211),
.Y(n_246)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_246),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_238),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_252),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_219),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_255),
.C(n_256),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_148),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_254),
.Y(n_259)
);

NAND4xp25_ASAP7_75t_SL g254 ( 
.A(n_244),
.B(n_165),
.C(n_167),
.D(n_153),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_239),
.B(n_242),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_234),
.B1(n_245),
.B2(n_240),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_243),
.C(n_240),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_263),
.C(n_264),
.Y(n_267)
);

NOR2xp67_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_227),
.Y(n_262)
);

AOI31xp33_ASAP7_75t_L g266 ( 
.A1(n_262),
.A2(n_247),
.A3(n_251),
.B(n_222),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_221),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_265),
.B(n_11),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_268),
.Y(n_273)
);

OAI221xp5_ASAP7_75t_L g268 ( 
.A1(n_257),
.A2(n_221),
.B1(n_9),
.B2(n_10),
.C(n_15),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_259),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_271),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_258),
.A2(n_14),
.B(n_12),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_270),
.A2(n_272),
.B(n_11),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_260),
.A2(n_11),
.B(n_10),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_274),
.A2(n_275),
.B(n_277),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_264),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_272),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_273),
.A2(n_263),
.B(n_265),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_276),
.Y(n_280)
);

AOI322xp5_ASAP7_75t_L g281 ( 
.A1(n_280),
.A2(n_278),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_281)
);

OAI321xp33_ASAP7_75t_L g282 ( 
.A1(n_281),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_3),
.Y(n_283)
);


endmodule