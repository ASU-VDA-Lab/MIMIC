module fake_jpeg_6581_n_335 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_3),
.B(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_37),
.Y(n_47)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_15),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_41),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_41),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_45),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_19),
.B1(n_24),
.B2(n_23),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_46),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_16),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_51),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_23),
.B1(n_24),
.B2(n_19),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_54),
.A2(n_60),
.B1(n_22),
.B2(n_21),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_19),
.B1(n_23),
.B2(n_24),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_16),
.B1(n_20),
.B2(n_21),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_35),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_57),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_38),
.A2(n_23),
.B1(n_24),
.B2(n_28),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_61),
.Y(n_74)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_64),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_20),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_69),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_78),
.Y(n_106)
);

AO22x1_ASAP7_75t_SL g73 ( 
.A1(n_46),
.A2(n_38),
.B1(n_42),
.B2(n_33),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_73),
.A2(n_82),
.B1(n_55),
.B2(n_50),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_75),
.A2(n_87),
.B1(n_28),
.B2(n_29),
.Y(n_95)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_11),
.B(n_13),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_65),
.B(n_64),
.Y(n_111)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_83),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_16),
.B1(n_31),
.B2(n_17),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_85),
.A2(n_91),
.B1(n_93),
.B2(n_50),
.Y(n_101)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_90),
.Y(n_114)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_57),
.A2(n_28),
.B1(n_22),
.B2(n_21),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_95),
.B(n_113),
.Y(n_123)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_98),
.Y(n_120)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_102),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_SL g100 ( 
.A1(n_94),
.A2(n_49),
.B(n_51),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_100),
.A2(n_112),
.B1(n_72),
.B2(n_90),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_101),
.A2(n_111),
.B1(n_22),
.B2(n_62),
.Y(n_146)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_109),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_48),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_105),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_84),
.B(n_48),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_73),
.A2(n_63),
.B1(n_50),
.B2(n_55),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_110),
.B1(n_118),
.B2(n_62),
.Y(n_129)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

FAx1_ASAP7_75t_SL g113 ( 
.A(n_84),
.B(n_70),
.CI(n_47),
.CON(n_113),
.SN(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_115),
.B(n_116),
.Y(n_147)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_71),
.A2(n_31),
.B(n_17),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_29),
.B(n_27),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_73),
.A2(n_55),
.B1(n_58),
.B2(n_69),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_47),
.Y(n_119)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_77),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_121),
.B(n_131),
.C(n_143),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_116),
.A2(n_73),
.B1(n_71),
.B2(n_86),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_122),
.A2(n_146),
.B1(n_107),
.B2(n_113),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_114),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_134),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_129),
.A2(n_62),
.B1(n_91),
.B2(n_83),
.Y(n_170)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_133),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_77),
.C(n_58),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_132),
.B(n_135),
.Y(n_148)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_139),
.Y(n_160)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_138),
.Y(n_174)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_141),
.A2(n_111),
.B(n_123),
.Y(n_152)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_145),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_58),
.C(n_89),
.Y(n_143)
);

A2O1A1O1Ixp25_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_90),
.B(n_67),
.C(n_74),
.D(n_30),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_144),
.B(n_74),
.Y(n_169)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_97),
.Y(n_145)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_153),
.Y(n_194)
);

FAx1_ASAP7_75t_SL g180 ( 
.A(n_152),
.B(n_175),
.CI(n_141),
.CON(n_180),
.SN(n_180)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_118),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_154),
.A2(n_162),
.B1(n_170),
.B2(n_132),
.Y(n_189)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_156),
.B(n_163),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_103),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_159),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_122),
.B(n_102),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_142),
.B(n_109),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_167),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_115),
.B1(n_98),
.B2(n_110),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_165),
.Y(n_176)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_92),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_131),
.C(n_144),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_166),
.C(n_152),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_169),
.B(n_157),
.Y(n_186)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_151),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_89),
.Y(n_173)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_173),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_SL g175 ( 
.A1(n_126),
.A2(n_25),
.B(n_26),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_174),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_182),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_185),
.C(n_188),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_180),
.B(n_181),
.Y(n_221)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_149),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_200),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_165),
.C(n_168),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_155),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_135),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_189),
.A2(n_193),
.B1(n_195),
.B2(n_156),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_139),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_192),
.C(n_198),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_137),
.C(n_134),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_162),
.A2(n_89),
.B1(n_80),
.B2(n_78),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_154),
.A2(n_133),
.B1(n_130),
.B2(n_17),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_167),
.B(n_67),
.Y(n_196)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_173),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_197),
.B(n_199),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_67),
.Y(n_198)
);

FAx1_ASAP7_75t_SL g199 ( 
.A(n_172),
.B(n_67),
.CI(n_34),
.CON(n_199),
.SN(n_199)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_153),
.B(n_27),
.Y(n_200)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_201),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_42),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_203),
.C(n_170),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_136),
.C(n_42),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_193),
.A2(n_158),
.B1(n_163),
.B2(n_150),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_204),
.A2(n_224),
.B1(n_25),
.B2(n_26),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_203),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_206),
.A2(n_218),
.B1(n_226),
.B2(n_229),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_148),
.Y(n_208)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_208),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_176),
.A2(n_148),
.B(n_155),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_211),
.A2(n_228),
.B1(n_179),
.B2(n_29),
.Y(n_244)
);

FAx1_ASAP7_75t_SL g251 ( 
.A(n_213),
.B(n_227),
.CI(n_30),
.CON(n_251),
.SN(n_251)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_187),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_216),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_215),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_199),
.Y(n_245)
);

NAND2x1_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_160),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_219),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_190),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_222),
.Y(n_241)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_184),
.A2(n_171),
.B(n_151),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_227),
.Y(n_237)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_184),
.B(n_174),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_195),
.A2(n_17),
.B1(n_31),
.B2(n_26),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_177),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_185),
.C(n_178),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_232),
.C(n_240),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_191),
.C(n_186),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_218),
.B(n_188),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_237),
.Y(n_261)
);

OA21x2_ASAP7_75t_L g234 ( 
.A1(n_216),
.A2(n_199),
.B(n_180),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_234),
.A2(n_210),
.B(n_27),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_223),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_212),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_218),
.C(n_209),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_198),
.C(n_202),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_242),
.B(n_245),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_180),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_243),
.B(n_246),
.Y(n_263)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_136),
.C(n_68),
.Y(n_246)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_247),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_136),
.C(n_68),
.Y(n_248)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_248),
.Y(n_257)
);

AOI21xp33_ASAP7_75t_L g249 ( 
.A1(n_211),
.A2(n_30),
.B(n_25),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_249),
.A2(n_220),
.B(n_228),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_88),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_208),
.Y(n_252)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_252),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_238),
.A2(n_224),
.B1(n_214),
.B2(n_213),
.Y(n_253)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_254),
.A2(n_258),
.B(n_260),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_235),
.A2(n_212),
.B1(n_229),
.B2(n_219),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_267),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_230),
.A2(n_31),
.B(n_1),
.Y(n_264)
);

NOR3xp33_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_0),
.C(n_1),
.Y(n_279)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_269),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_239),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_250),
.A2(n_30),
.B1(n_53),
.B2(n_2),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_270),
.A2(n_242),
.B1(n_14),
.B2(n_13),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_241),
.B(n_252),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_271),
.Y(n_276)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_236),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_257),
.Y(n_282)
);

OAI321xp33_ASAP7_75t_L g273 ( 
.A1(n_259),
.A2(n_234),
.A3(n_251),
.B1(n_245),
.B2(n_243),
.C(n_233),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_273),
.A2(n_278),
.B(n_288),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_232),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_266),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_254),
.B(n_248),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_277),
.A2(n_281),
.B(n_263),
.Y(n_292)
);

OAI321xp33_ASAP7_75t_L g278 ( 
.A1(n_260),
.A2(n_268),
.A3(n_255),
.B1(n_264),
.B2(n_234),
.C(n_253),
.Y(n_278)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_257),
.B(n_240),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_289),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_53),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_283),
.B(n_2),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_284),
.A2(n_267),
.B1(n_262),
.B2(n_265),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_231),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_266),
.C(n_256),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_262),
.B(n_14),
.Y(n_288)
);

FAx1_ASAP7_75t_L g289 ( 
.A(n_261),
.B(n_30),
.CI(n_1),
.CON(n_289),
.SN(n_289)
);

AOI31xp33_ASAP7_75t_L g291 ( 
.A1(n_289),
.A2(n_286),
.A3(n_285),
.B(n_276),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_291),
.A2(n_292),
.B(n_298),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_289),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_294),
.B(n_296),
.Y(n_314)
);

BUFx24_ASAP7_75t_SL g297 ( 
.A(n_274),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_297),
.B(n_299),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_272),
.Y(n_298)
);

BUFx24_ASAP7_75t_SL g299 ( 
.A(n_285),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_0),
.C(n_2),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_300),
.A2(n_303),
.B(n_3),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_280),
.A2(n_13),
.B1(n_11),
.B2(n_3),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_302),
.B(n_304),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_0),
.Y(n_303)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_305),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_307),
.B(n_312),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_290),
.B(n_10),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_311),
.C(n_313),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_301),
.A2(n_4),
.B(n_5),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_4),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_5),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_296),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_315),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_5),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_317),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_5),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_6),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_10),
.Y(n_328)
);

O2A1O1Ixp33_ASAP7_75t_SL g327 ( 
.A1(n_320),
.A2(n_322),
.B(n_318),
.C(n_9),
.Y(n_327)
);

A2O1A1Ixp33_ASAP7_75t_SL g322 ( 
.A1(n_306),
.A2(n_6),
.B(n_7),
.C(n_9),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_310),
.Y(n_325)
);

NAND2xp33_ASAP7_75t_SL g332 ( 
.A(n_325),
.B(n_326),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_308),
.Y(n_326)
);

NAND3xp33_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_329),
.C(n_10),
.Y(n_331)
);

INVxp33_ASAP7_75t_L g330 ( 
.A(n_328),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_322),
.A2(n_6),
.B(n_9),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_331),
.B(n_324),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_330),
.C(n_332),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_322),
.Y(n_335)
);


endmodule