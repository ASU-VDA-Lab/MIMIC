module fake_jpeg_23851_n_242 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_242);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_242;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_12),
.B(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_42),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_39),
.B(n_43),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_1),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_24),
.B(n_1),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_16),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_61),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_43),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_52),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_27),
.B1(n_20),
.B2(n_33),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_53),
.A2(n_63),
.B1(n_18),
.B2(n_75),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_27),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_54),
.B(n_80),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_56),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_27),
.B1(n_16),
.B2(n_20),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_38),
.A2(n_29),
.B1(n_34),
.B2(n_26),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_60),
.A2(n_76),
.B1(n_18),
.B2(n_55),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_22),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_35),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_67),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_19),
.B1(n_25),
.B2(n_33),
.Y(n_63)
);

NOR2x1_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_29),
.Y(n_65)
);

NOR2x1_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_26),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_35),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_31),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_79),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_70),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_37),
.B(n_34),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_30),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_77),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_41),
.A2(n_31),
.B1(n_19),
.B2(n_25),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_40),
.B(n_30),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_28),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g81 ( 
.A1(n_44),
.A2(n_1),
.B(n_2),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_3),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_84),
.A2(n_97),
.B1(n_98),
.B2(n_102),
.Y(n_136)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_89),
.Y(n_114)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_65),
.B(n_44),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_66),
.C(n_64),
.Y(n_135)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_103),
.Y(n_119)
);

OAI32xp33_ASAP7_75t_L g95 ( 
.A1(n_65),
.A2(n_48),
.A3(n_46),
.B1(n_28),
.B2(n_17),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_63),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_48),
.B1(n_46),
.B2(n_28),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_96),
.A2(n_72),
.B1(n_49),
.B2(n_61),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_2),
.Y(n_101)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_57),
.A2(n_48),
.B1(n_28),
.B2(n_5),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_52),
.A2(n_60),
.B1(n_51),
.B2(n_53),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_104),
.A2(n_62),
.B1(n_79),
.B2(n_58),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_59),
.B(n_3),
.Y(n_105)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_110),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_107),
.A2(n_83),
.B(n_84),
.Y(n_123)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_112),
.A2(n_120),
.B1(n_108),
.B2(n_111),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_54),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_113),
.B(n_116),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_56),
.Y(n_115)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_50),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_134),
.B1(n_135),
.B2(n_138),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_121),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_78),
.Y(n_122)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_125),
.C(n_127),
.Y(n_158)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_131),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_50),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_78),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_129),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_83),
.B(n_64),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_91),
.B(n_67),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_72),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_132),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_91),
.B(n_64),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_86),
.B(n_75),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_100),
.A2(n_72),
.B1(n_82),
.B2(n_75),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_107),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_100),
.A2(n_82),
.B1(n_69),
.B2(n_74),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_93),
.B(n_69),
.C(n_74),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_106),
.B(n_103),
.Y(n_162)
);

AOI22x1_ASAP7_75t_SL g142 ( 
.A1(n_112),
.A2(n_130),
.B1(n_136),
.B2(n_95),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_143),
.B(n_144),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_145),
.A2(n_149),
.B1(n_163),
.B2(n_118),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_116),
.A2(n_111),
.B(n_108),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_125),
.B(n_127),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_121),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_152),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_137),
.A2(n_96),
.B1(n_110),
.B2(n_85),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_151),
.B(n_154),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_121),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_99),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_133),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_155),
.B(n_157),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_92),
.Y(n_157)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_139),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_113),
.A2(n_69),
.B1(n_94),
.B2(n_14),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_117),
.B(n_4),
.Y(n_164)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_174),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_173),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_132),
.Y(n_170)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_131),
.Y(n_171)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_141),
.A2(n_130),
.B(n_126),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_140),
.B(n_122),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_179),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_135),
.B1(n_138),
.B2(n_134),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_178),
.A2(n_182),
.B1(n_158),
.B2(n_146),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_183),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_142),
.A2(n_146),
.B1(n_141),
.B2(n_163),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_158),
.A2(n_143),
.B(n_160),
.Y(n_183)
);

NAND3xp33_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_150),
.C(n_160),
.Y(n_184)
);

AOI21xp33_ASAP7_75t_L g201 ( 
.A1(n_184),
.A2(n_154),
.B(n_157),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_186),
.B(n_182),
.Y(n_199)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_192),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_175),
.A2(n_140),
.B1(n_150),
.B2(n_115),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_195),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_179),
.A2(n_155),
.B1(n_149),
.B2(n_129),
.Y(n_191)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_172),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_170),
.Y(n_198)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_198),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_178),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_177),
.C(n_186),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_202),
.C(n_207),
.Y(n_213)
);

NAND4xp25_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_190),
.C(n_180),
.D(n_191),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_183),
.C(n_167),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_166),
.C(n_173),
.Y(n_207)
);

XNOR2x1_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_175),
.Y(n_209)
);

XNOR2x1_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_189),
.Y(n_214)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_193),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_194),
.C(n_123),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_216),
.C(n_217),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_214),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_215),
.B(n_203),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_193),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_204),
.A2(n_197),
.B1(n_196),
.B2(n_165),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_218),
.A2(n_205),
.B1(n_206),
.B2(n_199),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_181),
.C(n_196),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_220),
.C(n_208),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_117),
.C(n_176),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_156),
.C(n_7),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_223),
.B(n_224),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_152),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_226),
.A2(n_176),
.B(n_148),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_217),
.C(n_214),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_213),
.C(n_164),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_229),
.C(n_231),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_156),
.C(n_161),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_6),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_233),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_230),
.A2(n_226),
.B(n_225),
.Y(n_234)
);

NOR3xp33_ASAP7_75t_SL g237 ( 
.A(n_234),
.B(n_236),
.C(n_7),
.Y(n_237)
);

OAI321xp33_ASAP7_75t_L g236 ( 
.A1(n_229),
.A2(n_69),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_239),
.C(n_9),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_235),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_241),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_69),
.C(n_9),
.Y(n_241)
);


endmodule