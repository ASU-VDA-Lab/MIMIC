module real_jpeg_25490_n_30 (n_17, n_8, n_0, n_21, n_141, n_2, n_142, n_29, n_143, n_10, n_9, n_12, n_147, n_24, n_146, n_6, n_28, n_23, n_11, n_14, n_25, n_7, n_22, n_18, n_3, n_145, n_144, n_5, n_4, n_150, n_1, n_26, n_27, n_20, n_19, n_148, n_149, n_16, n_15, n_13, n_30);

input n_17;
input n_8;
input n_0;
input n_21;
input n_141;
input n_2;
input n_142;
input n_29;
input n_143;
input n_10;
input n_9;
input n_12;
input n_147;
input n_24;
input n_146;
input n_6;
input n_28;
input n_23;
input n_11;
input n_14;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_145;
input n_144;
input n_5;
input n_4;
input n_150;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_148;
input n_149;
input n_16;
input n_15;
input n_13;

output n_30;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_0),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_0),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_1),
.B(n_55),
.C(n_76),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_2),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_3),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_4),
.B(n_43),
.C(n_125),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_5),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_6),
.B(n_57),
.C(n_68),
.Y(n_56)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_7),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_8),
.B(n_51),
.C(n_92),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_9),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_10),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_11),
.B(n_49),
.C(n_101),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_12),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_13),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_14),
.B(n_41),
.C(n_135),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_17),
.Y(n_139)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_19),
.B(n_47),
.C(n_110),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_20),
.Y(n_121)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_22),
.Y(n_115)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_24),
.B(n_45),
.C(n_116),
.Y(n_44)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_25),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_26),
.B(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_27),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_28),
.B(n_53),
.C(n_83),
.Y(n_52)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_39),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_36),
.B(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_36),
.B(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_36),
.B(n_117),
.Y(n_116)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_37),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_40),
.C(n_137),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_42),
.C(n_131),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_118),
.C(n_119),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_112),
.C(n_113),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_104),
.C(n_105),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_95),
.C(n_96),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_86),
.C(n_87),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_78),
.C(n_79),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_71),
.C(n_72),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_63),
.C(n_64),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_141),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_142),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_143),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_144),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_145),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_146),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_147),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_148),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_149),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_150),
.Y(n_98)
);


endmodule