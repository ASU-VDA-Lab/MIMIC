module fake_aes_8644_n_13 (n_1, n_2, n_0, n_13);
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
CKINVDCx8_ASAP7_75t_R g3 ( .A(n_2), .Y(n_3) );
INVx2_ASAP7_75t_L g4 ( .A(n_0), .Y(n_4) );
INVx1_ASAP7_75t_SL g5 ( .A(n_4), .Y(n_5) );
AND2x4_ASAP7_75t_L g6 ( .A(n_3), .B(n_0), .Y(n_6) );
OAI21xp5_ASAP7_75t_L g7 ( .A1(n_5), .A2(n_0), .B(n_1), .Y(n_7) );
OAI221xp5_ASAP7_75t_L g8 ( .A1(n_5), .A2(n_0), .B1(n_1), .B2(n_2), .C(n_6), .Y(n_8) );
INVx1_ASAP7_75t_SL g9 ( .A(n_7), .Y(n_9) );
AOI22xp5_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_6), .B1(n_8), .B2(n_2), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_9), .Y(n_11) );
NAND3xp33_ASAP7_75t_L g12 ( .A(n_10), .B(n_6), .C(n_1), .Y(n_12) );
AOI22x1_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_6), .B1(n_11), .B2(n_1), .Y(n_13) );
endmodule