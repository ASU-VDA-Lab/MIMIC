module fake_ibex_273_n_1470 (n_151, n_147, n_85, n_167, n_128, n_208, n_234, n_84, n_64, n_244, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_247, n_55, n_130, n_63, n_98, n_129, n_161, n_237, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_233, n_8, n_118, n_224, n_183, n_245, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_27, n_165, n_242, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_240, n_61, n_201, n_14, n_0, n_239, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_80, n_172, n_215, n_49, n_40, n_66, n_17, n_74, n_90, n_235, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_236, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_248, n_92, n_144, n_170, n_213, n_101, n_190, n_113, n_138, n_230, n_96, n_185, n_241, n_68, n_117, n_214, n_238, n_79, n_81, n_35, n_159, n_202, n_231, n_158, n_211, n_218, n_132, n_174, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_246, n_31, n_56, n_23, n_146, n_232, n_91, n_207, n_54, n_243, n_19, n_228, n_1470);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_208;
input n_234;
input n_84;
input n_64;
input n_244;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_247;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_237;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_233;
input n_8;
input n_118;
input n_224;
input n_183;
input n_245;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_242;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_240;
input n_61;
input n_201;
input n_14;
input n_0;
input n_239;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_80;
input n_172;
input n_215;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_235;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_236;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_248;
input n_92;
input n_144;
input n_170;
input n_213;
input n_101;
input n_190;
input n_113;
input n_138;
input n_230;
input n_96;
input n_185;
input n_241;
input n_68;
input n_117;
input n_214;
input n_238;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_158;
input n_211;
input n_218;
input n_132;
input n_174;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_246;
input n_31;
input n_56;
input n_23;
input n_146;
input n_232;
input n_91;
input n_207;
input n_54;
input n_243;
input n_19;
input n_228;

output n_1470;

wire n_1084;
wire n_1295;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_1382;
wire n_273;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1134;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_280;
wire n_375;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_1463;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_641;
wire n_557;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_279;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_1449;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_359;
wire n_1466;
wire n_1412;
wire n_262;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_1401;
wire n_369;
wire n_1301;
wire n_257;
wire n_869;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_562;
wire n_564;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_314;
wire n_563;
wire n_881;
wire n_734;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_288;
wire n_379;
wire n_551;
wire n_729;
wire n_1434;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_1467;
wire n_544;
wire n_1281;
wire n_1447;
wire n_695;
wire n_639;
wire n_1332;
wire n_482;
wire n_282;
wire n_1424;
wire n_870;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_252;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_1425;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_256;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_258;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1452;
wire n_1318;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_840;
wire n_1421;
wire n_1203;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1364;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_295;
wire n_1120;
wire n_576;
wire n_388;
wire n_1279;
wire n_290;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_267;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_998;
wire n_1115;
wire n_1395;
wire n_801;
wire n_1046;
wire n_882;
wire n_942;
wire n_1431;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_444;
wire n_986;
wire n_495;
wire n_1420;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_272;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_1439;
wire n_863;
wire n_597;
wire n_285;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_318;
wire n_291;
wire n_268;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_303;
wire n_717;
wire n_1357;
wire n_668;
wire n_871;
wire n_266;
wire n_1339;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_460;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_260;
wire n_836;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1163;
wire n_677;
wire n_964;
wire n_916;
wire n_503;
wire n_292;
wire n_895;
wire n_687;
wire n_1035;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_281;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_255;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_991;
wire n_961;
wire n_1331;
wire n_1349;
wire n_1223;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1429;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_317;
wire n_1458;
wire n_1460;
wire n_326;
wire n_270;
wire n_1340;
wire n_259;
wire n_276;
wire n_339;
wire n_348;
wire n_674;
wire n_287;
wire n_552;
wire n_251;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_400;
wire n_1055;
wire n_673;
wire n_798;
wire n_278;
wire n_404;
wire n_1177;
wire n_1025;
wire n_296;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_289;
wire n_716;
wire n_923;
wire n_642;
wire n_286;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1188;
wire n_261;
wire n_742;
wire n_1191;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_595;
wire n_1001;
wire n_269;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_922;
wire n_851;
wire n_993;
wire n_253;
wire n_300;
wire n_1135;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_1066;
wire n_648;
wire n_571;
wire n_1169;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_1337;
wire n_839;
wire n_768;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_1406;
wire n_804;
wire n_484;
wire n_1455;
wire n_480;
wire n_1057;
wire n_354;
wire n_516;
wire n_1403;
wire n_329;
wire n_1149;
wire n_1176;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_277;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_1371;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1221;
wire n_284;
wire n_1047;
wire n_1374;
wire n_1435;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_302;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_298;
wire n_1256;
wire n_587;
wire n_1303;
wire n_764;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1257;
wire n_274;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1362;
wire n_1097;
wire n_293;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_1330;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_249;
wire n_1443;
wire n_478;
wire n_336;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_828;
wire n_1438;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_265;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1297;
wire n_1369;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_898;
wire n_928;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1381;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_1419;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1074;
wire n_759;
wire n_1379;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_335;
wire n_263;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_305;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1089;
wire n_392;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_283;
wire n_366;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_322;
wire n_888;
wire n_1325;
wire n_582;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_264;
wire n_1145;
wire n_537;
wire n_1113;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1354;
wire n_1277;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_294;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_1287;
wire n_860;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_297;
wire n_921;
wire n_489;
wire n_254;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_271;
wire n_1393;
wire n_984;
wire n_394;
wire n_364;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

BUFx2_ASAP7_75t_L g249 ( 
.A(n_35),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_206),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_205),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_33),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_226),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_6),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_57),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_159),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_236),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_88),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_54),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_201),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_154),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_26),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_4),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_179),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_172),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_93),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_120),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_47),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_186),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_41),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_196),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_191),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_173),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_202),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_162),
.Y(n_276)
);

BUFx8_ASAP7_75t_SL g277 ( 
.A(n_165),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_24),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_11),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_112),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_82),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_176),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_13),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_5),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_38),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_63),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_82),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_66),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_184),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_174),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_12),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_83),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_213),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_144),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_46),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_58),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_225),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_2),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_43),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_177),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_30),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_183),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_138),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_247),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_170),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_96),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_195),
.Y(n_307)
);

INVxp33_ASAP7_75t_L g308 ( 
.A(n_43),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_190),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_42),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_42),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_125),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_24),
.Y(n_313)
);

INVxp33_ASAP7_75t_L g314 ( 
.A(n_32),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_217),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_113),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_31),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_74),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_220),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_101),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_16),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_28),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_66),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_209),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_233),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_142),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_232),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_222),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_239),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_135),
.Y(n_330)
);

NOR2xp67_ASAP7_75t_L g331 ( 
.A(n_31),
.B(n_175),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_134),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_123),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_110),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_235),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_15),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_28),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_15),
.Y(n_338)
);

BUFx2_ASAP7_75t_SL g339 ( 
.A(n_5),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_17),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_129),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_53),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_30),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_178),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_163),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_153),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_180),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_224),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_198),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_223),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_3),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_87),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_143),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_203),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_12),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_151),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_133),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_76),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_88),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_84),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_242),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_156),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_61),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_116),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_60),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_23),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_51),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_72),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_67),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_166),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_193),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_81),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_41),
.Y(n_373)
);

OR2x2_ASAP7_75t_L g374 ( 
.A(n_234),
.B(n_103),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_139),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_36),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_13),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_240),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_25),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_59),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_130),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_237),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_185),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_168),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_50),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_69),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_181),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_20),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_R g389 ( 
.A(n_57),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_145),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_192),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_54),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_117),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_95),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_218),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_32),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_119),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_99),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_56),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_22),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_97),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_230),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_33),
.Y(n_403)
);

INVx1_ASAP7_75t_SL g404 ( 
.A(n_29),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_169),
.B(n_7),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_149),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_64),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_212),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_211),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_219),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_107),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_115),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_35),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_131),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_238),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_157),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_216),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_171),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_200),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_6),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_221),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_34),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_160),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_36),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_231),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_244),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_245),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_215),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_78),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_246),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_23),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_78),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_53),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_208),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_38),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_167),
.Y(n_436)
);

BUFx10_ASAP7_75t_L g437 ( 
.A(n_121),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_204),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_227),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_114),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_194),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_18),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_241),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_249),
.B(n_292),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_297),
.B(n_0),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_256),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_308),
.B(n_0),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_266),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_266),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_258),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_308),
.B(n_1),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_300),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_258),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_429),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_277),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_256),
.Y(n_456)
);

OAI21x1_ASAP7_75t_L g457 ( 
.A1(n_300),
.A2(n_100),
.B(n_98),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_304),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_255),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_406),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_406),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_414),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_411),
.B(n_415),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_256),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_255),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_414),
.Y(n_466)
);

OA21x2_ASAP7_75t_L g467 ( 
.A1(n_416),
.A2(n_104),
.B(n_102),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_265),
.B(n_250),
.Y(n_468)
);

BUFx2_ASAP7_75t_L g469 ( 
.A(n_389),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_301),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_416),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_265),
.B(n_8),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_304),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_301),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_277),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_322),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_256),
.Y(n_477)
);

INVx5_ASAP7_75t_L g478 ( 
.A(n_276),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_314),
.B(n_9),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_280),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_389),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_314),
.B(n_10),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_322),
.Y(n_483)
);

OA21x2_ASAP7_75t_L g484 ( 
.A1(n_419),
.A2(n_106),
.B(n_105),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_343),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_419),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_304),
.Y(n_487)
);

BUFx8_ASAP7_75t_L g488 ( 
.A(n_374),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_298),
.B(n_14),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_437),
.Y(n_490)
);

INVx6_ASAP7_75t_L g491 ( 
.A(n_437),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_437),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_429),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_343),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_290),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_359),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_427),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_264),
.B(n_14),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_253),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_288),
.B(n_16),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_253),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_359),
.Y(n_502)
);

OA21x2_ASAP7_75t_L g503 ( 
.A1(n_427),
.A2(n_109),
.B(n_108),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_288),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_295),
.B(n_17),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_276),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_363),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_290),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_264),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_276),
.Y(n_510)
);

OAI22x1_ASAP7_75t_L g511 ( 
.A1(n_267),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_295),
.B(n_19),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_276),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_357),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_363),
.Y(n_515)
);

BUFx8_ASAP7_75t_L g516 ( 
.A(n_344),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_403),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_357),
.Y(n_518)
);

INVx5_ASAP7_75t_L g519 ( 
.A(n_344),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_403),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_251),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_385),
.Y(n_522)
);

OAI22x1_ASAP7_75t_L g523 ( 
.A1(n_267),
.A2(n_21),
.B1(n_22),
.B2(n_25),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_385),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_431),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_269),
.A2(n_21),
.B1(n_26),
.B2(n_27),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_431),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_257),
.Y(n_528)
);

BUFx12f_ASAP7_75t_L g529 ( 
.A(n_260),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_261),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_262),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_252),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_254),
.B(n_27),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_269),
.B(n_29),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_268),
.B(n_34),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_270),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_285),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_271),
.B(n_37),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_273),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_274),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_344),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_371),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_443),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_491),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_533),
.Y(n_545)
);

INVxp33_ASAP7_75t_L g546 ( 
.A(n_469),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_446),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_446),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_456),
.Y(n_549)
);

OAI22xp33_ASAP7_75t_L g550 ( 
.A1(n_465),
.A2(n_386),
.B1(n_394),
.B2(n_271),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_469),
.B(n_260),
.Y(n_551)
);

BUFx2_ASAP7_75t_L g552 ( 
.A(n_459),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_491),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_533),
.Y(n_554)
);

BUFx2_ASAP7_75t_L g555 ( 
.A(n_529),
.Y(n_555)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_444),
.B(n_386),
.Y(n_556)
);

BUFx6f_ASAP7_75t_SL g557 ( 
.A(n_505),
.Y(n_557)
);

INVxp33_ASAP7_75t_L g558 ( 
.A(n_509),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_533),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_516),
.Y(n_560)
);

BUFx2_ASAP7_75t_L g561 ( 
.A(n_529),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_488),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_504),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_504),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_541),
.Y(n_565)
);

NAND3xp33_ASAP7_75t_L g566 ( 
.A(n_447),
.B(n_396),
.C(n_394),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_541),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_542),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_504),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_542),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_542),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_458),
.B(n_272),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_504),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_458),
.B(n_272),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_525),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_525),
.Y(n_576)
);

AND3x2_ASAP7_75t_L g577 ( 
.A(n_447),
.B(n_263),
.C(n_259),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_525),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_458),
.B(n_396),
.Y(n_579)
);

OAI22xp33_ASAP7_75t_L g580 ( 
.A1(n_465),
.A2(n_413),
.B1(n_424),
.B2(n_407),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_478),
.Y(n_581)
);

INVx4_ASAP7_75t_L g582 ( 
.A(n_505),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_478),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_491),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_525),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_478),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_533),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_505),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_505),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_488),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_519),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_512),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_458),
.B(n_407),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_451),
.A2(n_424),
.B1(n_413),
.B2(n_320),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_488),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_519),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_473),
.B(n_328),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g598 ( 
.A(n_463),
.B(n_404),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_512),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_500),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_519),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_448),
.Y(n_602)
);

INVxp33_ASAP7_75t_L g603 ( 
.A(n_479),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_519),
.Y(n_604)
);

INVx4_ASAP7_75t_L g605 ( 
.A(n_473),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_500),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_524),
.Y(n_607)
);

NAND2xp33_ASAP7_75t_L g608 ( 
.A(n_530),
.B(n_371),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_482),
.A2(n_296),
.B1(n_310),
.B2(n_283),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_487),
.B(n_328),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_449),
.Y(n_611)
);

OAI22xp33_ASAP7_75t_SL g612 ( 
.A1(n_526),
.A2(n_279),
.B1(n_281),
.B2(n_278),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_519),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_487),
.B(n_329),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_452),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_524),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_452),
.Y(n_617)
);

INVxp67_ASAP7_75t_L g618 ( 
.A(n_538),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_490),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_490),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_527),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_490),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_456),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_527),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_490),
.B(n_329),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_460),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_538),
.A2(n_532),
.B1(n_530),
.B2(n_531),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_456),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_492),
.B(n_468),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_456),
.Y(n_630)
);

NAND2x1p5_ASAP7_75t_L g631 ( 
.A(n_467),
.B(n_275),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_464),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_492),
.B(n_330),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_531),
.B(n_330),
.Y(n_634)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_455),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_464),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_522),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_522),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_464),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_464),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_536),
.B(n_390),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_477),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_536),
.B(n_390),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_495),
.Y(n_644)
);

NAND3xp33_ASAP7_75t_L g645 ( 
.A(n_445),
.B(n_286),
.C(n_284),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_461),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_539),
.B(n_398),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_477),
.Y(n_648)
);

NAND2xp33_ASAP7_75t_R g649 ( 
.A(n_475),
.B(n_287),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_461),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_462),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_506),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_516),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_506),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_539),
.B(n_398),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_540),
.A2(n_317),
.B1(n_318),
.B2(n_311),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_506),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_495),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_540),
.B(n_409),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_498),
.A2(n_336),
.B1(n_337),
.B2(n_323),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_488),
.B(n_409),
.Y(n_661)
);

INVxp67_ASAP7_75t_SL g662 ( 
.A(n_534),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_480),
.B(n_303),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_462),
.Y(n_664)
);

OAI22x1_ASAP7_75t_L g665 ( 
.A1(n_526),
.A2(n_299),
.B1(n_313),
.B2(n_291),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_466),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_466),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_506),
.Y(n_668)
);

BUFx10_ASAP7_75t_L g669 ( 
.A(n_472),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_506),
.Y(n_670)
);

OR2x6_ASAP7_75t_L g671 ( 
.A(n_511),
.B(n_339),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_543),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_521),
.B(n_418),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_521),
.B(n_528),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_510),
.Y(n_675)
);

INVxp67_ASAP7_75t_SL g676 ( 
.A(n_516),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_528),
.B(n_340),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_508),
.B(n_418),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_471),
.Y(n_679)
);

OAI22xp33_ASAP7_75t_L g680 ( 
.A1(n_481),
.A2(n_320),
.B1(n_345),
.B2(n_293),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_510),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_510),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_471),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_510),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_510),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_510),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_513),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_514),
.B(n_282),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_514),
.B(n_518),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_535),
.A2(n_293),
.B1(n_354),
.B2(n_345),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_518),
.B(n_289),
.Y(n_691)
);

OR2x6_ASAP7_75t_L g692 ( 
.A(n_511),
.B(n_342),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_513),
.Y(n_693)
);

BUFx2_ASAP7_75t_L g694 ( 
.A(n_501),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_486),
.Y(n_695)
);

AND2x6_ASAP7_75t_L g696 ( 
.A(n_486),
.B(n_306),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_513),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_497),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_579),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_618),
.A2(n_354),
.B1(n_391),
.B2(n_489),
.Y(n_700)
);

OR2x2_ASAP7_75t_L g701 ( 
.A(n_598),
.B(n_454),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_673),
.B(n_450),
.Y(n_702)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_598),
.B(n_454),
.Y(n_703)
);

NAND2xp33_ASAP7_75t_L g704 ( 
.A(n_545),
.B(n_294),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_673),
.B(n_450),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_554),
.A2(n_457),
.B(n_467),
.Y(n_706)
);

NOR3xp33_ASAP7_75t_L g707 ( 
.A(n_612),
.B(n_358),
.C(n_338),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_662),
.B(n_453),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_579),
.Y(n_709)
);

NAND2xp33_ASAP7_75t_L g710 ( 
.A(n_559),
.B(n_302),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_641),
.B(n_453),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_643),
.B(n_470),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_637),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_593),
.B(n_470),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_560),
.B(n_305),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_552),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_638),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_602),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_602),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_629),
.B(n_572),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_605),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_653),
.B(n_307),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_611),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_574),
.B(n_474),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_562),
.B(n_391),
.Y(n_725)
);

AND2x2_ASAP7_75t_SL g726 ( 
.A(n_562),
.B(n_467),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_603),
.A2(n_366),
.B1(n_367),
.B2(n_365),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_611),
.Y(n_728)
);

AND2x6_ASAP7_75t_SL g729 ( 
.A(n_671),
.B(n_692),
.Y(n_729)
);

NOR2x1p5_ASAP7_75t_L g730 ( 
.A(n_556),
.B(n_493),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_644),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_546),
.B(n_476),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_590),
.B(n_315),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_597),
.B(n_483),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_626),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_614),
.B(n_483),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_605),
.B(n_485),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_626),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_605),
.B(n_485),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_646),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_619),
.B(n_494),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_SL g742 ( 
.A1(n_692),
.A2(n_352),
.B1(n_355),
.B2(n_351),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_619),
.B(n_494),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_625),
.B(n_496),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_590),
.B(n_319),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_610),
.B(n_502),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_646),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_595),
.B(n_332),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_595),
.B(n_333),
.Y(n_749)
);

NOR2xp67_ASAP7_75t_L g750 ( 
.A(n_665),
.B(n_523),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_658),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_588),
.A2(n_523),
.B1(n_515),
.B2(n_517),
.Y(n_752)
);

INVx1_ASAP7_75t_SL g753 ( 
.A(n_552),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_633),
.B(n_507),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_650),
.Y(n_755)
);

NOR2x1p5_ASAP7_75t_L g756 ( 
.A(n_566),
.B(n_369),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_SL g757 ( 
.A(n_676),
.B(n_373),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_SL g758 ( 
.A1(n_692),
.A2(n_671),
.B1(n_557),
.B2(n_589),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_603),
.B(n_515),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_627),
.B(n_517),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_550),
.A2(n_379),
.B1(n_435),
.B2(n_376),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_580),
.A2(n_368),
.B1(n_372),
.B2(n_360),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_600),
.B(n_520),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_606),
.B(n_520),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_650),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_577),
.Y(n_766)
);

XOR2xp5_ASAP7_75t_L g767 ( 
.A(n_690),
.B(n_37),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_669),
.B(n_334),
.Y(n_768)
);

OR2x6_ASAP7_75t_L g769 ( 
.A(n_555),
.B(n_377),
.Y(n_769)
);

A2O1A1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_587),
.A2(n_388),
.B(n_392),
.C(n_380),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_634),
.B(n_309),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_555),
.Y(n_772)
);

OAI22xp5_ASAP7_75t_L g773 ( 
.A1(n_609),
.A2(n_420),
.B1(n_422),
.B2(n_400),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_557),
.A2(n_558),
.B1(n_661),
.B2(n_582),
.Y(n_774)
);

NAND3xp33_ASAP7_75t_L g775 ( 
.A(n_660),
.B(n_503),
.C(n_484),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_546),
.B(n_432),
.Y(n_776)
);

INVx4_ASAP7_75t_L g777 ( 
.A(n_557),
.Y(n_777)
);

BUFx8_ASAP7_75t_L g778 ( 
.A(n_561),
.Y(n_778)
);

O2A1O1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_592),
.A2(n_442),
.B(n_316),
.C(n_324),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_582),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_651),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_651),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_669),
.B(n_346),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_620),
.B(n_347),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_599),
.A2(n_503),
.B(n_484),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_558),
.B(n_285),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_620),
.B(n_348),
.Y(n_787)
);

AND2x6_ASAP7_75t_SL g788 ( 
.A(n_671),
.B(n_405),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_622),
.B(n_349),
.Y(n_789)
);

NAND2xp33_ASAP7_75t_SL g790 ( 
.A(n_561),
.B(n_665),
.Y(n_790)
);

CKINVDCx11_ASAP7_75t_R g791 ( 
.A(n_635),
.Y(n_791)
);

OR2x2_ASAP7_75t_L g792 ( 
.A(n_594),
.B(n_694),
.Y(n_792)
);

NOR3xp33_ASAP7_75t_L g793 ( 
.A(n_680),
.B(n_325),
.C(n_312),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_679),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_683),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_589),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_551),
.B(n_335),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_647),
.B(n_375),
.Y(n_798)
);

A2O1A1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_589),
.A2(n_387),
.B(n_326),
.C(n_327),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_692),
.A2(n_616),
.B1(n_621),
.B2(n_607),
.Y(n_800)
);

NAND2xp33_ASAP7_75t_L g801 ( 
.A(n_672),
.B(n_382),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_624),
.A2(n_399),
.B1(n_285),
.B2(n_321),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_683),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_669),
.B(n_383),
.Y(n_804)
);

BUFx6f_ASAP7_75t_SL g805 ( 
.A(n_671),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_645),
.B(n_384),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_655),
.B(n_428),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_659),
.B(n_430),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_678),
.B(n_341),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_544),
.Y(n_810)
);

INVxp67_ASAP7_75t_L g811 ( 
.A(n_674),
.Y(n_811)
);

INVxp33_ASAP7_75t_L g812 ( 
.A(n_694),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_544),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_677),
.B(n_412),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_SL g815 ( 
.A1(n_663),
.A2(n_436),
.B1(n_425),
.B2(n_439),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_553),
.B(n_350),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_664),
.Y(n_817)
);

HB1xp67_ASAP7_75t_L g818 ( 
.A(n_677),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_615),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_553),
.B(n_584),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_656),
.B(n_321),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_666),
.B(n_667),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_688),
.B(n_353),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_615),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_691),
.B(n_356),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_617),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_617),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_617),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_696),
.A2(n_399),
.B1(n_433),
.B2(n_362),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_563),
.A2(n_402),
.B1(n_378),
.B2(n_361),
.Y(n_830)
);

NOR2xp67_ASAP7_75t_L g831 ( 
.A(n_695),
.B(n_537),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_695),
.Y(n_832)
);

OAI22xp33_ASAP7_75t_L g833 ( 
.A1(n_698),
.A2(n_399),
.B1(n_433),
.B2(n_331),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_563),
.B(n_364),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_564),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_569),
.B(n_573),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_689),
.B(n_433),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_575),
.Y(n_838)
);

NOR3xp33_ASAP7_75t_L g839 ( 
.A(n_575),
.B(n_393),
.C(n_370),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_696),
.B(n_395),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_576),
.B(n_397),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_576),
.B(n_401),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_SL g843 ( 
.A1(n_696),
.A2(n_433),
.B1(n_408),
.B2(n_410),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_578),
.B(n_417),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_696),
.A2(n_434),
.B1(n_421),
.B2(n_423),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_585),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_696),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_631),
.A2(n_438),
.B1(n_440),
.B2(n_441),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_547),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_631),
.B(n_371),
.Y(n_850)
);

OR2x2_ASAP7_75t_L g851 ( 
.A(n_649),
.B(n_39),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_581),
.B(n_537),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_608),
.B(n_371),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_608),
.B(n_381),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_547),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_548),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_548),
.Y(n_857)
);

AND2x6_ASAP7_75t_L g858 ( 
.A(n_583),
.B(n_381),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_583),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_586),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_753),
.B(n_716),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_812),
.B(n_39),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_777),
.B(n_40),
.Y(n_863)
);

AO22x1_ASAP7_75t_L g864 ( 
.A1(n_778),
.A2(n_426),
.B1(n_44),
.B2(n_45),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_699),
.B(n_709),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_777),
.B(n_40),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_811),
.B(n_591),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_811),
.B(n_596),
.Y(n_868)
);

A2O1A1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_746),
.A2(n_613),
.B(n_604),
.C(n_601),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_778),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_758),
.A2(n_613),
.B1(n_604),
.B2(n_601),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_818),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_780),
.Y(n_873)
);

A2O1A1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_746),
.A2(n_565),
.B(n_570),
.C(n_568),
.Y(n_874)
);

OAI22xp5_ASAP7_75t_SL g875 ( 
.A1(n_767),
.A2(n_426),
.B1(n_46),
.B2(n_47),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_720),
.B(n_714),
.Y(n_876)
);

INVx1_ASAP7_75t_SL g877 ( 
.A(n_791),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_780),
.Y(n_878)
);

AO22x1_ASAP7_75t_L g879 ( 
.A1(n_725),
.A2(n_426),
.B1(n_48),
.B2(n_49),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_725),
.B(n_45),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_769),
.Y(n_881)
);

O2A1O1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_770),
.A2(n_567),
.B(n_570),
.C(n_571),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_769),
.B(n_48),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_732),
.B(n_759),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_759),
.B(n_49),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_835),
.Y(n_886)
);

CKINVDCx20_ASAP7_75t_R g887 ( 
.A(n_772),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_838),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_726),
.A2(n_628),
.B(n_623),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_769),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_721),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_818),
.B(n_50),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_703),
.B(n_51),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_708),
.B(n_52),
.Y(n_894)
);

INVxp67_ASAP7_75t_L g895 ( 
.A(n_757),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_SL g896 ( 
.A(n_805),
.B(n_513),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_846),
.Y(n_897)
);

INVxp67_ASAP7_75t_L g898 ( 
.A(n_776),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_796),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_727),
.B(n_52),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_758),
.B(n_774),
.Y(n_901)
);

O2A1O1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_773),
.A2(n_697),
.B(n_693),
.C(n_687),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_850),
.A2(n_632),
.B(n_630),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_796),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_702),
.B(n_55),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_714),
.B(n_55),
.Y(n_906)
);

BUFx4f_ASAP7_75t_L g907 ( 
.A(n_766),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_839),
.A2(n_707),
.B1(n_756),
.B2(n_750),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_700),
.A2(n_693),
.B1(n_686),
.B2(n_685),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_792),
.B(n_56),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_763),
.Y(n_911)
);

O2A1O1Ixp33_ASAP7_75t_SL g912 ( 
.A1(n_799),
.A2(n_685),
.B(n_684),
.C(n_681),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_815),
.B(n_58),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_850),
.A2(n_640),
.B(n_636),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_764),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_797),
.B(n_59),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_786),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_768),
.B(n_783),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_800),
.B(n_60),
.Y(n_919)
);

INVx1_ASAP7_75t_SL g920 ( 
.A(n_851),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_737),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_739),
.Y(n_922)
);

NOR2x1_ASAP7_75t_L g923 ( 
.A(n_804),
.B(n_642),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_836),
.A2(n_743),
.B(n_741),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_705),
.Y(n_925)
);

O2A1O1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_760),
.A2(n_684),
.B(n_681),
.C(n_675),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_848),
.A2(n_648),
.B1(n_652),
.B2(n_654),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_718),
.B(n_61),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_SL g929 ( 
.A(n_805),
.B(n_652),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_719),
.B(n_723),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_860),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_728),
.B(n_62),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_852),
.Y(n_933)
);

NAND3xp33_ASAP7_75t_SL g934 ( 
.A(n_752),
.B(n_654),
.C(n_657),
.Y(n_934)
);

INVxp67_ASAP7_75t_L g935 ( 
.A(n_814),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_733),
.B(n_745),
.Y(n_936)
);

BUFx12f_ASAP7_75t_L g937 ( 
.A(n_729),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_822),
.A2(n_657),
.B1(n_668),
.B2(n_670),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_748),
.B(n_62),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_735),
.B(n_738),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_740),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_747),
.B(n_63),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_755),
.B(n_64),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_749),
.B(n_65),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_713),
.Y(n_945)
);

INVx4_ASAP7_75t_L g946 ( 
.A(n_824),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_761),
.B(n_65),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_798),
.B(n_807),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_779),
.A2(n_682),
.B(n_639),
.C(n_549),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_704),
.A2(n_710),
.B(n_711),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_712),
.A2(n_682),
.B(n_639),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_765),
.B(n_67),
.Y(n_952)
);

INVx1_ASAP7_75t_SL g953 ( 
.A(n_821),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_844),
.A2(n_782),
.B(n_781),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_717),
.B(n_68),
.Y(n_955)
);

NOR2xp67_ASAP7_75t_L g956 ( 
.A(n_762),
.B(n_69),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_825),
.B(n_70),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_SL g958 ( 
.A1(n_820),
.A2(n_549),
.B(n_161),
.C(n_164),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_730),
.B(n_70),
.Y(n_959)
);

NOR3xp33_ASAP7_75t_L g960 ( 
.A(n_790),
.B(n_71),
.C(n_72),
.Y(n_960)
);

NOR2x1p5_ASAP7_75t_SL g961 ( 
.A(n_849),
.B(n_111),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_R g962 ( 
.A(n_801),
.B(n_71),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_794),
.B(n_73),
.Y(n_963)
);

NAND3xp33_ASAP7_75t_L g964 ( 
.A(n_742),
.B(n_73),
.C(n_74),
.Y(n_964)
);

NOR3xp33_ASAP7_75t_L g965 ( 
.A(n_742),
.B(n_806),
.C(n_808),
.Y(n_965)
);

O2A1O1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_795),
.A2(n_75),
.B(n_76),
.C(n_77),
.Y(n_966)
);

O2A1O1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_803),
.A2(n_75),
.B(n_77),
.C(n_79),
.Y(n_967)
);

OAI21xp33_ASAP7_75t_SL g968 ( 
.A1(n_752),
.A2(n_80),
.B(n_81),
.Y(n_968)
);

OR2x2_ASAP7_75t_L g969 ( 
.A(n_823),
.B(n_80),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_SL g970 ( 
.A(n_847),
.B(n_83),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_784),
.B(n_84),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_817),
.B(n_85),
.Y(n_972)
);

AOI221xp5_ASAP7_75t_L g973 ( 
.A1(n_754),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.C(n_89),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_844),
.B(n_86),
.Y(n_974)
);

NOR3xp33_ASAP7_75t_L g975 ( 
.A(n_771),
.B(n_754),
.C(n_809),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_724),
.B(n_89),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_787),
.B(n_90),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_789),
.B(n_90),
.Y(n_978)
);

NOR3xp33_ASAP7_75t_L g979 ( 
.A(n_771),
.B(n_91),
.C(n_92),
.Y(n_979)
);

INVxp67_ASAP7_75t_L g980 ( 
.A(n_809),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_724),
.B(n_91),
.Y(n_981)
);

BUFx4f_ASAP7_75t_L g982 ( 
.A(n_810),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_845),
.A2(n_736),
.B1(n_734),
.B2(n_744),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_788),
.B(n_92),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_734),
.A2(n_744),
.B(n_736),
.Y(n_985)
);

NOR2x1_ASAP7_75t_L g986 ( 
.A(n_715),
.B(n_93),
.Y(n_986)
);

INVx3_ASAP7_75t_L g987 ( 
.A(n_824),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_841),
.A2(n_182),
.B(n_229),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_842),
.B(n_94),
.Y(n_989)
);

BUFx4f_ASAP7_75t_L g990 ( 
.A(n_813),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_830),
.B(n_94),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_SL g992 ( 
.A(n_858),
.B(n_118),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_816),
.B(n_122),
.Y(n_993)
);

INVx6_ASAP7_75t_L g994 ( 
.A(n_859),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_816),
.B(n_248),
.Y(n_995)
);

AO221x2_ASAP7_75t_L g996 ( 
.A1(n_833),
.A2(n_124),
.B1(n_126),
.B2(n_127),
.C(n_128),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_731),
.A2(n_132),
.B(n_136),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_834),
.A2(n_137),
.B1(n_140),
.B2(n_141),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_837),
.Y(n_999)
);

AO21x1_ASAP7_75t_L g1000 ( 
.A1(n_833),
.A2(n_146),
.B(n_147),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_751),
.A2(n_148),
.B(n_150),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_826),
.A2(n_152),
.B(n_155),
.C(n_158),
.Y(n_1002)
);

CKINVDCx10_ASAP7_75t_R g1003 ( 
.A(n_843),
.Y(n_1003)
);

BUFx12f_ASAP7_75t_L g1004 ( 
.A(n_858),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_843),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_855),
.A2(n_197),
.B(n_199),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_856),
.A2(n_207),
.B(n_210),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_925),
.B(n_722),
.Y(n_1008)
);

OAI21x1_ASAP7_75t_SL g1009 ( 
.A1(n_930),
.A2(n_840),
.B(n_827),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_911),
.B(n_819),
.Y(n_1010)
);

AO31x2_ASAP7_75t_L g1011 ( 
.A1(n_1000),
.A2(n_854),
.A3(n_853),
.B(n_828),
.Y(n_1011)
);

INVxp67_ASAP7_75t_SL g1012 ( 
.A(n_861),
.Y(n_1012)
);

AO22x2_ASAP7_75t_L g1013 ( 
.A1(n_955),
.A2(n_832),
.B1(n_857),
.B2(n_829),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_870),
.Y(n_1014)
);

OAI22xp33_ASAP7_75t_L g1015 ( 
.A1(n_890),
.A2(n_831),
.B1(n_859),
.B2(n_854),
.Y(n_1015)
);

AO31x2_ASAP7_75t_L g1016 ( 
.A1(n_889),
.A2(n_853),
.A3(n_829),
.B(n_802),
.Y(n_1016)
);

NOR2xp67_ASAP7_75t_L g1017 ( 
.A(n_937),
.B(n_214),
.Y(n_1017)
);

OR2x6_ASAP7_75t_L g1018 ( 
.A(n_881),
.B(n_228),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_948),
.A2(n_950),
.B(n_916),
.C(n_954),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_945),
.Y(n_1020)
);

AO21x2_ASAP7_75t_L g1021 ( 
.A1(n_934),
.A2(n_988),
.B(n_1006),
.Y(n_1021)
);

INVx1_ASAP7_75t_SL g1022 ( 
.A(n_887),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_865),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_936),
.B(n_872),
.Y(n_1024)
);

OAI21xp33_ASAP7_75t_L g1025 ( 
.A1(n_884),
.A2(n_910),
.B(n_893),
.Y(n_1025)
);

INVxp67_ASAP7_75t_SL g1026 ( 
.A(n_955),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_877),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_935),
.B(n_980),
.Y(n_1028)
);

BUFx12f_ASAP7_75t_L g1029 ( 
.A(n_863),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_930),
.A2(n_940),
.B1(n_922),
.B2(n_921),
.Y(n_1030)
);

BUFx2_ASAP7_75t_L g1031 ( 
.A(n_863),
.Y(n_1031)
);

INVxp67_ASAP7_75t_SL g1032 ( 
.A(n_867),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_1004),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_940),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_907),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_975),
.A2(n_906),
.B(n_974),
.C(n_968),
.Y(n_1036)
);

AO32x2_ASAP7_75t_L g1037 ( 
.A1(n_871),
.A2(n_983),
.A3(n_909),
.B1(n_1005),
.B2(n_938),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_951),
.A2(n_914),
.B(n_903),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_898),
.B(n_941),
.Y(n_1039)
);

BUFx4_ASAP7_75t_SL g1040 ( 
.A(n_964),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_906),
.A2(n_974),
.B(n_985),
.C(n_885),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_895),
.B(n_962),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_865),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_SL g1044 ( 
.A1(n_996),
.A2(n_866),
.B(n_1007),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_880),
.B(n_908),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_SL g1046 ( 
.A1(n_919),
.A2(n_868),
.B(n_867),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_886),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_899),
.B(n_904),
.Y(n_1048)
);

HB1xp67_ASAP7_75t_L g1049 ( 
.A(n_866),
.Y(n_1049)
);

AO31x2_ASAP7_75t_L g1050 ( 
.A1(n_869),
.A2(n_949),
.A3(n_1002),
.B(n_952),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_946),
.Y(n_1051)
);

AOI21xp33_ASAP7_75t_L g1052 ( 
.A1(n_920),
.A2(n_918),
.B(n_892),
.Y(n_1052)
);

BUFx2_ASAP7_75t_R g1053 ( 
.A(n_901),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_913),
.B(n_883),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_953),
.B(n_900),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_989),
.A2(n_991),
.B(n_905),
.C(n_967),
.Y(n_1056)
);

OR2x6_ASAP7_75t_L g1057 ( 
.A(n_879),
.B(n_864),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_888),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_SL g1059 ( 
.A1(n_996),
.A2(n_993),
.B(n_995),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_936),
.B(n_965),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_947),
.B(n_868),
.Y(n_1061)
);

INVx5_ASAP7_75t_L g1062 ( 
.A(n_931),
.Y(n_1062)
);

OR2x2_ASAP7_75t_L g1063 ( 
.A(n_933),
.B(n_969),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_874),
.A2(n_926),
.B(n_902),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_999),
.B(n_956),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_989),
.A2(n_981),
.B(n_976),
.C(n_919),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_959),
.B(n_862),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_928),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_976),
.A2(n_981),
.B(n_966),
.C(n_894),
.Y(n_1069)
);

INVxp67_ASAP7_75t_L g1070 ( 
.A(n_957),
.Y(n_1070)
);

AO22x2_ASAP7_75t_L g1071 ( 
.A1(n_957),
.A2(n_960),
.B1(n_1003),
.B2(n_979),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_982),
.B(n_990),
.Y(n_1072)
);

AO32x2_ASAP7_75t_L g1073 ( 
.A1(n_875),
.A2(n_917),
.A3(n_927),
.B1(n_961),
.B2(n_912),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_932),
.A2(n_963),
.B(n_942),
.C(n_943),
.Y(n_1074)
);

OR2x2_ASAP7_75t_L g1075 ( 
.A(n_991),
.B(n_972),
.Y(n_1075)
);

INVx1_ASAP7_75t_SL g1076 ( 
.A(n_942),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_943),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_971),
.Y(n_1078)
);

BUFx12f_ASAP7_75t_L g1079 ( 
.A(n_982),
.Y(n_1079)
);

NAND3x1_ASAP7_75t_L g1080 ( 
.A(n_984),
.B(n_973),
.C(n_986),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_990),
.B(n_944),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_939),
.B(n_977),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_978),
.Y(n_1083)
);

INVx4_ASAP7_75t_L g1084 ( 
.A(n_891),
.Y(n_1084)
);

AO31x2_ASAP7_75t_L g1085 ( 
.A1(n_997),
.A2(n_1001),
.A3(n_958),
.B(n_878),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_873),
.A2(n_882),
.B(n_923),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_987),
.B(n_929),
.Y(n_1087)
);

O2A1O1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_970),
.A2(n_896),
.B(n_992),
.C(n_998),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_994),
.A2(n_753),
.B1(n_501),
.B2(n_499),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_911),
.B(n_915),
.Y(n_1090)
);

AO31x2_ASAP7_75t_L g1091 ( 
.A1(n_1000),
.A2(n_706),
.A3(n_785),
.B(n_889),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_930),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_925),
.B(n_911),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_911),
.B(n_915),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_881),
.B(n_701),
.Y(n_1095)
);

INVx2_ASAP7_75t_SL g1096 ( 
.A(n_870),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_911),
.B(n_915),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_925),
.B(n_911),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_911),
.A2(n_915),
.B1(n_876),
.B2(n_925),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_911),
.A2(n_915),
.B1(n_876),
.B2(n_925),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_876),
.A2(n_775),
.B(n_924),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_1004),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_911),
.B(n_915),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_930),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_R g1105 ( 
.A(n_887),
.B(n_778),
.Y(n_1105)
);

AO31x2_ASAP7_75t_L g1106 ( 
.A1(n_1000),
.A2(n_706),
.A3(n_785),
.B(n_889),
.Y(n_1106)
);

NAND3xp33_ASAP7_75t_L g1107 ( 
.A(n_916),
.B(n_707),
.C(n_488),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_930),
.Y(n_1108)
);

INVx1_ASAP7_75t_SL g1109 ( 
.A(n_861),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_870),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_876),
.A2(n_775),
.B(n_924),
.Y(n_1111)
);

NAND2xp33_ASAP7_75t_R g1112 ( 
.A(n_870),
.B(n_499),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_911),
.B(n_915),
.Y(n_1113)
);

NAND3x1_ASAP7_75t_L g1114 ( 
.A(n_984),
.B(n_465),
.C(n_793),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_930),
.Y(n_1115)
);

OAI21xp33_ASAP7_75t_SL g1116 ( 
.A1(n_930),
.A2(n_940),
.B(n_876),
.Y(n_1116)
);

INVx4_ASAP7_75t_L g1117 ( 
.A(n_870),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_876),
.A2(n_775),
.B(n_924),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_911),
.B(n_915),
.Y(n_1119)
);

AO31x2_ASAP7_75t_L g1120 ( 
.A1(n_1000),
.A2(n_706),
.A3(n_785),
.B(n_889),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_890),
.B(n_757),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_SL g1122 ( 
.A1(n_930),
.A2(n_940),
.B(n_954),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_890),
.B(n_757),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_945),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_890),
.B(n_757),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_R g1126 ( 
.A(n_887),
.B(n_778),
.Y(n_1126)
);

NAND3x1_ASAP7_75t_L g1127 ( 
.A(n_984),
.B(n_465),
.C(n_793),
.Y(n_1127)
);

CKINVDCx20_ASAP7_75t_R g1128 ( 
.A(n_887),
.Y(n_1128)
);

OA22x2_ASAP7_75t_L g1129 ( 
.A1(n_890),
.A2(n_690),
.B1(n_700),
.B2(n_499),
.Y(n_1129)
);

NOR2xp67_ASAP7_75t_L g1130 ( 
.A(n_937),
.B(n_772),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_890),
.B(n_757),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_861),
.B(n_753),
.Y(n_1132)
);

AO31x2_ASAP7_75t_L g1133 ( 
.A1(n_1000),
.A2(n_706),
.A3(n_785),
.B(n_889),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_911),
.B(n_915),
.Y(n_1134)
);

BUFx10_ASAP7_75t_L g1135 ( 
.A(n_890),
.Y(n_1135)
);

NAND2x1p5_ASAP7_75t_L g1136 ( 
.A(n_870),
.B(n_753),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_890),
.B(n_757),
.Y(n_1137)
);

AOI211x1_ASAP7_75t_L g1138 ( 
.A1(n_876),
.A2(n_985),
.B(n_964),
.C(n_991),
.Y(n_1138)
);

AO31x2_ASAP7_75t_L g1139 ( 
.A1(n_1000),
.A2(n_706),
.A3(n_785),
.B(n_889),
.Y(n_1139)
);

AND3x4_ASAP7_75t_L g1140 ( 
.A(n_956),
.B(n_750),
.C(n_793),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_911),
.A2(n_915),
.B1(n_876),
.B2(n_925),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_890),
.B(n_757),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_897),
.Y(n_1143)
);

AO31x2_ASAP7_75t_L g1144 ( 
.A1(n_1000),
.A2(n_706),
.A3(n_785),
.B(n_889),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_881),
.B(n_701),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_945),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_861),
.B(n_753),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_861),
.B(n_753),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1116),
.A2(n_1030),
.B(n_1122),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1090),
.Y(n_1150)
);

BUFx2_ASAP7_75t_L g1151 ( 
.A(n_1128),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1043),
.B(n_1023),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_1136),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1132),
.B(n_1147),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_1032),
.A2(n_1099),
.B1(n_1141),
.B2(n_1100),
.Y(n_1155)
);

INVx3_ASAP7_75t_L g1156 ( 
.A(n_1093),
.Y(n_1156)
);

INVx4_ASAP7_75t_L g1157 ( 
.A(n_1079),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1094),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1097),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_1105),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_1092),
.Y(n_1161)
);

OA21x2_ASAP7_75t_L g1162 ( 
.A1(n_1064),
.A2(n_1111),
.B(n_1101),
.Y(n_1162)
);

NAND3xp33_ASAP7_75t_L g1163 ( 
.A(n_1107),
.B(n_1138),
.C(n_1019),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_SL g1164 ( 
.A1(n_1046),
.A2(n_1009),
.B(n_1088),
.Y(n_1164)
);

OR2x2_ASAP7_75t_L g1165 ( 
.A(n_1109),
.B(n_1028),
.Y(n_1165)
);

AO21x2_ASAP7_75t_L g1166 ( 
.A1(n_1059),
.A2(n_1021),
.B(n_1118),
.Y(n_1166)
);

AO31x2_ASAP7_75t_L g1167 ( 
.A1(n_1036),
.A2(n_1069),
.A3(n_1038),
.B(n_1068),
.Y(n_1167)
);

OAI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1056),
.A2(n_1061),
.B(n_1080),
.Y(n_1168)
);

BUFx2_ASAP7_75t_L g1169 ( 
.A(n_1126),
.Y(n_1169)
);

OR2x6_ASAP7_75t_L g1170 ( 
.A(n_1029),
.B(n_1018),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1104),
.B(n_1108),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_1104),
.B(n_1108),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1103),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_1033),
.Y(n_1174)
);

INVx1_ASAP7_75t_SL g1175 ( 
.A(n_1022),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1113),
.Y(n_1176)
);

OR2x2_ASAP7_75t_L g1177 ( 
.A(n_1148),
.B(n_1012),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1119),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1134),
.Y(n_1179)
);

AO31x2_ASAP7_75t_L g1180 ( 
.A1(n_1068),
.A2(n_1086),
.A3(n_1060),
.B(n_1077),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1020),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1124),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1087),
.A2(n_1044),
.B(n_1051),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1054),
.B(n_1095),
.Y(n_1184)
);

HB1xp67_ASAP7_75t_L g1185 ( 
.A(n_1115),
.Y(n_1185)
);

OA21x2_ASAP7_75t_L g1186 ( 
.A1(n_1082),
.A2(n_1078),
.B(n_1083),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_SL g1187 ( 
.A1(n_1084),
.A2(n_1075),
.B(n_1143),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1047),
.Y(n_1188)
);

OAI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1076),
.A2(n_1045),
.B(n_1065),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1071),
.A2(n_1140),
.B1(n_1129),
.B2(n_1055),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1145),
.B(n_1039),
.Y(n_1191)
);

AO31x2_ASAP7_75t_L g1192 ( 
.A1(n_1058),
.A2(n_1037),
.A3(n_1011),
.B(n_1146),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1048),
.Y(n_1193)
);

OR2x2_ASAP7_75t_L g1194 ( 
.A(n_1089),
.B(n_1031),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1026),
.B(n_1070),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_1008),
.B(n_1024),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1013),
.A2(n_1010),
.B(n_1052),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_1062),
.Y(n_1198)
);

CKINVDCx20_ASAP7_75t_R g1199 ( 
.A(n_1027),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1008),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1015),
.A2(n_1125),
.B(n_1142),
.Y(n_1201)
);

INVx6_ASAP7_75t_L g1202 ( 
.A(n_1062),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_1049),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1121),
.A2(n_1137),
.B(n_1131),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1114),
.A2(n_1127),
.B(n_1067),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_1024),
.B(n_1063),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1018),
.Y(n_1207)
);

AOI21xp33_ASAP7_75t_SL g1208 ( 
.A1(n_1071),
.A2(n_1112),
.B(n_1042),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1091),
.A2(n_1144),
.B(n_1139),
.Y(n_1209)
);

INVx2_ASAP7_75t_SL g1210 ( 
.A(n_1135),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_1057),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1040),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1081),
.B(n_1123),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1033),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1096),
.B(n_1110),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_1062),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_1033),
.Y(n_1217)
);

OAI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1057),
.A2(n_1017),
.B(n_1072),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1106),
.Y(n_1219)
);

INVxp67_ASAP7_75t_L g1220 ( 
.A(n_1053),
.Y(n_1220)
);

BUFx8_ASAP7_75t_SL g1221 ( 
.A(n_1014),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1037),
.A2(n_1130),
.B(n_1073),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1135),
.B(n_1117),
.Y(n_1223)
);

INVx2_ASAP7_75t_SL g1224 ( 
.A(n_1035),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1117),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1050),
.Y(n_1226)
);

INVx6_ASAP7_75t_L g1227 ( 
.A(n_1102),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1102),
.B(n_1011),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1120),
.A2(n_1133),
.B(n_1085),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1120),
.A2(n_1085),
.B(n_1073),
.Y(n_1230)
);

AO31x2_ASAP7_75t_L g1231 ( 
.A1(n_1085),
.A2(n_1066),
.A3(n_1041),
.B(n_1074),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1016),
.Y(n_1232)
);

INVx3_ASAP7_75t_SL g1233 ( 
.A(n_1128),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1025),
.A2(n_793),
.B1(n_1030),
.B2(n_1099),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_1034),
.B(n_1092),
.Y(n_1235)
);

OR2x6_ASAP7_75t_L g1236 ( 
.A(n_1029),
.B(n_1018),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1116),
.A2(n_1030),
.B(n_1122),
.Y(n_1237)
);

NOR2x1_ASAP7_75t_R g1238 ( 
.A(n_1029),
.B(n_791),
.Y(n_1238)
);

CKINVDCx11_ASAP7_75t_R g1239 ( 
.A(n_1128),
.Y(n_1239)
);

CKINVDCx11_ASAP7_75t_R g1240 ( 
.A(n_1128),
.Y(n_1240)
);

NAND2x1p5_ASAP7_75t_L g1241 ( 
.A(n_1093),
.B(n_1098),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1043),
.B(n_1023),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1030),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1043),
.B(n_1023),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_SL g1245 ( 
.A1(n_1116),
.A2(n_501),
.B1(n_1026),
.B2(n_1030),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_1154),
.Y(n_1246)
);

INVx1_ASAP7_75t_SL g1247 ( 
.A(n_1161),
.Y(n_1247)
);

OR2x2_ASAP7_75t_L g1248 ( 
.A(n_1161),
.B(n_1185),
.Y(n_1248)
);

BUFx3_ASAP7_75t_L g1249 ( 
.A(n_1241),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1243),
.Y(n_1250)
);

OR2x2_ASAP7_75t_L g1251 ( 
.A(n_1185),
.B(n_1177),
.Y(n_1251)
);

OR2x6_ASAP7_75t_L g1252 ( 
.A(n_1149),
.B(n_1237),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1188),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1243),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1171),
.B(n_1172),
.Y(n_1255)
);

OR2x2_ASAP7_75t_L g1256 ( 
.A(n_1172),
.B(n_1235),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1180),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1219),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_1165),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1167),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1167),
.Y(n_1261)
);

CKINVDCx6p67_ASAP7_75t_R g1262 ( 
.A(n_1233),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1153),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1150),
.B(n_1158),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_SL g1265 ( 
.A1(n_1155),
.A2(n_1236),
.B(n_1170),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1167),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1198),
.Y(n_1267)
);

INVx1_ASAP7_75t_SL g1268 ( 
.A(n_1198),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1245),
.B(n_1159),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1192),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1192),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1192),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_1202),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1245),
.B(n_1173),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1192),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1152),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1242),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1244),
.Y(n_1278)
);

NOR2xp67_ASAP7_75t_L g1279 ( 
.A(n_1163),
.B(n_1222),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1209),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1183),
.B(n_1211),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1176),
.Y(n_1282)
);

OR2x6_ASAP7_75t_L g1283 ( 
.A(n_1164),
.B(n_1211),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1178),
.B(n_1179),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1187),
.Y(n_1285)
);

INVxp67_ASAP7_75t_L g1286 ( 
.A(n_1285),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1247),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1253),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_1285),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1247),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1246),
.B(n_1233),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1276),
.B(n_1168),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1269),
.A2(n_1205),
.B1(n_1190),
.B2(n_1170),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1260),
.B(n_1261),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1260),
.B(n_1226),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1281),
.B(n_1229),
.Y(n_1296)
);

OR2x2_ASAP7_75t_L g1297 ( 
.A(n_1248),
.B(n_1228),
.Y(n_1297)
);

BUFx3_ASAP7_75t_L g1298 ( 
.A(n_1285),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_1248),
.Y(n_1299)
);

BUFx2_ASAP7_75t_L g1300 ( 
.A(n_1281),
.Y(n_1300)
);

BUFx2_ASAP7_75t_L g1301 ( 
.A(n_1283),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_L g1302 ( 
.A(n_1258),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1266),
.B(n_1232),
.Y(n_1303)
);

OAI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1262),
.A2(n_1170),
.B1(n_1236),
.B2(n_1220),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1269),
.A2(n_1190),
.B1(n_1236),
.B2(n_1234),
.Y(n_1305)
);

OA222x2_ASAP7_75t_L g1306 ( 
.A1(n_1251),
.A2(n_1256),
.B1(n_1255),
.B2(n_1283),
.C1(n_1265),
.C2(n_1249),
.Y(n_1306)
);

OR2x2_ASAP7_75t_L g1307 ( 
.A(n_1251),
.B(n_1162),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1270),
.B(n_1162),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1257),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1277),
.B(n_1278),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1277),
.B(n_1234),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1252),
.B(n_1166),
.Y(n_1312)
);

AND2x4_ASAP7_75t_L g1313 ( 
.A(n_1252),
.B(n_1230),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1257),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1250),
.B(n_1231),
.Y(n_1315)
);

OAI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1262),
.A2(n_1220),
.B1(n_1194),
.B2(n_1156),
.Y(n_1316)
);

NAND3xp33_ASAP7_75t_L g1317 ( 
.A(n_1265),
.B(n_1204),
.C(n_1208),
.Y(n_1317)
);

AOI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1274),
.A2(n_1184),
.B1(n_1191),
.B2(n_1193),
.Y(n_1318)
);

NOR2xp67_ASAP7_75t_L g1319 ( 
.A(n_1267),
.B(n_1197),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1270),
.B(n_1231),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1309),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1309),
.Y(n_1322)
);

OR2x2_ASAP7_75t_L g1323 ( 
.A(n_1307),
.B(n_1250),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1314),
.Y(n_1324)
);

INVx1_ASAP7_75t_SL g1325 ( 
.A(n_1289),
.Y(n_1325)
);

INVx3_ASAP7_75t_L g1326 ( 
.A(n_1312),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1308),
.B(n_1271),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1308),
.B(n_1271),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1314),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1308),
.B(n_1272),
.Y(n_1330)
);

OR2x2_ASAP7_75t_L g1331 ( 
.A(n_1307),
.B(n_1254),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1320),
.B(n_1272),
.Y(n_1332)
);

INVx3_ASAP7_75t_L g1333 ( 
.A(n_1312),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1288),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1320),
.B(n_1275),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1318),
.B(n_1207),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1320),
.B(n_1275),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1294),
.B(n_1313),
.Y(n_1338)
);

OR2x2_ASAP7_75t_L g1339 ( 
.A(n_1297),
.B(n_1254),
.Y(n_1339)
);

INVx2_ASAP7_75t_SL g1340 ( 
.A(n_1289),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1302),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1318),
.B(n_1274),
.Y(n_1342)
);

BUFx2_ASAP7_75t_L g1343 ( 
.A(n_1286),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1294),
.B(n_1313),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1313),
.B(n_1280),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1286),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1296),
.B(n_1295),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1296),
.B(n_1252),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1323),
.B(n_1299),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1323),
.B(n_1299),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1334),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1321),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1323),
.B(n_1297),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1342),
.B(n_1311),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1321),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1348),
.Y(n_1356)
);

INVxp67_ASAP7_75t_L g1357 ( 
.A(n_1343),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1322),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1322),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1324),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1341),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1338),
.B(n_1303),
.Y(n_1362)
);

NOR2x1p5_ASAP7_75t_L g1363 ( 
.A(n_1326),
.B(n_1317),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1324),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1329),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1334),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1338),
.B(n_1344),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1338),
.B(n_1303),
.Y(n_1368)
);

OR2x2_ASAP7_75t_L g1369 ( 
.A(n_1331),
.B(n_1315),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_1353),
.Y(n_1370)
);

AOI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1354),
.A2(n_1342),
.B1(n_1336),
.B2(n_1305),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1361),
.B(n_1332),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1352),
.Y(n_1373)
);

AOI322xp5_ASAP7_75t_L g1374 ( 
.A1(n_1362),
.A2(n_1304),
.A3(n_1293),
.B1(n_1336),
.B2(n_1316),
.C1(n_1291),
.C2(n_1344),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1352),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1355),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1369),
.B(n_1331),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1369),
.B(n_1331),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1355),
.Y(n_1379)
);

OA21x2_ASAP7_75t_L g1380 ( 
.A1(n_1357),
.A2(n_1319),
.B(n_1345),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_SL g1381 ( 
.A(n_1356),
.B(n_1340),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1367),
.B(n_1344),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1353),
.B(n_1332),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1362),
.B(n_1332),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1356),
.B(n_1348),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1358),
.Y(n_1386)
);

INVxp67_ASAP7_75t_L g1387 ( 
.A(n_1349),
.Y(n_1387)
);

AOI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1371),
.A2(n_1363),
.B1(n_1368),
.B2(n_1317),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1387),
.B(n_1370),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1377),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1377),
.A2(n_1356),
.B1(n_1349),
.B2(n_1350),
.Y(n_1391)
);

AOI321xp33_ASAP7_75t_SL g1392 ( 
.A1(n_1374),
.A2(n_1175),
.A3(n_1306),
.B1(n_1325),
.B2(n_1238),
.C(n_1240),
.Y(n_1392)
);

INVx2_ASAP7_75t_SL g1393 ( 
.A(n_1381),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1378),
.Y(n_1394)
);

AOI322xp5_ASAP7_75t_L g1395 ( 
.A1(n_1383),
.A2(n_1367),
.A3(n_1368),
.B1(n_1347),
.B2(n_1259),
.C1(n_1282),
.C2(n_1337),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1378),
.A2(n_1350),
.B1(n_1340),
.B2(n_1325),
.Y(n_1396)
);

AO22x1_ASAP7_75t_L g1397 ( 
.A1(n_1385),
.A2(n_1306),
.B1(n_1340),
.B2(n_1343),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1382),
.B(n_1347),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1382),
.B(n_1347),
.Y(n_1399)
);

AOI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1372),
.A2(n_1348),
.B1(n_1337),
.B2(n_1335),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1376),
.Y(n_1401)
);

INVxp67_ASAP7_75t_L g1402 ( 
.A(n_1376),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1385),
.B(n_1348),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1384),
.B(n_1339),
.Y(n_1404)
);

AOI322xp5_ASAP7_75t_L g1405 ( 
.A1(n_1385),
.A2(n_1337),
.A3(n_1335),
.B1(n_1348),
.B2(n_1327),
.C1(n_1328),
.C2(n_1330),
.Y(n_1405)
);

XOR2x2_ASAP7_75t_L g1406 ( 
.A(n_1381),
.B(n_1151),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1395),
.A2(n_1199),
.B(n_1169),
.C(n_1218),
.Y(n_1407)
);

OAI21xp5_ASAP7_75t_SL g1408 ( 
.A1(n_1388),
.A2(n_1212),
.B(n_1343),
.Y(n_1408)
);

AOI221xp5_ASAP7_75t_L g1409 ( 
.A1(n_1397),
.A2(n_1386),
.B1(n_1373),
.B2(n_1379),
.C(n_1375),
.Y(n_1409)
);

OAI321xp33_ASAP7_75t_L g1410 ( 
.A1(n_1392),
.A2(n_1301),
.A3(n_1346),
.B1(n_1339),
.B2(n_1300),
.C(n_1252),
.Y(n_1410)
);

A2O1A1Ixp33_ASAP7_75t_L g1411 ( 
.A1(n_1405),
.A2(n_1298),
.B(n_1289),
.C(n_1346),
.Y(n_1411)
);

INVx1_ASAP7_75t_SL g1412 ( 
.A(n_1406),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1401),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1403),
.B(n_1326),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1390),
.Y(n_1415)
);

AOI32xp33_ASAP7_75t_L g1416 ( 
.A1(n_1396),
.A2(n_1346),
.A3(n_1326),
.B1(n_1333),
.B2(n_1298),
.Y(n_1416)
);

AOI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1406),
.A2(n_1326),
.B1(n_1333),
.B2(n_1335),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1394),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1414),
.B(n_1398),
.Y(n_1419)
);

AOI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1418),
.A2(n_1393),
.B(n_1391),
.Y(n_1420)
);

AOI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1412),
.A2(n_1389),
.B1(n_1393),
.B2(n_1400),
.Y(n_1421)
);

AND4x1_ASAP7_75t_L g1422 ( 
.A(n_1407),
.B(n_1389),
.C(n_1240),
.D(n_1239),
.Y(n_1422)
);

OAI221xp5_ASAP7_75t_L g1423 ( 
.A1(n_1408),
.A2(n_1402),
.B1(n_1404),
.B2(n_1380),
.C(n_1333),
.Y(n_1423)
);

AOI221xp5_ASAP7_75t_L g1424 ( 
.A1(n_1410),
.A2(n_1402),
.B1(n_1399),
.B2(n_1351),
.C(n_1366),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_1417),
.Y(n_1425)
);

AOI222xp33_ASAP7_75t_L g1426 ( 
.A1(n_1409),
.A2(n_1284),
.B1(n_1365),
.B2(n_1364),
.C1(n_1360),
.C2(n_1359),
.Y(n_1426)
);

AOI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1407),
.A2(n_1333),
.B1(n_1326),
.B2(n_1380),
.Y(n_1427)
);

AOI211xp5_ASAP7_75t_SL g1428 ( 
.A1(n_1409),
.A2(n_1199),
.B(n_1311),
.C(n_1279),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1411),
.A2(n_1290),
.B(n_1287),
.Y(n_1429)
);

AOI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1415),
.A2(n_1333),
.B1(n_1380),
.B2(n_1312),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1413),
.B(n_1416),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1422),
.B(n_1239),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1426),
.B(n_1358),
.Y(n_1433)
);

NAND4xp25_ASAP7_75t_L g1434 ( 
.A(n_1428),
.B(n_1157),
.C(n_1217),
.D(n_1174),
.Y(n_1434)
);

AOI211x1_ASAP7_75t_SL g1435 ( 
.A1(n_1431),
.A2(n_1189),
.B(n_1279),
.C(n_1310),
.Y(n_1435)
);

NAND3xp33_ASAP7_75t_L g1436 ( 
.A(n_1424),
.B(n_1427),
.C(n_1421),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1425),
.Y(n_1437)
);

O2A1O1Ixp33_ASAP7_75t_L g1438 ( 
.A1(n_1423),
.A2(n_1213),
.B(n_1263),
.C(n_1225),
.Y(n_1438)
);

AND4x1_ASAP7_75t_L g1439 ( 
.A(n_1429),
.B(n_1160),
.C(n_1221),
.D(n_1157),
.Y(n_1439)
);

NAND4xp25_ASAP7_75t_L g1440 ( 
.A(n_1429),
.B(n_1217),
.C(n_1214),
.D(n_1174),
.Y(n_1440)
);

AOI31xp33_ASAP7_75t_L g1441 ( 
.A1(n_1432),
.A2(n_1160),
.A3(n_1430),
.B(n_1221),
.Y(n_1441)
);

NAND4xp75_ASAP7_75t_L g1442 ( 
.A(n_1433),
.B(n_1223),
.C(n_1210),
.D(n_1419),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1437),
.B(n_1420),
.Y(n_1443)
);

NOR3xp33_ASAP7_75t_L g1444 ( 
.A(n_1436),
.B(n_1224),
.C(n_1214),
.Y(n_1444)
);

OR2x6_ASAP7_75t_L g1445 ( 
.A(n_1439),
.B(n_1227),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_1440),
.B(n_1227),
.Y(n_1446)
);

XOR2xp5_ASAP7_75t_L g1447 ( 
.A(n_1434),
.B(n_1215),
.Y(n_1447)
);

NOR3x1_ASAP7_75t_L g1448 ( 
.A(n_1435),
.B(n_1301),
.C(n_1292),
.Y(n_1448)
);

NOR2x1_ASAP7_75t_L g1449 ( 
.A(n_1438),
.B(n_1216),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1433),
.Y(n_1450)
);

NAND3xp33_ASAP7_75t_SL g1451 ( 
.A(n_1443),
.B(n_1201),
.C(n_1268),
.Y(n_1451)
);

NAND4xp75_ASAP7_75t_L g1452 ( 
.A(n_1448),
.B(n_1186),
.C(n_1200),
.D(n_1284),
.Y(n_1452)
);

NAND4xp75_ASAP7_75t_L g1453 ( 
.A(n_1450),
.B(n_1449),
.C(n_1446),
.D(n_1444),
.Y(n_1453)
);

AND3x4_ASAP7_75t_L g1454 ( 
.A(n_1442),
.B(n_1298),
.C(n_1196),
.Y(n_1454)
);

INVxp33_ASAP7_75t_L g1455 ( 
.A(n_1447),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1445),
.Y(n_1456)
);

NOR4xp75_ASAP7_75t_SL g1457 ( 
.A(n_1441),
.B(n_1264),
.C(n_1310),
.D(n_1292),
.Y(n_1457)
);

NAND4xp75_ASAP7_75t_L g1458 ( 
.A(n_1443),
.B(n_1186),
.C(n_1206),
.D(n_1195),
.Y(n_1458)
);

INVxp67_ASAP7_75t_SL g1459 ( 
.A(n_1455),
.Y(n_1459)
);

NAND2xp33_ASAP7_75t_L g1460 ( 
.A(n_1456),
.B(n_1273),
.Y(n_1460)
);

OAI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1453),
.A2(n_1206),
.B(n_1283),
.Y(n_1461)
);

NOR2x1p5_ASAP7_75t_L g1462 ( 
.A(n_1451),
.B(n_1273),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1459),
.Y(n_1463)
);

OAI21xp5_ASAP7_75t_SL g1464 ( 
.A1(n_1461),
.A2(n_1457),
.B(n_1454),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1463),
.A2(n_1460),
.B(n_1457),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1465),
.A2(n_1464),
.B1(n_1458),
.B2(n_1462),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1466),
.B(n_1452),
.Y(n_1467)
);

OAI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1467),
.A2(n_1216),
.B(n_1203),
.Y(n_1468)
);

OR2x6_ASAP7_75t_L g1469 ( 
.A(n_1468),
.B(n_1227),
.Y(n_1469)
);

AO21x2_ASAP7_75t_L g1470 ( 
.A1(n_1469),
.A2(n_1182),
.B(n_1181),
.Y(n_1470)
);


endmodule