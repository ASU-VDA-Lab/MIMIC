module real_aes_7259_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_673;
wire n_386;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_504;
wire n_455;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_691;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_681;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_0), .Y(n_428) );
CKINVDCx20_ASAP7_75t_R g660 ( .A(n_1), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_2), .A2(n_12), .B1(n_366), .B2(n_551), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_3), .A2(n_137), .B1(n_283), .B2(n_304), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_4), .B(n_477), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_5), .A2(n_42), .B1(n_328), .B2(n_329), .Y(n_327) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_6), .Y(n_547) );
INVx1_ASAP7_75t_L g615 ( .A(n_7), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g276 ( .A1(n_8), .A2(n_189), .B1(n_277), .B2(n_282), .Y(n_276) );
CKINVDCx20_ASAP7_75t_R g306 ( .A(n_9), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_10), .B(n_619), .Y(n_618) );
AOI22xp33_ASAP7_75t_SL g400 ( .A1(n_11), .A2(n_78), .B1(n_282), .B2(n_304), .Y(n_400) );
AOI22xp33_ASAP7_75t_SL g483 ( .A1(n_13), .A2(n_47), .B1(n_484), .B2(n_485), .Y(n_483) );
AOI22xp33_ASAP7_75t_SL g375 ( .A1(n_14), .A2(n_180), .B1(n_376), .B2(n_377), .Y(n_375) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_15), .Y(n_424) );
INVx1_ASAP7_75t_L g683 ( .A(n_16), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_17), .A2(n_219), .B1(n_332), .B2(n_359), .Y(n_478) );
INVx1_ASAP7_75t_L g337 ( .A(n_18), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_19), .A2(n_59), .B1(n_367), .B2(n_510), .Y(n_509) );
AO22x2_ASAP7_75t_L g252 ( .A1(n_20), .A2(n_64), .B1(n_243), .B2(n_248), .Y(n_252) );
INVx1_ASAP7_75t_L g646 ( .A(n_20), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_21), .A2(n_120), .B1(n_238), .B2(n_253), .Y(n_237) );
AOI22xp33_ASAP7_75t_SL g364 ( .A1(n_22), .A2(n_26), .B1(n_365), .B2(n_366), .Y(n_364) );
AOI222xp33_ASAP7_75t_L g408 ( .A1(n_23), .A2(n_77), .B1(n_97), .B2(n_348), .C1(n_409), .C2(n_410), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g631 ( .A(n_24), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_25), .A2(n_185), .B1(n_403), .B2(n_404), .Y(n_402) );
INVx1_ASAP7_75t_L g605 ( .A(n_27), .Y(n_605) );
AOI222xp33_ASAP7_75t_L g296 ( .A1(n_28), .A2(n_70), .B1(n_201), .B2(n_297), .C1(n_300), .C2(n_303), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_29), .A2(n_149), .B1(n_300), .B2(n_339), .Y(n_338) );
AOI22xp33_ASAP7_75t_SL g357 ( .A1(n_30), .A2(n_46), .B1(n_358), .B2(n_359), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g318 ( .A1(n_31), .A2(n_38), .B1(n_319), .B2(n_320), .Y(n_318) );
AOI22xp5_ASAP7_75t_L g310 ( .A1(n_32), .A2(n_169), .B1(n_239), .B2(n_288), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_33), .A2(n_125), .B1(n_367), .B2(n_390), .Y(n_389) );
AO22x2_ASAP7_75t_L g250 ( .A1(n_34), .A2(n_66), .B1(n_243), .B2(n_244), .Y(n_250) );
INVx1_ASAP7_75t_L g647 ( .A(n_34), .Y(n_647) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_35), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_36), .A2(n_102), .B1(n_379), .B2(n_630), .Y(n_629) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_37), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_39), .A2(n_115), .B1(n_484), .B2(n_485), .Y(n_674) );
INVx1_ASAP7_75t_L g517 ( .A(n_40), .Y(n_517) );
AOI22xp5_ASAP7_75t_SL g311 ( .A1(n_41), .A2(n_208), .B1(n_312), .B2(n_314), .Y(n_311) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_43), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_44), .A2(n_92), .B1(n_379), .B2(n_673), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_45), .A2(n_171), .B1(n_421), .B2(n_422), .Y(n_420) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_48), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_49), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_50), .A2(n_202), .B1(n_332), .B2(n_333), .Y(n_331) );
AOI22xp33_ASAP7_75t_SL g616 ( .A1(n_51), .A2(n_213), .B1(n_300), .B2(n_351), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_52), .B(n_361), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_53), .A2(n_69), .B1(n_514), .B2(n_583), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_54), .A2(n_127), .B1(n_406), .B2(n_407), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_55), .B(n_329), .Y(n_475) );
INVx1_ASAP7_75t_L g462 ( .A(n_56), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_57), .A2(n_150), .B1(n_323), .B2(n_510), .Y(n_569) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_58), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_60), .A2(n_124), .B1(n_426), .B2(n_514), .Y(n_513) );
AOI22xp33_ASAP7_75t_SL g480 ( .A1(n_61), .A2(n_90), .B1(n_259), .B2(n_481), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_62), .A2(n_207), .B1(n_361), .B2(n_362), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_63), .A2(n_215), .B1(n_270), .B2(n_275), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_65), .A2(n_114), .B1(n_315), .B2(n_421), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_67), .A2(n_210), .B1(n_259), .B2(n_264), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g322 ( .A1(n_68), .A2(n_168), .B1(n_323), .B2(n_325), .Y(n_322) );
AND2x2_ASAP7_75t_L g229 ( .A(n_71), .B(n_230), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_72), .A2(n_98), .B1(n_373), .B2(n_403), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g355 ( .A(n_73), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_74), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g226 ( .A(n_75), .Y(n_226) );
INVx1_ASAP7_75t_L g340 ( .A(n_76), .Y(n_340) );
AOI22xp33_ASAP7_75t_SL g372 ( .A1(n_79), .A2(n_214), .B1(n_290), .B2(n_373), .Y(n_372) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_80), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_81), .A2(n_116), .B1(n_426), .B2(n_628), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_82), .A2(n_136), .B1(n_293), .B2(n_295), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_83), .A2(n_93), .B1(n_288), .B2(n_290), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_84), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_85), .Y(n_497) );
INVx1_ASAP7_75t_L g607 ( .A(n_86), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_87), .B(n_354), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_88), .A2(n_131), .B1(n_277), .B2(n_300), .Y(n_502) );
AOI222xp33_ASAP7_75t_L g559 ( .A1(n_89), .A2(n_101), .B1(n_176), .B2(n_453), .C1(n_560), .C2(n_561), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_91), .Y(n_543) );
INVx1_ASAP7_75t_L g601 ( .A(n_94), .Y(n_601) );
CKINVDCx20_ASAP7_75t_R g696 ( .A(n_95), .Y(n_696) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_96), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_99), .Y(n_703) );
AO22x2_ASAP7_75t_L g526 ( .A1(n_100), .A2(n_527), .B1(n_562), .B2(n_563), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_100), .Y(n_562) );
AOI22xp33_ASAP7_75t_SL g368 ( .A1(n_103), .A2(n_198), .B1(n_314), .B2(n_369), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_104), .A2(n_107), .B1(n_510), .B2(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g603 ( .A(n_105), .Y(n_603) );
CKINVDCx20_ASAP7_75t_R g349 ( .A(n_106), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_108), .A2(n_133), .B1(n_571), .B2(n_572), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_109), .B(n_453), .Y(n_452) );
AOI222xp33_ASAP7_75t_L g608 ( .A1(n_110), .A2(n_147), .B1(n_154), .B2(n_277), .C1(n_298), .C2(n_354), .Y(n_608) );
AOI221xp5_ASAP7_75t_L g553 ( .A1(n_111), .A2(n_221), .B1(n_362), .B2(n_554), .C(n_555), .Y(n_553) );
AOI222xp33_ASAP7_75t_L g584 ( .A1(n_112), .A2(n_138), .B1(n_173), .B2(n_298), .C1(n_351), .C2(n_585), .Y(n_584) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_113), .Y(n_698) );
AOI22xp33_ASAP7_75t_SL g490 ( .A1(n_117), .A2(n_151), .B1(n_325), .B2(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g230 ( .A(n_118), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_119), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_121), .A2(n_204), .B1(n_392), .B2(n_393), .Y(n_391) );
CKINVDCx20_ASAP7_75t_R g655 ( .A(n_122), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_123), .A2(n_177), .B1(n_404), .B2(n_436), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_126), .A2(n_190), .B1(n_359), .B2(n_576), .Y(n_575) );
AND2x6_ASAP7_75t_L g225 ( .A(n_128), .B(n_226), .Y(n_225) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_128), .Y(n_640) );
AO22x2_ASAP7_75t_L g242 ( .A1(n_129), .A2(n_184), .B1(n_243), .B2(n_244), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_130), .A2(n_211), .B1(n_572), .B2(n_592), .Y(n_591) );
AOI22xp33_ASAP7_75t_SL g470 ( .A1(n_132), .A2(n_163), .B1(n_354), .B2(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_134), .B(n_270), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_135), .A2(n_183), .B1(n_404), .B2(n_516), .Y(n_515) );
AOI22xp33_ASAP7_75t_SL g487 ( .A1(n_139), .A2(n_205), .B1(n_319), .B2(n_488), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_140), .Y(n_557) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_141), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_142), .A2(n_216), .B1(n_390), .B2(n_580), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_143), .A2(n_200), .B1(n_359), .B2(n_576), .Y(n_709) );
INVx1_ASAP7_75t_L g595 ( .A(n_144), .Y(n_595) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_145), .A2(n_223), .B(n_231), .C(n_648), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_146), .B(n_707), .Y(n_706) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_148), .Y(n_412) );
INVx1_ASAP7_75t_L g609 ( .A(n_152), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_153), .A2(n_199), .B1(n_315), .B2(n_692), .Y(n_691) );
AO22x2_ASAP7_75t_L g247 ( .A1(n_155), .A2(n_191), .B1(n_243), .B2(n_248), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_156), .Y(n_443) );
AOI22xp33_ASAP7_75t_SL g624 ( .A1(n_157), .A2(n_196), .B1(n_516), .B2(n_580), .Y(n_624) );
XOR2x2_ASAP7_75t_L g566 ( .A(n_158), .B(n_567), .Y(n_566) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_159), .Y(n_665) );
AOI22xp33_ASAP7_75t_SL g704 ( .A1(n_160), .A2(n_174), .B1(n_473), .B2(n_585), .Y(n_704) );
AOI22xp33_ASAP7_75t_SL g625 ( .A1(n_161), .A2(n_162), .B1(n_264), .B2(n_421), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g666 ( .A(n_164), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_165), .A2(n_197), .B1(n_303), .B2(n_576), .Y(n_598) );
INVx1_ASAP7_75t_L g506 ( .A(n_166), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_167), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g662 ( .A(n_170), .Y(n_662) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_172), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_175), .B(n_597), .Y(n_596) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_178), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_179), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_181), .Y(n_455) );
XOR2x2_ASAP7_75t_L g465 ( .A(n_182), .B(n_466), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_184), .B(n_645), .Y(n_644) );
CKINVDCx20_ASAP7_75t_R g395 ( .A(n_186), .Y(n_395) );
CKINVDCx20_ASAP7_75t_R g556 ( .A(n_187), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_188), .A2(n_193), .B1(n_582), .B2(n_583), .Y(n_581) );
INVx1_ASAP7_75t_L g643 ( .A(n_191), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_192), .A2(n_218), .B1(n_329), .B2(n_554), .Y(n_574) );
INVx1_ASAP7_75t_L g469 ( .A(n_194), .Y(n_469) );
OA22x2_ASAP7_75t_L g342 ( .A1(n_195), .A2(n_343), .B1(n_344), .B2(n_380), .Y(n_342) );
CKINVDCx20_ASAP7_75t_R g343 ( .A(n_195), .Y(n_343) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_203), .Y(n_352) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_206), .A2(n_650), .B1(n_675), .B2(n_676), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_206), .Y(n_675) );
INVx1_ASAP7_75t_L g243 ( .A(n_209), .Y(n_243) );
INVx1_ASAP7_75t_L g245 ( .A(n_209), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g653 ( .A(n_212), .Y(n_653) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_217), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_220), .Y(n_498) );
INVx1_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_227), .Y(n_224) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_226), .Y(n_639) );
OAI21xp5_ASAP7_75t_L g681 ( .A1(n_227), .A2(n_638), .B(n_682), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_228), .Y(n_227) );
INVxp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AOI221xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_521), .B1(n_633), .B2(n_634), .C(n_635), .Y(n_231) );
INVx1_ASAP7_75t_L g633 ( .A(n_232), .Y(n_633) );
XNOR2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_341), .Y(n_232) );
XNOR2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_307), .Y(n_233) );
XOR2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_306), .Y(n_234) );
NAND4xp75_ASAP7_75t_L g235 ( .A(n_236), .B(n_268), .C(n_286), .D(n_296), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_258), .Y(n_236) );
BUFx3_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
BUFx3_ASAP7_75t_L g365 ( .A(n_239), .Y(n_365) );
BUFx3_ASAP7_75t_L g407 ( .A(n_239), .Y(n_407) );
INVx6_ASAP7_75t_L g427 ( .A(n_239), .Y(n_427) );
AND2x4_ASAP7_75t_L g239 ( .A(n_240), .B(n_249), .Y(n_239) );
AND2x2_ASAP7_75t_L g294 ( .A(n_240), .B(n_261), .Y(n_294) );
AND2x6_ASAP7_75t_L g295 ( .A(n_240), .B(n_273), .Y(n_295) );
AND2x6_ASAP7_75t_L g298 ( .A(n_240), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_246), .Y(n_240) );
AND2x2_ASAP7_75t_L g263 ( .A(n_241), .B(n_247), .Y(n_263) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g256 ( .A(n_242), .B(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_242), .B(n_247), .Y(n_267) );
AND2x2_ASAP7_75t_L g281 ( .A(n_242), .B(n_252), .Y(n_281) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g248 ( .A(n_245), .Y(n_248) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g257 ( .A(n_247), .Y(n_257) );
INVx1_ASAP7_75t_L g280 ( .A(n_247), .Y(n_280) );
AND2x2_ASAP7_75t_L g255 ( .A(n_249), .B(n_256), .Y(n_255) );
AND2x6_ASAP7_75t_L g275 ( .A(n_249), .B(n_263), .Y(n_275) );
NAND2x1p5_ASAP7_75t_L g398 ( .A(n_249), .B(n_263), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_249), .B(n_256), .Y(n_538) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
INVx2_ASAP7_75t_L g262 ( .A(n_250), .Y(n_262) );
OR2x2_ASAP7_75t_L g274 ( .A(n_250), .B(n_251), .Y(n_274) );
INVx1_ASAP7_75t_L g285 ( .A(n_250), .Y(n_285) );
AND2x2_ASAP7_75t_L g299 ( .A(n_250), .B(n_252), .Y(n_299) );
AND2x2_ASAP7_75t_L g261 ( .A(n_251), .B(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
BUFx2_ASAP7_75t_L g484 ( .A(n_253), .Y(n_484) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_253), .Y(n_571) );
INVx5_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx4_ASAP7_75t_L g313 ( .A(n_254), .Y(n_313) );
INVx1_ASAP7_75t_L g370 ( .A(n_254), .Y(n_370) );
INVx3_ASAP7_75t_L g392 ( .A(n_254), .Y(n_392) );
INVx2_ASAP7_75t_L g421 ( .A(n_254), .Y(n_421) );
BUFx3_ASAP7_75t_L g593 ( .A(n_254), .Y(n_593) );
INVx8_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g289 ( .A(n_256), .B(n_261), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_256), .B(n_261), .Y(n_431) );
INVx1_ASAP7_75t_L g305 ( .A(n_257), .Y(n_305) );
INVx4_ASAP7_75t_L g324 ( .A(n_259), .Y(n_324) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
BUFx3_ASAP7_75t_L g379 ( .A(n_260), .Y(n_379) );
BUFx3_ASAP7_75t_L g404 ( .A(n_260), .Y(n_404) );
AND2x4_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
AND2x4_ASAP7_75t_L g291 ( .A(n_261), .B(n_266), .Y(n_291) );
INVx1_ASAP7_75t_L g265 ( .A(n_262), .Y(n_265) );
AND2x2_ASAP7_75t_L g279 ( .A(n_262), .B(n_280), .Y(n_279) );
AND2x4_ASAP7_75t_L g272 ( .A(n_263), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g458 ( .A(n_263), .Y(n_458) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
NAND2x1p5_ASAP7_75t_L g442 ( .A(n_265), .B(n_281), .Y(n_442) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OR2x6_ASAP7_75t_L g316 ( .A(n_267), .B(n_285), .Y(n_316) );
AND2x2_ASAP7_75t_SL g268 ( .A(n_269), .B(n_276), .Y(n_268) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_270), .Y(n_554) );
INVx5_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g328 ( .A(n_271), .Y(n_328) );
INVx2_ASAP7_75t_L g361 ( .A(n_271), .Y(n_361) );
INVx2_ASAP7_75t_L g477 ( .A(n_271), .Y(n_477) );
INVx4_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g457 ( .A(n_274), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_SL g330 ( .A(n_275), .Y(n_330) );
BUFx2_ASAP7_75t_L g362 ( .A(n_275), .Y(n_362) );
BUFx4f_ASAP7_75t_L g619 ( .A(n_275), .Y(n_619) );
BUFx2_ASAP7_75t_L g707 ( .A(n_275), .Y(n_707) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_277), .Y(n_409) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
BUFx2_ASAP7_75t_L g339 ( .A(n_278), .Y(n_339) );
BUFx4f_ASAP7_75t_SL g351 ( .A(n_278), .Y(n_351) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_278), .Y(n_453) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_278), .Y(n_473) );
AND2x4_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
INVx1_ASAP7_75t_L g302 ( .A(n_280), .Y(n_302) );
AND2x4_ASAP7_75t_L g283 ( .A(n_281), .B(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_L g301 ( .A(n_281), .B(n_302), .Y(n_301) );
BUFx3_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx2_ASAP7_75t_L g332 ( .A(n_283), .Y(n_332) );
BUFx2_ASAP7_75t_L g358 ( .A(n_283), .Y(n_358) );
INVx1_ASAP7_75t_L g577 ( .A(n_283), .Y(n_577) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_292), .Y(n_286) );
INVx1_ASAP7_75t_L g489 ( .A(n_288), .Y(n_489) );
BUFx3_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx3_ASAP7_75t_L g367 ( .A(n_289), .Y(n_367) );
BUFx3_ASAP7_75t_L g580 ( .A(n_289), .Y(n_580) );
BUFx3_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
BUFx2_ASAP7_75t_SL g325 ( .A(n_291), .Y(n_325) );
BUFx3_ASAP7_75t_L g390 ( .A(n_291), .Y(n_390) );
BUFx2_ASAP7_75t_SL g436 ( .A(n_291), .Y(n_436) );
BUFx2_ASAP7_75t_L g516 ( .A(n_291), .Y(n_516) );
BUFx3_ASAP7_75t_L g552 ( .A(n_291), .Y(n_552) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_293), .Y(n_319) );
BUFx3_ASAP7_75t_L g376 ( .A(n_293), .Y(n_376) );
BUFx3_ASAP7_75t_L g673 ( .A(n_293), .Y(n_673) );
INVx3_ASAP7_75t_L g699 ( .A(n_293), .Y(n_699) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
BUFx2_ASAP7_75t_SL g403 ( .A(n_294), .Y(n_403) );
BUFx2_ASAP7_75t_SL g510 ( .A(n_294), .Y(n_510) );
INVx2_ASAP7_75t_L g531 ( .A(n_294), .Y(n_531) );
INVx11_ASAP7_75t_L g321 ( .A(n_295), .Y(n_321) );
INVx11_ASAP7_75t_L g374 ( .A(n_295), .Y(n_374) );
INVx3_ASAP7_75t_L g501 ( .A(n_297), .Y(n_501) );
BUFx3_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx4_ASAP7_75t_L g336 ( .A(n_298), .Y(n_336) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_298), .Y(n_659) );
AND2x4_ASAP7_75t_L g304 ( .A(n_299), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g445 ( .A(n_299), .Y(n_445) );
INVx2_ASAP7_75t_L g411 ( .A(n_300), .Y(n_411) );
BUFx4f_ASAP7_75t_SL g585 ( .A(n_300), .Y(n_585) );
BUFx12f_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_301), .Y(n_354) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_301), .Y(n_450) );
BUFx3_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_304), .Y(n_333) );
BUFx2_ASAP7_75t_SL g359 ( .A(n_304), .Y(n_359) );
INVx1_ASAP7_75t_L g446 ( .A(n_305), .Y(n_446) );
XOR2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_340), .Y(n_307) );
NOR4xp75_ASAP7_75t_L g308 ( .A(n_309), .B(n_317), .C(n_326), .D(n_334), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g309 ( .A(n_310), .B(n_311), .Y(n_309) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g693 ( .A(n_313), .Y(n_693) );
INVxp67_ASAP7_75t_L g540 ( .A(n_314), .Y(n_540) );
BUFx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
BUFx2_ASAP7_75t_L g393 ( .A(n_315), .Y(n_393) );
BUFx2_ASAP7_75t_L g485 ( .A(n_315), .Y(n_485) );
BUFx2_ASAP7_75t_L g572 ( .A(n_315), .Y(n_572) );
INVx6_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g422 ( .A(n_316), .Y(n_422) );
NAND2x1_ASAP7_75t_L g317 ( .A(n_318), .B(n_322), .Y(n_317) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_SL g406 ( .A(n_321), .Y(n_406) );
INVx4_ASAP7_75t_L g514 ( .A(n_321), .Y(n_514) );
INVx1_ASAP7_75t_L g582 ( .A(n_321), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_321), .A2(n_427), .B1(n_695), .B2(n_696), .Y(n_694) );
INVx4_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_324), .A2(n_433), .B1(n_434), .B2(n_435), .Y(n_432) );
INVx3_ASAP7_75t_L g590 ( .A(n_324), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g326 ( .A(n_327), .B(n_331), .Y(n_326) );
INVx1_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
OAI21xp5_ASAP7_75t_SL g334 ( .A1(n_335), .A2(n_337), .B(n_338), .Y(n_334) );
INVx1_ASAP7_75t_L g560 ( .A(n_335), .Y(n_560) );
BUFx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx4_ASAP7_75t_L g348 ( .A(n_336), .Y(n_348) );
OAI221xp5_ASAP7_75t_L g447 ( .A1(n_336), .A2(n_448), .B1(n_449), .B2(n_451), .C(n_452), .Y(n_447) );
OAI21xp5_ASAP7_75t_SL g702 ( .A1(n_336), .A2(n_703), .B(n_704), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_381), .B1(n_382), .B2(n_520), .Y(n_341) );
INVx1_ASAP7_75t_L g520 ( .A(n_342), .Y(n_520) );
INVx2_ASAP7_75t_L g380 ( .A(n_344), .Y(n_380) );
NAND3x1_ASAP7_75t_L g344 ( .A(n_345), .B(n_363), .C(n_371), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_346), .B(n_356), .Y(n_345) );
OAI222xp33_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_349), .B1(n_350), .B2(n_352), .C1(n_353), .C2(n_355), .Y(n_346) );
OAI21xp5_ASAP7_75t_SL g468 ( .A1(n_347), .A2(n_469), .B(n_470), .Y(n_468) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_357), .B(n_360), .Y(n_356) );
BUFx2_ASAP7_75t_L g597 ( .A(n_361), .Y(n_597) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_368), .Y(n_363) );
BUFx3_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_375), .Y(n_371) );
INVx1_ASAP7_75t_L g606 ( .A(n_373), .Y(n_606) );
INVx3_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_374), .A2(n_543), .B1(n_544), .B2(n_545), .Y(n_542) );
INVx4_ASAP7_75t_L g628 ( .A(n_374), .Y(n_628) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_384), .B1(n_463), .B2(n_519), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OAI22xp5_ASAP7_75t_SL g384 ( .A1(n_385), .A2(n_386), .B1(n_413), .B2(n_414), .Y(n_384) );
INVx3_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
XOR2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_412), .Y(n_386) );
NAND4xp75_ASAP7_75t_L g387 ( .A(n_388), .B(n_394), .C(n_401), .D(n_408), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_391), .Y(n_388) );
INVxp67_ASAP7_75t_L g602 ( .A(n_390), .Y(n_602) );
OA211x2_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B(n_399), .C(n_400), .Y(n_394) );
OA211x2_ASAP7_75t_L g594 ( .A1(n_396), .A2(n_595), .B(n_596), .C(n_598), .Y(n_594) );
BUFx3_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
BUFx3_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g461 ( .A(n_398), .Y(n_461) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_405), .Y(n_401) );
BUFx2_ASAP7_75t_L g534 ( .A(n_404), .Y(n_534) );
INVx1_ASAP7_75t_L g482 ( .A(n_406), .Y(n_482) );
INVx1_ASAP7_75t_L g545 ( .A(n_407), .Y(n_545) );
INVx2_ASAP7_75t_SL g661 ( .A(n_409), .Y(n_661) );
INVx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
XOR2xp5_ASAP7_75t_SL g415 ( .A(n_416), .B(n_462), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_437), .Y(n_416) );
NOR3xp33_ASAP7_75t_L g417 ( .A(n_418), .B(n_423), .C(n_432), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_425), .B1(n_428), .B2(n_429), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_425), .A2(n_605), .B1(n_606), .B2(n_607), .Y(n_604) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx3_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g491 ( .A(n_427), .Y(n_491) );
INVx2_ASAP7_75t_L g583 ( .A(n_427), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_429), .A2(n_601), .B1(n_602), .B2(n_603), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_429), .A2(n_698), .B1(n_699), .B2(n_700), .Y(n_697) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g548 ( .A(n_430), .Y(n_548) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
NOR3xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_447), .C(n_454), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_440), .B1(n_443), .B2(n_444), .Y(n_438) );
INVx3_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
INVx4_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx3_ASAP7_75t_L g505 ( .A(n_442), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_442), .A2(n_558), .B1(n_665), .B2(n_666), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_444), .A2(n_504), .B1(n_505), .B2(n_506), .Y(n_503) );
BUFx2_ASAP7_75t_L g558 ( .A(n_444), .Y(n_558) );
OR2x6_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
BUFx3_ASAP7_75t_L g561 ( .A(n_450), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_456), .B1(n_459), .B2(n_460), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_456), .A2(n_460), .B1(n_497), .B2(n_498), .Y(n_496) );
BUFx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_457), .Y(n_654) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_SL g656 ( .A(n_461), .Y(n_656) );
INVx1_ASAP7_75t_L g519 ( .A(n_463), .Y(n_519) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_492), .B1(n_493), .B2(n_518), .Y(n_464) );
INVx2_ASAP7_75t_L g518 ( .A(n_465), .Y(n_518) );
NAND3x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_479), .C(n_486), .Y(n_466) );
NOR2x1_ASAP7_75t_SL g467 ( .A(n_468), .B(n_474), .Y(n_467) );
INVx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx4_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NAND3xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .C(n_478), .Y(n_474) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_483), .Y(n_479) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_490), .Y(n_486) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_SL g492 ( .A(n_493), .Y(n_492) );
XOR2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_517), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_507), .Y(n_494) );
NOR3xp33_ASAP7_75t_L g495 ( .A(n_496), .B(n_499), .C(n_503), .Y(n_495) );
OAI21xp33_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_501), .B(n_502), .Y(n_499) );
OAI21xp5_ASAP7_75t_SL g614 ( .A1(n_501), .A2(n_615), .B(n_616), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_505), .A2(n_556), .B1(n_557), .B2(n_558), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_508), .B(n_512), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_511), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_515), .Y(n_512) );
INVx1_ASAP7_75t_L g634 ( .A(n_521), .Y(n_634) );
AOI22xp5_ASAP7_75t_SL g521 ( .A1(n_522), .A2(n_610), .B1(n_611), .B2(n_632), .Y(n_521) );
INVx1_ASAP7_75t_L g632 ( .A(n_522), .Y(n_632) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_526), .B1(n_564), .B2(n_565), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g563 ( .A(n_527), .Y(n_563) );
AND4x1_ASAP7_75t_L g527 ( .A(n_528), .B(n_541), .C(n_553), .D(n_559), .Y(n_527) );
NOR2xp33_ASAP7_75t_SL g528 ( .A(n_529), .B(n_535), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B1(n_532), .B2(n_533), .Y(n_529) );
INVx3_ASAP7_75t_L g630 ( .A(n_531), .Y(n_630) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_537), .B1(n_539), .B2(n_540), .Y(n_535) );
BUFx2_ASAP7_75t_R g537 ( .A(n_538), .Y(n_537) );
NOR2xp33_ASAP7_75t_SL g541 ( .A(n_542), .B(n_546), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B1(n_549), .B2(n_550), .Y(n_546) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
XOR2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_586), .Y(n_565) );
NAND4xp75_ASAP7_75t_L g567 ( .A(n_568), .B(n_573), .C(n_578), .D(n_584), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
AND2x2_ASAP7_75t_SL g573 ( .A(n_574), .B(n_575), .Y(n_573) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
XOR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_609), .Y(n_586) );
NAND4xp75_ASAP7_75t_L g587 ( .A(n_588), .B(n_594), .C(n_599), .D(n_608), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .Y(n_588) );
INVx3_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_600), .B(n_604), .Y(n_599) );
INVx3_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
XOR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_631), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g612 ( .A(n_613), .B(n_622), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_614), .B(n_617), .Y(n_613) );
NAND3xp33_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .C(n_621), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_626), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
INVx1_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
NOR2x1_ASAP7_75t_L g636 ( .A(n_637), .B(n_641), .Y(n_636) );
OR2x2_ASAP7_75t_SL g712 ( .A(n_637), .B(n_642), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_639), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_639), .B(n_679), .Y(n_682) );
CKINVDCx16_ASAP7_75t_R g679 ( .A(n_640), .Y(n_679) );
CKINVDCx20_ASAP7_75t_R g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
OAI322xp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_677), .A3(n_678), .B1(n_680), .B2(n_683), .C1(n_684), .C2(n_710), .Y(n_648) );
INVx1_ASAP7_75t_L g676 ( .A(n_650), .Y(n_676) );
AND2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_667), .Y(n_650) );
NOR3xp33_ASAP7_75t_L g651 ( .A(n_652), .B(n_657), .C(n_664), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_654), .B1(n_655), .B2(n_656), .Y(n_652) );
OAI221xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_660), .B1(n_661), .B2(n_662), .C(n_663), .Y(n_657) );
INVx2_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_668), .B(n_671), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_674), .Y(n_671) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
CKINVDCx16_ASAP7_75t_R g680 ( .A(n_681), .Y(n_680) );
XOR2x2_ASAP7_75t_L g686 ( .A(n_683), .B(n_687), .Y(n_686) );
CKINVDCx16_ASAP7_75t_R g684 ( .A(n_685), .Y(n_684) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_SL g687 ( .A(n_688), .B(n_701), .Y(n_687) );
NOR3xp33_ASAP7_75t_L g688 ( .A(n_689), .B(n_694), .C(n_697), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
INVx3_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_702), .B(n_705), .Y(n_701) );
NAND3xp33_ASAP7_75t_L g705 ( .A(n_706), .B(n_708), .C(n_709), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_711), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_712), .Y(n_711) );
endmodule