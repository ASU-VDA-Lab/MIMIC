module fake_ariane_25_n_2136 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_499, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_522, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_528, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_511, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_234, n_492, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_30, n_494, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_127, n_531, n_2136);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_499;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_522;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_528;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_234;
input n_492;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_127;
input n_531;

output n_2136;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_1383;
wire n_603;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_690;
wire n_1109;
wire n_1430;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_1682;
wire n_1836;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_813;
wire n_1985;
wire n_995;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_559;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_661;
wire n_2098;
wire n_1751;
wire n_1917;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_1112;
wire n_1159;
wire n_700;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2116;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_1432;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_696;
wire n_1442;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_2087;
wire n_931;
wire n_669;
wire n_1491;
wire n_619;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_1340;
wire n_1240;
wire n_1087;
wire n_632;
wire n_650;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_976;
wire n_712;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_1578;
wire n_1455;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_706;
wire n_2120;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_552;
wire n_670;
wire n_1826;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_1899;
wire n_1467;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_677;
wire n_604;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_1015;
wire n_545;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_1156;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_957;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_1005;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_1708;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_1281;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1733;
wire n_1476;
wire n_1524;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_1165;
wire n_1641;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_1038;
wire n_1978;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_2014;
wire n_975;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_1775;
wire n_908;
wire n_788;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_1537;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_917;
wire n_1271;
wire n_2096;
wire n_1530;
wire n_631;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_1813;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_1344;
wire n_1390;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_1150;
wire n_977;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_1136;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_954;
wire n_596;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_574;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_1063;
wire n_991;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_937;
wire n_1474;
wire n_2081;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_548;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_849;
wire n_2095;
wire n_1820;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_573;
wire n_796;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_147),
.Y(n_540)
);

BUFx2_ASAP7_75t_SL g541 ( 
.A(n_354),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_517),
.Y(n_542)
);

BUFx10_ASAP7_75t_L g543 ( 
.A(n_178),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_468),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_363),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_153),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_101),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_223),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_344),
.Y(n_549)
);

INVx1_ASAP7_75t_SL g550 ( 
.A(n_125),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_103),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_326),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_32),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_461),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_200),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_92),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_71),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_248),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_533),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_198),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_280),
.Y(n_561)
);

BUFx2_ASAP7_75t_SL g562 ( 
.A(n_222),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_272),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_510),
.Y(n_564)
);

BUFx8_ASAP7_75t_SL g565 ( 
.A(n_189),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_478),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_482),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_519),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_95),
.Y(n_569)
);

CKINVDCx16_ASAP7_75t_R g570 ( 
.A(n_39),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_57),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_509),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_104),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_407),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_294),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_373),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_3),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_347),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_251),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_507),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_531),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_323),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_480),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_431),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_227),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_52),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_371),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_515),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_170),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_83),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_31),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_177),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_194),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_532),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_41),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_303),
.Y(n_596)
);

CKINVDCx16_ASAP7_75t_R g597 ( 
.A(n_276),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_316),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_415),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_378),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_360),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_295),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_278),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_529),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_504),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_255),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_486),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_228),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_293),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_51),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_21),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_457),
.Y(n_612)
);

CKINVDCx16_ASAP7_75t_R g613 ( 
.A(n_1),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_79),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_29),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_534),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_479),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_254),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_435),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_122),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_539),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_14),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_105),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_506),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_387),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_155),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_390),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_300),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_19),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_352),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_249),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_325),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_1),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_116),
.Y(n_634)
);

INVxp33_ASAP7_75t_L g635 ( 
.A(n_398),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_204),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_113),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_301),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_423),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_69),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_257),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_481),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_92),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_50),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_424),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_403),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_124),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_289),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_477),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_343),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_52),
.Y(n_651)
);

BUFx10_ASAP7_75t_L g652 ( 
.A(n_466),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_157),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_456),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_155),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_530),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_432),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_71),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_154),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_513),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_0),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_508),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_164),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_452),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_512),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_143),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_314),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_112),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_45),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g670 ( 
.A(n_217),
.Y(n_670)
);

BUFx10_ASAP7_75t_L g671 ( 
.A(n_537),
.Y(n_671)
);

CKINVDCx20_ASAP7_75t_R g672 ( 
.A(n_88),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_74),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_238),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_310),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_404),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_332),
.Y(n_677)
);

INVxp67_ASAP7_75t_SL g678 ( 
.A(n_280),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_32),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_36),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_224),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_458),
.Y(n_682)
);

CKINVDCx14_ASAP7_75t_R g683 ( 
.A(n_397),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_180),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_22),
.Y(n_685)
);

BUFx5_ASAP7_75t_L g686 ( 
.A(n_427),
.Y(n_686)
);

INVxp67_ASAP7_75t_L g687 ( 
.A(n_448),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_455),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_329),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_236),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_72),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_10),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_75),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_243),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_490),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_183),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_511),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_78),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_523),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_204),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_505),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_462),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_119),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_7),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_368),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_476),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_472),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_212),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_400),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_272),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_250),
.Y(n_711)
);

INVx1_ASAP7_75t_SL g712 ( 
.A(n_181),
.Y(n_712)
);

BUFx10_ASAP7_75t_L g713 ( 
.A(n_182),
.Y(n_713)
);

HB1xp67_ASAP7_75t_L g714 ( 
.A(n_522),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_444),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_391),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_346),
.Y(n_717)
);

INVx1_ASAP7_75t_SL g718 ( 
.A(n_525),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_536),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_526),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_6),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_518),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_125),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_144),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_503),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_233),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_357),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_263),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_142),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_191),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_514),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_470),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_467),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_520),
.Y(n_734)
);

CKINVDCx16_ASAP7_75t_R g735 ( 
.A(n_291),
.Y(n_735)
);

BUFx5_ASAP7_75t_L g736 ( 
.A(n_535),
.Y(n_736)
);

BUFx2_ASAP7_75t_SL g737 ( 
.A(n_216),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_119),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_229),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_153),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_120),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_318),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_100),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_14),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_340),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_31),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_527),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_524),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_11),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_306),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_500),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_226),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_7),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_133),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_475),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_149),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_473),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_441),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_411),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_487),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_516),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_76),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_401),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_185),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_425),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_350),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_137),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_41),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_169),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_251),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_528),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_56),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_413),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_74),
.Y(n_774)
);

HB1xp67_ASAP7_75t_L g775 ( 
.A(n_50),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_151),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_261),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_337),
.Y(n_778)
);

CKINVDCx20_ASAP7_75t_R g779 ( 
.A(n_412),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_203),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_383),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_145),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_393),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_193),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_521),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_252),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_189),
.Y(n_787)
);

CKINVDCx20_ASAP7_75t_R g788 ( 
.A(n_202),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_224),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_127),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_150),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_140),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_420),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_56),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_133),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_283),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_166),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_317),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_44),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_379),
.Y(n_800)
);

CKINVDCx20_ASAP7_75t_R g801 ( 
.A(n_250),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_114),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_246),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_159),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_298),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_333),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_236),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_429),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_115),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_704),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_704),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_739),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_739),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_791),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_540),
.Y(n_815)
);

INVxp67_ASAP7_75t_L g816 ( 
.A(n_775),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_791),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_701),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_802),
.Y(n_819)
);

INVxp67_ASAP7_75t_SL g820 ( 
.A(n_540),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_546),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_540),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_551),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_553),
.Y(n_824)
);

CKINVDCx20_ASAP7_75t_R g825 ( 
.A(n_548),
.Y(n_825)
);

INVxp33_ASAP7_75t_SL g826 ( 
.A(n_714),
.Y(n_826)
);

CKINVDCx16_ASAP7_75t_R g827 ( 
.A(n_570),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_558),
.Y(n_828)
);

INVxp67_ASAP7_75t_SL g829 ( 
.A(n_540),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_577),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_585),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_548),
.Y(n_832)
);

CKINVDCx14_ASAP7_75t_R g833 ( 
.A(n_683),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_591),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_555),
.Y(n_835)
);

INVxp33_ASAP7_75t_SL g836 ( 
.A(n_547),
.Y(n_836)
);

CKINVDCx16_ASAP7_75t_R g837 ( 
.A(n_597),
.Y(n_837)
);

CKINVDCx20_ASAP7_75t_R g838 ( 
.A(n_555),
.Y(n_838)
);

BUFx2_ASAP7_75t_L g839 ( 
.A(n_565),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_606),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_592),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_595),
.Y(n_842)
);

INVxp33_ASAP7_75t_SL g843 ( 
.A(n_557),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_610),
.Y(n_844)
);

INVxp33_ASAP7_75t_SL g845 ( 
.A(n_560),
.Y(n_845)
);

INVxp67_ASAP7_75t_SL g846 ( 
.A(n_606),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_618),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_626),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_565),
.Y(n_849)
);

CKINVDCx20_ASAP7_75t_R g850 ( 
.A(n_670),
.Y(n_850)
);

INVxp67_ASAP7_75t_SL g851 ( 
.A(n_606),
.Y(n_851)
);

CKINVDCx20_ASAP7_75t_R g852 ( 
.A(n_670),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_631),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_636),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_637),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_640),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_647),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_648),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_679),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_684),
.Y(n_860)
);

CKINVDCx14_ASAP7_75t_R g861 ( 
.A(n_683),
.Y(n_861)
);

INVxp67_ASAP7_75t_SL g862 ( 
.A(n_606),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_685),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_698),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_613),
.Y(n_865)
);

BUFx3_ASAP7_75t_L g866 ( 
.A(n_701),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_735),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_708),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_723),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_729),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_743),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_744),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_746),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_754),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_745),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_767),
.Y(n_876)
);

INVxp67_ASAP7_75t_SL g877 ( 
.A(n_563),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_721),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_552),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_567),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_770),
.Y(n_881)
);

INVxp67_ASAP7_75t_SL g882 ( 
.A(n_563),
.Y(n_882)
);

CKINVDCx20_ASAP7_75t_R g883 ( 
.A(n_721),
.Y(n_883)
);

INVxp33_ASAP7_75t_SL g884 ( 
.A(n_561),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_772),
.Y(n_885)
);

INVxp67_ASAP7_75t_SL g886 ( 
.A(n_579),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_599),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_632),
.Y(n_888)
);

INVxp33_ASAP7_75t_SL g889 ( 
.A(n_569),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_573),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_786),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_586),
.Y(n_892)
);

CKINVDCx20_ASAP7_75t_R g893 ( 
.A(n_726),
.Y(n_893)
);

INVxp67_ASAP7_75t_SL g894 ( 
.A(n_579),
.Y(n_894)
);

INVxp33_ASAP7_75t_SL g895 ( 
.A(n_589),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_552),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_745),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_795),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_796),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_818),
.B(n_590),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_816),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_833),
.B(n_559),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_815),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_815),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_826),
.B(n_635),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_822),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_822),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_820),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_892),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_829),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_840),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_861),
.B(n_635),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_846),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_840),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_880),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_827),
.B(n_543),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_818),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_866),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_851),
.Y(n_919)
);

OAI22x1_ASAP7_75t_SL g920 ( 
.A1(n_825),
.A2(n_801),
.B1(n_726),
.B2(n_556),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_862),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_866),
.B(n_564),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_875),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_875),
.B(n_590),
.Y(n_924)
);

BUFx12f_ASAP7_75t_L g925 ( 
.A(n_849),
.Y(n_925)
);

INVx6_ASAP7_75t_L g926 ( 
.A(n_897),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_826),
.A2(n_719),
.B1(n_732),
.B2(n_646),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_821),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_897),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_823),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_890),
.B(n_836),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_867),
.A2(n_719),
.B1(n_732),
.B2(n_646),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_836),
.B(n_639),
.Y(n_933)
);

NOR2x1_ASAP7_75t_L g934 ( 
.A(n_810),
.B(n_541),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_811),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_824),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_828),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_830),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_831),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_834),
.Y(n_940)
);

CKINVDCx16_ASAP7_75t_R g941 ( 
.A(n_837),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_867),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_877),
.B(n_543),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_841),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_842),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_SL g946 ( 
.A1(n_825),
.A2(n_801),
.B1(n_571),
.B2(n_641),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_844),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_847),
.Y(n_948)
);

INVx5_ASAP7_75t_L g949 ( 
.A(n_839),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_843),
.B(n_639),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_882),
.B(n_790),
.Y(n_951)
);

BUFx8_ASAP7_75t_L g952 ( 
.A(n_848),
.Y(n_952)
);

INVx5_ASAP7_75t_L g953 ( 
.A(n_886),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_894),
.B(n_812),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_843),
.B(n_549),
.Y(n_955)
);

INVx4_ASAP7_75t_L g956 ( 
.A(n_813),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_853),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_854),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_855),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_887),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_856),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_857),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_R g963 ( 
.A(n_915),
.B(n_888),
.Y(n_963)
);

CKINVDCx16_ASAP7_75t_R g964 ( 
.A(n_941),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_R g965 ( 
.A(n_915),
.B(n_849),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_901),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_960),
.Y(n_967)
);

CKINVDCx20_ASAP7_75t_R g968 ( 
.A(n_927),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_903),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_903),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_930),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_925),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_925),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_930),
.Y(n_974)
);

BUFx10_ASAP7_75t_L g975 ( 
.A(n_931),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_904),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_952),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_952),
.Y(n_978)
);

BUFx10_ASAP7_75t_L g979 ( 
.A(n_931),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_901),
.B(n_865),
.Y(n_980)
);

CKINVDCx20_ASAP7_75t_R g981 ( 
.A(n_932),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_952),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_933),
.B(n_895),
.Y(n_983)
);

INVxp67_ASAP7_75t_L g984 ( 
.A(n_905),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_942),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_949),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_938),
.Y(n_987)
);

CKINVDCx20_ASAP7_75t_R g988 ( 
.A(n_946),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_906),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_949),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_938),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_945),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_949),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_949),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_918),
.Y(n_995)
);

CKINVDCx11_ASAP7_75t_R g996 ( 
.A(n_945),
.Y(n_996)
);

INVxp67_ASAP7_75t_L g997 ( 
.A(n_905),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_918),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_947),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_947),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_918),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_955),
.B(n_845),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_906),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_909),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_904),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_959),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_959),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_955),
.B(n_845),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_R g1009 ( 
.A(n_917),
.B(n_879),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_916),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_918),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_944),
.Y(n_1012)
);

CKINVDCx16_ASAP7_75t_R g1013 ( 
.A(n_912),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_906),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_906),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_923),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_923),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_907),
.Y(n_1018)
);

INVxp67_ASAP7_75t_L g1019 ( 
.A(n_933),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_923),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_923),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_907),
.Y(n_1022)
);

HB1xp67_ASAP7_75t_L g1023 ( 
.A(n_917),
.Y(n_1023)
);

BUFx2_ASAP7_75t_L g1024 ( 
.A(n_943),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_920),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_961),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_926),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_926),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_926),
.Y(n_1029)
);

AOI21x1_ASAP7_75t_L g1030 ( 
.A1(n_922),
.A2(n_574),
.B(n_566),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_935),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_935),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_907),
.Y(n_1033)
);

BUFx2_ASAP7_75t_L g1034 ( 
.A(n_954),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_950),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_950),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_954),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_961),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_961),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_929),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_907),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_1034),
.B(n_954),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_1031),
.B(n_884),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_SL g1044 ( 
.A(n_975),
.Y(n_1044)
);

OAI22xp33_ASAP7_75t_L g1045 ( 
.A1(n_984),
.A2(n_896),
.B1(n_879),
.B2(n_634),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_971),
.Y(n_1046)
);

AND2x4_ASAP7_75t_L g1047 ( 
.A(n_1037),
.B(n_951),
.Y(n_1047)
);

INVx4_ASAP7_75t_L g1048 ( 
.A(n_1027),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_1031),
.B(n_884),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_989),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_974),
.Y(n_1051)
);

AND2x4_ASAP7_75t_L g1052 ( 
.A(n_1027),
.B(n_951),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_997),
.B(n_953),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_989),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_989),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_963),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_987),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_969),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_1019),
.B(n_889),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_991),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1035),
.B(n_1036),
.Y(n_1061)
);

INVx5_ASAP7_75t_L g1062 ( 
.A(n_1013),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_992),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_999),
.Y(n_1064)
);

INVx4_ASAP7_75t_SL g1065 ( 
.A(n_1024),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_980),
.B(n_896),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_970),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_1004),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_R g1069 ( 
.A(n_967),
.B(n_832),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1000),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1006),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1007),
.Y(n_1072)
);

AOI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_970),
.A2(n_951),
.B1(n_779),
.B2(n_761),
.Y(n_1073)
);

XOR2x2_ASAP7_75t_L g1074 ( 
.A(n_1002),
.B(n_832),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_976),
.Y(n_1075)
);

AND2x6_ASAP7_75t_L g1076 ( 
.A(n_1012),
.B(n_934),
.Y(n_1076)
);

INVx4_ASAP7_75t_L g1077 ( 
.A(n_1028),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_972),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1005),
.Y(n_1079)
);

NAND3xp33_ASAP7_75t_L g1080 ( 
.A(n_983),
.B(n_956),
.C(n_953),
.Y(n_1080)
);

INVx5_ASAP7_75t_L g1081 ( 
.A(n_975),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_1003),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1040),
.B(n_953),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_1032),
.B(n_889),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1023),
.B(n_953),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1008),
.B(n_919),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_975),
.B(n_895),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1005),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1028),
.B(n_919),
.Y(n_1089)
);

INVxp67_ASAP7_75t_L g1090 ( 
.A(n_966),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_968),
.A2(n_900),
.B1(n_924),
.B2(n_643),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_1009),
.Y(n_1092)
);

BUFx10_ASAP7_75t_L g1093 ( 
.A(n_972),
.Y(n_1093)
);

INVx4_ASAP7_75t_L g1094 ( 
.A(n_995),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_985),
.B(n_902),
.Y(n_1095)
);

NAND3x1_ASAP7_75t_L g1096 ( 
.A(n_964),
.B(n_838),
.C(n_835),
.Y(n_1096)
);

OR2x2_ASAP7_75t_L g1097 ( 
.A(n_1010),
.B(n_819),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_1029),
.B(n_900),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_1003),
.Y(n_1099)
);

OR2x2_ASAP7_75t_L g1100 ( 
.A(n_977),
.B(n_900),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1026),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1038),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_986),
.B(n_990),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1039),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1014),
.Y(n_1105)
);

INVx1_ASAP7_75t_SL g1106 ( 
.A(n_996),
.Y(n_1106)
);

NAND2x1p5_ASAP7_75t_L g1107 ( 
.A(n_1003),
.B(n_929),
.Y(n_1107)
);

INVx6_ASAP7_75t_L g1108 ( 
.A(n_979),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_965),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_979),
.B(n_993),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_979),
.B(n_924),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_994),
.B(n_924),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_998),
.B(n_908),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_973),
.Y(n_1114)
);

INVx6_ASAP7_75t_L g1115 ( 
.A(n_996),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1018),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1018),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1001),
.B(n_921),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1041),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1011),
.B(n_921),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1041),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_1018),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_978),
.B(n_948),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1041),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1014),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_968),
.A2(n_691),
.B1(n_762),
.B2(n_672),
.Y(n_1126)
);

AND2x4_ASAP7_75t_L g1127 ( 
.A(n_982),
.B(n_956),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1033),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1015),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_1016),
.B(n_910),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_1017),
.Y(n_1131)
);

INVx6_ASAP7_75t_L g1132 ( 
.A(n_1020),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1015),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_1021),
.B(n_913),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1033),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_981),
.B(n_956),
.Y(n_1136)
);

INVx4_ASAP7_75t_L g1137 ( 
.A(n_1033),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_981),
.A2(n_788),
.B1(n_948),
.B2(n_936),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_1022),
.Y(n_1139)
);

AND2x6_ASAP7_75t_L g1140 ( 
.A(n_1022),
.B(n_948),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_1030),
.B(n_928),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_988),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_988),
.Y(n_1143)
);

AND2x6_ASAP7_75t_L g1144 ( 
.A(n_1025),
.B(n_572),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_1004),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_989),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_984),
.B(n_937),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_1019),
.B(n_835),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_1004),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_971),
.Y(n_1150)
);

HB1xp67_ASAP7_75t_L g1151 ( 
.A(n_1004),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_967),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_1031),
.B(n_939),
.Y(n_1153)
);

INVx5_ASAP7_75t_L g1154 ( 
.A(n_1034),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_1034),
.A2(n_957),
.B1(n_958),
.B2(n_940),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_971),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_989),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_1019),
.B(n_838),
.Y(n_1158)
);

OR2x2_ASAP7_75t_L g1159 ( 
.A(n_966),
.B(n_962),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_963),
.Y(n_1160)
);

INVxp67_ASAP7_75t_SL g1161 ( 
.A(n_1023),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_989),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1019),
.B(n_850),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_969),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_1031),
.B(n_593),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1147),
.B(n_678),
.Y(n_1166)
);

NOR2xp67_ASAP7_75t_L g1167 ( 
.A(n_1056),
.B(n_814),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_1061),
.B(n_878),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1066),
.B(n_850),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1046),
.B(n_582),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1051),
.Y(n_1171)
);

NAND2x1_ASAP7_75t_L g1172 ( 
.A(n_1137),
.B(n_911),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_1148),
.B(n_878),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_1081),
.B(n_603),
.Y(n_1174)
);

NOR2xp67_ASAP7_75t_L g1175 ( 
.A(n_1160),
.B(n_817),
.Y(n_1175)
);

NAND2x1_ASAP7_75t_L g1176 ( 
.A(n_1137),
.B(n_1140),
.Y(n_1176)
);

NOR2xp67_ASAP7_75t_L g1177 ( 
.A(n_1109),
.B(n_858),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1053),
.A2(n_687),
.B(n_583),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1087),
.A2(n_1158),
.B(n_1163),
.C(n_1110),
.Y(n_1179)
);

INVx2_ASAP7_75t_SL g1180 ( 
.A(n_1062),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1089),
.B(n_550),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1057),
.Y(n_1182)
);

NAND2xp33_ASAP7_75t_L g1183 ( 
.A(n_1081),
.B(n_608),
.Y(n_1183)
);

NAND2x1p5_ASAP7_75t_L g1184 ( 
.A(n_1131),
.B(n_911),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1108),
.A2(n_803),
.B1(n_807),
.B2(n_799),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1113),
.B(n_644),
.Y(n_1186)
);

INVxp33_ASAP7_75t_SL g1187 ( 
.A(n_1069),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1060),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1063),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1067),
.Y(n_1190)
);

NOR2xp67_ASAP7_75t_L g1191 ( 
.A(n_1062),
.B(n_859),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_1048),
.B(n_614),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1045),
.B(n_1059),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1064),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1130),
.B(n_1134),
.Y(n_1195)
);

INVx2_ASAP7_75t_SL g1196 ( 
.A(n_1062),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1070),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1111),
.A2(n_712),
.B1(n_653),
.B2(n_883),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1052),
.B(n_883),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_1149),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_1068),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1164),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1048),
.B(n_615),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_1052),
.B(n_893),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1071),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1047),
.B(n_790),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1108),
.A2(n_1159),
.B1(n_1138),
.B2(n_1073),
.Y(n_1207)
);

INVx2_ASAP7_75t_SL g1208 ( 
.A(n_1132),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1047),
.B(n_797),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1042),
.A2(n_893),
.B1(n_852),
.B2(n_652),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1042),
.B(n_797),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1126),
.A2(n_852),
.B1(n_652),
.B2(n_671),
.Y(n_1212)
);

AND2x6_ASAP7_75t_L g1213 ( 
.A(n_1139),
.B(n_1078),
.Y(n_1213)
);

INVxp67_ASAP7_75t_SL g1214 ( 
.A(n_1145),
.Y(n_1214)
);

O2A1O1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1043),
.A2(n_611),
.B(n_809),
.C(n_860),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1136),
.B(n_863),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1072),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1150),
.B(n_588),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_SL g1219 ( 
.A(n_1077),
.B(n_1094),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1151),
.B(n_1090),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1075),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_1077),
.B(n_620),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1156),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1079),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_1094),
.B(n_622),
.Y(n_1225)
);

NAND2xp33_ASAP7_75t_SL g1226 ( 
.A(n_1044),
.B(n_623),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1049),
.B(n_629),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1088),
.Y(n_1228)
);

INVxp67_ASAP7_75t_L g1229 ( 
.A(n_1092),
.Y(n_1229)
);

INVx5_ASAP7_75t_L g1230 ( 
.A(n_1140),
.Y(n_1230)
);

AND3x1_ASAP7_75t_L g1231 ( 
.A(n_1123),
.B(n_868),
.C(n_864),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1086),
.B(n_612),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1162),
.B(n_617),
.Y(n_1233)
);

O2A1O1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1084),
.A2(n_870),
.B(n_871),
.C(n_869),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1085),
.A2(n_544),
.B(n_542),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1118),
.B(n_633),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1154),
.B(n_651),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_SL g1238 ( 
.A(n_1154),
.B(n_655),
.Y(n_1238)
);

INVx4_ASAP7_75t_L g1239 ( 
.A(n_1154),
.Y(n_1239)
);

NAND2xp33_ASAP7_75t_L g1240 ( 
.A(n_1140),
.B(n_658),
.Y(n_1240)
);

AOI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1153),
.A2(n_625),
.B1(n_642),
.B2(n_619),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1120),
.B(n_659),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1152),
.B(n_661),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1065),
.B(n_872),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1161),
.B(n_663),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1083),
.B(n_666),
.Y(n_1246)
);

NAND2xp33_ASAP7_75t_L g1247 ( 
.A(n_1140),
.B(n_668),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1101),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1155),
.B(n_1098),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1074),
.A2(n_671),
.B1(n_652),
.B2(n_562),
.Y(n_1250)
);

AOI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1095),
.A2(n_660),
.B1(n_664),
.B2(n_649),
.Y(n_1251)
);

OAI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1080),
.A2(n_676),
.B(n_665),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1098),
.B(n_669),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1102),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1112),
.B(n_673),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_1065),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1097),
.B(n_1091),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1165),
.B(n_674),
.Y(n_1258)
);

NOR2x1p5_ASAP7_75t_L g1259 ( 
.A(n_1114),
.B(n_873),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_1127),
.B(n_680),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1105),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1112),
.B(n_681),
.Y(n_1262)
);

INVxp67_ASAP7_75t_SL g1263 ( 
.A(n_1162),
.Y(n_1263)
);

NAND3xp33_ASAP7_75t_L g1264 ( 
.A(n_1116),
.B(n_756),
.C(n_710),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1100),
.B(n_690),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1104),
.A2(n_671),
.B1(n_737),
.B2(n_713),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_1127),
.B(n_692),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1076),
.B(n_693),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1076),
.B(n_1103),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1141),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1141),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1093),
.B(n_694),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1117),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1144),
.A2(n_1125),
.B1(n_1133),
.B2(n_1129),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1139),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1076),
.B(n_696),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1076),
.B(n_700),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1103),
.B(n_703),
.Y(n_1278)
);

AOI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1119),
.A2(n_697),
.B1(n_706),
.B2(n_677),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1121),
.A2(n_724),
.B1(n_728),
.B2(n_711),
.Y(n_1280)
);

NOR3xp33_ASAP7_75t_L g1281 ( 
.A(n_1106),
.B(n_738),
.C(n_730),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1124),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1128),
.B(n_740),
.Y(n_1283)
);

NAND2xp33_ASAP7_75t_L g1284 ( 
.A(n_1050),
.B(n_741),
.Y(n_1284)
);

O2A1O1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1135),
.A2(n_876),
.B(n_881),
.C(n_874),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1107),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1093),
.B(n_1082),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_1050),
.B(n_749),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1050),
.B(n_752),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1143),
.B(n_753),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1139),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1054),
.B(n_764),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1054),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1054),
.B(n_768),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1055),
.B(n_769),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1055),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1055),
.B(n_774),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1142),
.B(n_885),
.Y(n_1298)
);

NAND2xp33_ASAP7_75t_L g1299 ( 
.A(n_1082),
.B(n_776),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1082),
.B(n_1099),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1099),
.B(n_777),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1099),
.B(n_1122),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1122),
.B(n_780),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_SL g1304 ( 
.A(n_1122),
.B(n_782),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1146),
.B(n_784),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_SL g1306 ( 
.A(n_1115),
.B(n_543),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1146),
.B(n_787),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_SL g1308 ( 
.A(n_1146),
.B(n_789),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1157),
.B(n_707),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1157),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_1115),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1144),
.B(n_709),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_1144),
.B(n_792),
.Y(n_1313)
);

AOI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1144),
.A2(n_717),
.B1(n_722),
.B2(n_715),
.Y(n_1314)
);

NOR3xp33_ASAP7_75t_L g1315 ( 
.A(n_1096),
.B(n_804),
.C(n_794),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1066),
.B(n_891),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1138),
.A2(n_713),
.B1(n_899),
.B2(n_898),
.Y(n_1317)
);

AO221x1_ASAP7_75t_L g1318 ( 
.A1(n_1045),
.A2(n_638),
.B1(n_554),
.B2(n_731),
.C(n_725),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1147),
.B(n_742),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1147),
.B(n_750),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1058),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1147),
.B(n_755),
.Y(n_1322)
);

INVx8_ASAP7_75t_L g1323 ( 
.A(n_1062),
.Y(n_1323)
);

BUFx8_ASAP7_75t_L g1324 ( 
.A(n_1044),
.Y(n_1324)
);

INVx2_ASAP7_75t_SL g1325 ( 
.A(n_1062),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1046),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1061),
.B(n_713),
.Y(n_1327)
);

OAI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1061),
.A2(n_773),
.B1(n_785),
.B2(n_760),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1147),
.B(n_800),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1147),
.B(n_806),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_SL g1331 ( 
.A(n_1081),
.B(n_545),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1147),
.B(n_594),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1061),
.A2(n_598),
.B1(n_662),
.B2(n_572),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1147),
.B(n_718),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_1056),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1046),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1046),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1056),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1058),
.Y(n_1339)
);

NAND2x1p5_ASAP7_75t_L g1340 ( 
.A(n_1131),
.B(n_911),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1273),
.A2(n_662),
.B(n_598),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1195),
.B(n_911),
.Y(n_1342)
);

BUFx2_ASAP7_75t_L g1343 ( 
.A(n_1200),
.Y(n_1343)
);

OAI21xp33_ASAP7_75t_L g1344 ( 
.A1(n_1193),
.A2(n_748),
.B(n_575),
.Y(n_1344)
);

OAI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1282),
.A2(n_748),
.B(n_576),
.Y(n_1345)
);

BUFx4f_ASAP7_75t_L g1346 ( 
.A(n_1323),
.Y(n_1346)
);

NAND3xp33_ASAP7_75t_L g1347 ( 
.A(n_1173),
.B(n_914),
.C(n_578),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1216),
.B(n_914),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1300),
.A2(n_793),
.B(n_783),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1168),
.B(n_568),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_1230),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1179),
.B(n_914),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1186),
.B(n_914),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1316),
.B(n_0),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1171),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1332),
.B(n_2),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1323),
.Y(n_1357)
);

NAND3xp33_ASAP7_75t_SL g1358 ( 
.A(n_1327),
.B(n_624),
.C(n_601),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1323),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1319),
.A2(n_581),
.B(n_580),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1257),
.B(n_2),
.Y(n_1361)
);

BUFx4f_ASAP7_75t_L g1362 ( 
.A(n_1213),
.Y(n_1362)
);

AND2x4_ASAP7_75t_L g1363 ( 
.A(n_1239),
.B(n_3),
.Y(n_1363)
);

BUFx12f_ASAP7_75t_L g1364 ( 
.A(n_1324),
.Y(n_1364)
);

AOI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1233),
.A2(n_736),
.B(n_686),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1182),
.Y(n_1366)
);

INVxp67_ASAP7_75t_SL g1367 ( 
.A(n_1201),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1169),
.B(n_4),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1319),
.A2(n_587),
.B(n_584),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1334),
.B(n_4),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1188),
.Y(n_1371)
);

O2A1O1Ixp33_ASAP7_75t_L g1372 ( 
.A1(n_1328),
.A2(n_8),
.B(n_5),
.C(n_6),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1181),
.B(n_5),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1320),
.A2(n_600),
.B(n_596),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_SL g1375 ( 
.A(n_1220),
.B(n_602),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1166),
.B(n_8),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1322),
.B(n_9),
.Y(n_1377)
);

INVxp67_ASAP7_75t_L g1378 ( 
.A(n_1214),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1189),
.Y(n_1379)
);

BUFx6f_ASAP7_75t_L g1380 ( 
.A(n_1213),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1233),
.A2(n_605),
.B(n_604),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1322),
.A2(n_609),
.B(n_607),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1335),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1199),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1329),
.B(n_9),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1330),
.A2(n_621),
.B(n_616),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1330),
.B(n_10),
.Y(n_1387)
);

INVx8_ASAP7_75t_L g1388 ( 
.A(n_1213),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1248),
.Y(n_1389)
);

BUFx6f_ASAP7_75t_L g1390 ( 
.A(n_1213),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1254),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1298),
.B(n_11),
.Y(n_1392)
);

NOR3xp33_ASAP7_75t_L g1393 ( 
.A(n_1272),
.B(n_808),
.C(n_628),
.Y(n_1393)
);

AOI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1207),
.A2(n_627),
.B1(n_645),
.B2(n_630),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1194),
.Y(n_1395)
);

OAI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1197),
.A2(n_654),
.B(n_650),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1249),
.B(n_12),
.Y(n_1397)
);

AO21x1_ASAP7_75t_L g1398 ( 
.A1(n_1333),
.A2(n_1309),
.B(n_1252),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1204),
.B(n_656),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1207),
.A2(n_638),
.B1(n_554),
.B2(n_657),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_SL g1401 ( 
.A(n_1208),
.B(n_805),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1221),
.Y(n_1402)
);

BUFx12f_ASAP7_75t_L g1403 ( 
.A(n_1324),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1311),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1244),
.B(n_1265),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1263),
.A2(n_675),
.B(n_667),
.Y(n_1406)
);

CKINVDCx20_ASAP7_75t_R g1407 ( 
.A(n_1338),
.Y(n_1407)
);

AOI21xp33_ASAP7_75t_L g1408 ( 
.A1(n_1227),
.A2(n_688),
.B(n_682),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1211),
.B(n_13),
.Y(n_1409)
);

BUFx12f_ASAP7_75t_L g1410 ( 
.A(n_1259),
.Y(n_1410)
);

AND2x4_ASAP7_75t_L g1411 ( 
.A(n_1239),
.B(n_13),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1187),
.B(n_689),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1205),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1217),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1206),
.B(n_15),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1256),
.B(n_15),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1290),
.B(n_16),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1246),
.A2(n_699),
.B(n_695),
.Y(n_1418)
);

OAI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1223),
.A2(n_705),
.B(n_702),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1326),
.Y(n_1420)
);

INVx3_ASAP7_75t_L g1421 ( 
.A(n_1230),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1229),
.B(n_716),
.Y(n_1422)
);

O2A1O1Ixp33_ASAP7_75t_L g1423 ( 
.A1(n_1333),
.A2(n_18),
.B(n_16),
.C(n_17),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1336),
.Y(n_1424)
);

BUFx3_ASAP7_75t_L g1425 ( 
.A(n_1180),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1302),
.A2(n_727),
.B(n_720),
.Y(n_1426)
);

A2O1A1Ixp33_ASAP7_75t_L g1427 ( 
.A1(n_1258),
.A2(n_1252),
.B(n_1241),
.C(n_1178),
.Y(n_1427)
);

AOI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1231),
.A2(n_733),
.B1(n_747),
.B2(n_734),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1176),
.A2(n_1172),
.B(n_1240),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1209),
.B(n_17),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_SL g1431 ( 
.A(n_1177),
.B(n_751),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1236),
.B(n_1242),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1337),
.B(n_18),
.Y(n_1433)
);

AND2x4_ASAP7_75t_L g1434 ( 
.A(n_1269),
.B(n_1196),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1295),
.B(n_19),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1247),
.A2(n_758),
.B(n_757),
.Y(n_1436)
);

AOI21xp33_ASAP7_75t_L g1437 ( 
.A1(n_1237),
.A2(n_763),
.B(n_759),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_SL g1438 ( 
.A(n_1306),
.B(n_798),
.Y(n_1438)
);

AOI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1235),
.A2(n_1218),
.B(n_1170),
.Y(n_1439)
);

AND2x4_ASAP7_75t_L g1440 ( 
.A(n_1325),
.B(n_20),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1190),
.Y(n_1441)
);

INVx3_ASAP7_75t_L g1442 ( 
.A(n_1230),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1297),
.B(n_20),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1230),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1270),
.B(n_21),
.Y(n_1445)
);

INVx3_ASAP7_75t_L g1446 ( 
.A(n_1293),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1191),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_SL g1448 ( 
.A(n_1167),
.B(n_765),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1271),
.B(n_22),
.Y(n_1449)
);

O2A1O1Ixp33_ASAP7_75t_L g1450 ( 
.A1(n_1185),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1170),
.A2(n_771),
.B(n_766),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1198),
.B(n_778),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1313),
.B(n_23),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1218),
.A2(n_781),
.B(n_638),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1296),
.A2(n_638),
.B(n_554),
.Y(n_1455)
);

OAI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1224),
.A2(n_736),
.B(n_686),
.Y(n_1456)
);

OAI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1228),
.A2(n_736),
.B(n_686),
.Y(n_1457)
);

O2A1O1Ixp33_ASAP7_75t_L g1458 ( 
.A1(n_1185),
.A2(n_26),
.B(n_24),
.C(n_25),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1245),
.B(n_27),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1202),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1232),
.B(n_27),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1283),
.A2(n_554),
.B(n_292),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1275),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_L g1464 ( 
.A(n_1260),
.B(n_28),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1317),
.B(n_28),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1310),
.A2(n_296),
.B(n_290),
.Y(n_1466)
);

INVx3_ASAP7_75t_L g1467 ( 
.A(n_1291),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1232),
.B(n_29),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1274),
.B(n_30),
.Y(n_1469)
);

INVxp67_ASAP7_75t_L g1470 ( 
.A(n_1253),
.Y(n_1470)
);

OR2x6_ASAP7_75t_L g1471 ( 
.A(n_1267),
.B(n_30),
.Y(n_1471)
);

NOR2x1p5_ASAP7_75t_SL g1472 ( 
.A(n_1321),
.B(n_686),
.Y(n_1472)
);

INVx3_ASAP7_75t_L g1473 ( 
.A(n_1184),
.Y(n_1473)
);

INVx11_ASAP7_75t_L g1474 ( 
.A(n_1175),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1312),
.B(n_33),
.Y(n_1475)
);

OAI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1309),
.A2(n_736),
.B(n_686),
.Y(n_1476)
);

NAND3xp33_ASAP7_75t_L g1477 ( 
.A(n_1183),
.B(n_33),
.C(n_34),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1339),
.Y(n_1478)
);

AOI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1288),
.A2(n_736),
.B(n_686),
.Y(n_1479)
);

OAI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1278),
.A2(n_1219),
.B1(n_1262),
.B2(n_1255),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_1314),
.B(n_736),
.Y(n_1481)
);

A2O1A1Ixp33_ASAP7_75t_L g1482 ( 
.A1(n_1215),
.A2(n_736),
.B(n_36),
.C(n_34),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1261),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1287),
.B(n_35),
.Y(n_1484)
);

BUFx6f_ASAP7_75t_L g1485 ( 
.A(n_1184),
.Y(n_1485)
);

BUFx3_ASAP7_75t_L g1486 ( 
.A(n_1340),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1312),
.B(n_35),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1250),
.B(n_1212),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1280),
.B(n_37),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1268),
.B(n_37),
.Y(n_1490)
);

O2A1O1Ixp5_ASAP7_75t_L g1491 ( 
.A1(n_1292),
.A2(n_1308),
.B(n_1304),
.C(n_1331),
.Y(n_1491)
);

INVx2_ASAP7_75t_SL g1492 ( 
.A(n_1340),
.Y(n_1492)
);

OAI321xp33_ASAP7_75t_L g1493 ( 
.A1(n_1210),
.A2(n_40),
.A3(n_43),
.B1(n_38),
.B2(n_39),
.C(n_42),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1285),
.Y(n_1494)
);

AOI21x1_ASAP7_75t_L g1495 ( 
.A1(n_1289),
.A2(n_299),
.B(n_297),
.Y(n_1495)
);

AND2x4_ASAP7_75t_L g1496 ( 
.A(n_1286),
.B(n_38),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1280),
.B(n_40),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1294),
.A2(n_304),
.B(n_302),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1301),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1303),
.B(n_45),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1234),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_L g1502 ( 
.A(n_1276),
.B(n_46),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1305),
.Y(n_1503)
);

AO21x1_ASAP7_75t_L g1504 ( 
.A1(n_1277),
.A2(n_307),
.B(n_305),
.Y(n_1504)
);

NAND3xp33_ASAP7_75t_L g1505 ( 
.A(n_1251),
.B(n_46),
.C(n_47),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1307),
.A2(n_1203),
.B(n_1192),
.Y(n_1506)
);

AOI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1222),
.A2(n_309),
.B(n_308),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1266),
.B(n_47),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1279),
.B(n_48),
.Y(n_1509)
);

OAI21xp33_ASAP7_75t_L g1510 ( 
.A1(n_1225),
.A2(n_48),
.B(n_49),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1318),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1238),
.B(n_49),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1243),
.B(n_51),
.Y(n_1513)
);

A2O1A1Ixp33_ASAP7_75t_L g1514 ( 
.A1(n_1264),
.A2(n_1284),
.B(n_1299),
.C(n_1174),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1315),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1405),
.B(n_1281),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1343),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_SL g1518 ( 
.A(n_1362),
.B(n_1226),
.Y(n_1518)
);

A2O1A1Ixp33_ASAP7_75t_SL g1519 ( 
.A1(n_1513),
.A2(n_55),
.B(n_53),
.C(n_54),
.Y(n_1519)
);

AOI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1439),
.A2(n_312),
.B(n_311),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1342),
.A2(n_1432),
.B(n_1352),
.Y(n_1521)
);

A2O1A1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1427),
.A2(n_59),
.B(n_57),
.C(n_58),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1384),
.B(n_58),
.Y(n_1523)
);

O2A1O1Ixp5_ASAP7_75t_L g1524 ( 
.A1(n_1453),
.A2(n_61),
.B(n_59),
.C(n_60),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_SL g1525 ( 
.A(n_1362),
.B(n_313),
.Y(n_1525)
);

BUFx8_ASAP7_75t_SL g1526 ( 
.A(n_1364),
.Y(n_1526)
);

BUFx2_ASAP7_75t_L g1527 ( 
.A(n_1367),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1378),
.B(n_60),
.Y(n_1528)
);

AOI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1429),
.A2(n_319),
.B(n_315),
.Y(n_1529)
);

AOI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1381),
.A2(n_321),
.B(n_320),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1350),
.B(n_61),
.Y(n_1531)
);

OAI22x1_ASAP7_75t_L g1532 ( 
.A1(n_1394),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1361),
.B(n_62),
.Y(n_1533)
);

A2O1A1Ixp33_ASAP7_75t_L g1534 ( 
.A1(n_1344),
.A2(n_65),
.B(n_63),
.C(n_64),
.Y(n_1534)
);

CKINVDCx20_ASAP7_75t_R g1535 ( 
.A(n_1407),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1355),
.Y(n_1536)
);

AOI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1377),
.A2(n_324),
.B(n_322),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1399),
.B(n_65),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1385),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_1539)
);

AOI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1452),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1383),
.B(n_69),
.Y(n_1541)
);

AOI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1387),
.A2(n_328),
.B(n_327),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1456),
.A2(n_331),
.B(n_330),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1366),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_SL g1545 ( 
.A(n_1380),
.B(n_70),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1392),
.B(n_70),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1503),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_SL g1548 ( 
.A(n_1380),
.B(n_72),
.Y(n_1548)
);

OAI21xp33_ASAP7_75t_L g1549 ( 
.A1(n_1510),
.A2(n_73),
.B(n_75),
.Y(n_1549)
);

NAND3xp33_ASAP7_75t_L g1550 ( 
.A(n_1435),
.B(n_73),
.C(n_76),
.Y(n_1550)
);

NOR2xp67_ASAP7_75t_L g1551 ( 
.A(n_1470),
.B(n_334),
.Y(n_1551)
);

AOI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1457),
.A2(n_336),
.B(n_335),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1368),
.B(n_77),
.Y(n_1553)
);

NOR3xp33_ASAP7_75t_SL g1554 ( 
.A(n_1358),
.B(n_77),
.C(n_78),
.Y(n_1554)
);

AOI21xp5_ASAP7_75t_L g1555 ( 
.A1(n_1476),
.A2(n_339),
.B(n_338),
.Y(n_1555)
);

OA21x2_ASAP7_75t_L g1556 ( 
.A1(n_1365),
.A2(n_342),
.B(n_341),
.Y(n_1556)
);

INVx2_ASAP7_75t_SL g1557 ( 
.A(n_1346),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1462),
.A2(n_348),
.B(n_345),
.Y(n_1558)
);

BUFx10_ASAP7_75t_L g1559 ( 
.A(n_1412),
.Y(n_1559)
);

O2A1O1Ixp33_ASAP7_75t_L g1560 ( 
.A1(n_1443),
.A2(n_1497),
.B(n_1489),
.C(n_1417),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1371),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1379),
.B(n_79),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1395),
.Y(n_1563)
);

A2O1A1Ixp33_ASAP7_75t_SL g1564 ( 
.A1(n_1490),
.A2(n_82),
.B(n_80),
.C(n_81),
.Y(n_1564)
);

AO22x1_ASAP7_75t_L g1565 ( 
.A1(n_1488),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_1565)
);

AOI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1461),
.A2(n_351),
.B(n_349),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1496),
.B(n_84),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1438),
.B(n_85),
.Y(n_1568)
);

AOI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1468),
.A2(n_355),
.B(n_353),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1413),
.B(n_86),
.Y(n_1570)
);

O2A1O1Ixp33_ASAP7_75t_L g1571 ( 
.A1(n_1480),
.A2(n_1510),
.B(n_1373),
.C(n_1459),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1354),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.Y(n_1572)
);

AOI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1506),
.A2(n_358),
.B(n_356),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1414),
.B(n_87),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1420),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1424),
.Y(n_1576)
);

NOR2x1_ASAP7_75t_L g1577 ( 
.A(n_1404),
.B(n_359),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1389),
.B(n_89),
.Y(n_1578)
);

NOR2xp67_ASAP7_75t_L g1579 ( 
.A(n_1347),
.B(n_361),
.Y(n_1579)
);

A2O1A1Ixp33_ASAP7_75t_L g1580 ( 
.A1(n_1502),
.A2(n_91),
.B(n_89),
.C(n_90),
.Y(n_1580)
);

INVx3_ASAP7_75t_L g1581 ( 
.A(n_1388),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1391),
.B(n_90),
.Y(n_1582)
);

AOI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1348),
.A2(n_364),
.B(n_362),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1402),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1460),
.Y(n_1585)
);

NOR3xp33_ASAP7_75t_SL g1586 ( 
.A(n_1499),
.B(n_91),
.C(n_93),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_SL g1587 ( 
.A(n_1380),
.B(n_93),
.Y(n_1587)
);

OAI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1408),
.A2(n_94),
.B(n_95),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1446),
.Y(n_1589)
);

OAI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1494),
.A2(n_97),
.B1(n_94),
.B2(n_96),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1422),
.B(n_96),
.Y(n_1591)
);

BUFx6f_ASAP7_75t_L g1592 ( 
.A(n_1390),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1496),
.B(n_97),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1465),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1390),
.B(n_98),
.Y(n_1595)
);

INVx2_ASAP7_75t_SL g1596 ( 
.A(n_1346),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1376),
.B(n_99),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1396),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.Y(n_1598)
);

AOI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1454),
.A2(n_366),
.B(n_365),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1356),
.B(n_102),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_1403),
.Y(n_1601)
);

BUFx2_ASAP7_75t_L g1602 ( 
.A(n_1410),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1370),
.B(n_104),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_SL g1604 ( 
.A(n_1388),
.B(n_367),
.Y(n_1604)
);

INVx4_ASAP7_75t_L g1605 ( 
.A(n_1390),
.Y(n_1605)
);

NOR3xp33_ASAP7_75t_L g1606 ( 
.A(n_1493),
.B(n_105),
.C(n_106),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1397),
.B(n_106),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1393),
.B(n_107),
.Y(n_1608)
);

BUFx3_ASAP7_75t_L g1609 ( 
.A(n_1359),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1446),
.Y(n_1610)
);

O2A1O1Ixp33_ASAP7_75t_L g1611 ( 
.A1(n_1464),
.A2(n_109),
.B(n_107),
.C(n_108),
.Y(n_1611)
);

BUFx6f_ASAP7_75t_L g1612 ( 
.A(n_1357),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1434),
.B(n_108),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1341),
.A2(n_370),
.B(n_369),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1441),
.Y(n_1615)
);

BUFx3_ASAP7_75t_L g1616 ( 
.A(n_1357),
.Y(n_1616)
);

A2O1A1Ixp33_ASAP7_75t_L g1617 ( 
.A1(n_1345),
.A2(n_111),
.B(n_109),
.C(n_110),
.Y(n_1617)
);

AOI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1353),
.A2(n_374),
.B(n_372),
.Y(n_1618)
);

CKINVDCx10_ASAP7_75t_R g1619 ( 
.A(n_1471),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1434),
.B(n_110),
.Y(n_1620)
);

BUFx6f_ASAP7_75t_L g1621 ( 
.A(n_1357),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_SL g1622 ( 
.A(n_1416),
.B(n_375),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1498),
.A2(n_377),
.B(n_376),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_SL g1624 ( 
.A(n_1363),
.B(n_111),
.Y(n_1624)
);

OAI21x1_ASAP7_75t_L g1625 ( 
.A1(n_1479),
.A2(n_381),
.B(n_380),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_SL g1626 ( 
.A(n_1416),
.B(n_1486),
.Y(n_1626)
);

BUFx2_ASAP7_75t_L g1627 ( 
.A(n_1425),
.Y(n_1627)
);

INVx3_ASAP7_75t_L g1628 ( 
.A(n_1351),
.Y(n_1628)
);

O2A1O1Ixp33_ASAP7_75t_L g1629 ( 
.A1(n_1482),
.A2(n_114),
.B(n_112),
.C(n_113),
.Y(n_1629)
);

AOI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1514),
.A2(n_384),
.B(n_382),
.Y(n_1630)
);

INVx3_ASAP7_75t_L g1631 ( 
.A(n_1351),
.Y(n_1631)
);

O2A1O1Ixp33_ASAP7_75t_L g1632 ( 
.A1(n_1372),
.A2(n_117),
.B(n_115),
.C(n_116),
.Y(n_1632)
);

A2O1A1Ixp33_ASAP7_75t_L g1633 ( 
.A1(n_1500),
.A2(n_120),
.B(n_117),
.C(n_118),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1478),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1421),
.Y(n_1635)
);

BUFx6f_ASAP7_75t_L g1636 ( 
.A(n_1485),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1483),
.B(n_118),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1363),
.B(n_121),
.Y(n_1638)
);

AOI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1398),
.A2(n_386),
.B(n_385),
.Y(n_1639)
);

A2O1A1Ixp33_ASAP7_75t_L g1640 ( 
.A1(n_1475),
.A2(n_123),
.B(n_121),
.C(n_122),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1473),
.B(n_538),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1433),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1445),
.Y(n_1643)
);

OAI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1419),
.A2(n_126),
.B1(n_123),
.B2(n_124),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1449),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1409),
.Y(n_1646)
);

NAND2xp33_ASAP7_75t_L g1647 ( 
.A(n_1485),
.B(n_126),
.Y(n_1647)
);

BUFx6f_ASAP7_75t_L g1648 ( 
.A(n_1485),
.Y(n_1648)
);

AOI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1501),
.A2(n_389),
.B(n_388),
.Y(n_1649)
);

AOI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1466),
.A2(n_394),
.B(n_392),
.Y(n_1650)
);

OAI21xp33_ASAP7_75t_SL g1651 ( 
.A1(n_1509),
.A2(n_127),
.B(n_128),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_SL g1652 ( 
.A(n_1411),
.B(n_128),
.Y(n_1652)
);

A2O1A1Ixp33_ASAP7_75t_SL g1653 ( 
.A1(n_1507),
.A2(n_131),
.B(n_129),
.C(n_130),
.Y(n_1653)
);

NOR3xp33_ASAP7_75t_L g1654 ( 
.A(n_1450),
.B(n_129),
.C(n_130),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_SL g1655 ( 
.A(n_1411),
.B(n_131),
.Y(n_1655)
);

OAI22xp5_ASAP7_75t_L g1656 ( 
.A1(n_1428),
.A2(n_135),
.B1(n_132),
.B2(n_134),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1415),
.B(n_134),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1375),
.B(n_135),
.Y(n_1658)
);

BUFx3_ASAP7_75t_L g1659 ( 
.A(n_1463),
.Y(n_1659)
);

AO22x1_ASAP7_75t_L g1660 ( 
.A1(n_1512),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.Y(n_1660)
);

INVx3_ASAP7_75t_L g1661 ( 
.A(n_1421),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1536),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1544),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1567),
.B(n_1440),
.Y(n_1664)
);

AO31x2_ASAP7_75t_L g1665 ( 
.A1(n_1521),
.A2(n_1504),
.A3(n_1511),
.B(n_1455),
.Y(n_1665)
);

AO21x2_ASAP7_75t_L g1666 ( 
.A1(n_1639),
.A2(n_1487),
.B(n_1437),
.Y(n_1666)
);

INVx4_ASAP7_75t_L g1667 ( 
.A(n_1612),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1593),
.B(n_1440),
.Y(n_1668)
);

BUFx2_ASAP7_75t_SL g1669 ( 
.A(n_1535),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1527),
.B(n_1484),
.Y(n_1670)
);

AOI21x1_ASAP7_75t_L g1671 ( 
.A1(n_1520),
.A2(n_1495),
.B(n_1481),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1561),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1659),
.B(n_1473),
.Y(n_1673)
);

O2A1O1Ixp5_ASAP7_75t_L g1674 ( 
.A1(n_1522),
.A2(n_1491),
.B(n_1469),
.C(n_1430),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1563),
.Y(n_1675)
);

A2O1A1Ixp33_ASAP7_75t_L g1676 ( 
.A1(n_1560),
.A2(n_1458),
.B(n_1428),
.C(n_1423),
.Y(n_1676)
);

NOR3xp33_ASAP7_75t_L g1677 ( 
.A(n_1531),
.B(n_1477),
.C(n_1505),
.Y(n_1677)
);

AOI211x1_ASAP7_75t_L g1678 ( 
.A1(n_1660),
.A2(n_1508),
.B(n_1401),
.C(n_1431),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1517),
.B(n_1484),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1547),
.B(n_1512),
.Y(n_1680)
);

AOI21xp5_ASAP7_75t_SL g1681 ( 
.A1(n_1571),
.A2(n_1492),
.B(n_1471),
.Y(n_1681)
);

AOI21x1_ASAP7_75t_L g1682 ( 
.A1(n_1543),
.A2(n_1369),
.B(n_1360),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1643),
.B(n_1467),
.Y(n_1683)
);

INVxp67_ASAP7_75t_SL g1684 ( 
.A(n_1589),
.Y(n_1684)
);

AND2x2_ASAP7_75t_SL g1685 ( 
.A(n_1622),
.B(n_1400),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1575),
.Y(n_1686)
);

HB1xp67_ASAP7_75t_L g1687 ( 
.A(n_1610),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1645),
.B(n_1642),
.Y(n_1688)
);

NOR2xp67_ASAP7_75t_L g1689 ( 
.A(n_1557),
.B(n_1447),
.Y(n_1689)
);

A2O1A1Ixp33_ASAP7_75t_L g1690 ( 
.A1(n_1538),
.A2(n_1374),
.B(n_1386),
.C(n_1382),
.Y(n_1690)
);

A2O1A1Ixp33_ASAP7_75t_L g1691 ( 
.A1(n_1549),
.A2(n_1451),
.B(n_1515),
.C(n_1418),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1559),
.B(n_1463),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1576),
.Y(n_1693)
);

INVx8_ASAP7_75t_L g1694 ( 
.A(n_1526),
.Y(n_1694)
);

AOI21x1_ASAP7_75t_L g1695 ( 
.A1(n_1552),
.A2(n_1436),
.B(n_1349),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_R g1696 ( 
.A1(n_1601),
.A2(n_1474),
.B1(n_1448),
.B2(n_139),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1585),
.Y(n_1697)
);

A2O1A1Ixp33_ASAP7_75t_L g1698 ( 
.A1(n_1658),
.A2(n_1406),
.B(n_1426),
.C(n_1472),
.Y(n_1698)
);

OA21x2_ASAP7_75t_L g1699 ( 
.A1(n_1555),
.A2(n_1467),
.B(n_1463),
.Y(n_1699)
);

OAI21x1_ASAP7_75t_L g1700 ( 
.A1(n_1625),
.A2(n_1444),
.B(n_1442),
.Y(n_1700)
);

AOI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1530),
.A2(n_1444),
.B(n_1442),
.Y(n_1701)
);

INVx6_ASAP7_75t_SL g1702 ( 
.A(n_1559),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1630),
.A2(n_136),
.B(n_138),
.Y(n_1703)
);

OAI21x1_ASAP7_75t_SL g1704 ( 
.A1(n_1588),
.A2(n_139),
.B(n_140),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1626),
.B(n_141),
.Y(n_1705)
);

AOI21x1_ASAP7_75t_L g1706 ( 
.A1(n_1529),
.A2(n_396),
.B(n_395),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_SL g1707 ( 
.A1(n_1534),
.A2(n_141),
.B(n_142),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1646),
.B(n_143),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1516),
.B(n_144),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_SL g1710 ( 
.A(n_1592),
.B(n_145),
.Y(n_1710)
);

AOI21x1_ASAP7_75t_L g1711 ( 
.A1(n_1579),
.A2(n_402),
.B(n_399),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1546),
.B(n_146),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_SL g1713 ( 
.A(n_1604),
.B(n_405),
.Y(n_1713)
);

OAI21x1_ASAP7_75t_L g1714 ( 
.A1(n_1573),
.A2(n_408),
.B(n_406),
.Y(n_1714)
);

AND3x4_ASAP7_75t_L g1715 ( 
.A(n_1609),
.B(n_146),
.C(n_147),
.Y(n_1715)
);

OAI21x1_ASAP7_75t_L g1716 ( 
.A1(n_1558),
.A2(n_410),
.B(n_409),
.Y(n_1716)
);

OAI21x1_ASAP7_75t_L g1717 ( 
.A1(n_1623),
.A2(n_1599),
.B(n_1650),
.Y(n_1717)
);

A2O1A1Ixp33_ASAP7_75t_L g1718 ( 
.A1(n_1591),
.A2(n_150),
.B(n_148),
.C(n_149),
.Y(n_1718)
);

OAI21x1_ASAP7_75t_L g1719 ( 
.A1(n_1556),
.A2(n_416),
.B(n_414),
.Y(n_1719)
);

OAI21x1_ASAP7_75t_L g1720 ( 
.A1(n_1556),
.A2(n_418),
.B(n_417),
.Y(n_1720)
);

BUFx2_ASAP7_75t_L g1721 ( 
.A(n_1627),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1523),
.B(n_148),
.Y(n_1722)
);

INVx2_ASAP7_75t_SL g1723 ( 
.A(n_1616),
.Y(n_1723)
);

AO32x2_ASAP7_75t_L g1724 ( 
.A1(n_1539),
.A2(n_151),
.A3(n_152),
.B1(n_154),
.B2(n_156),
.Y(n_1724)
);

OAI21x1_ASAP7_75t_L g1725 ( 
.A1(n_1618),
.A2(n_421),
.B(n_419),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1533),
.B(n_152),
.Y(n_1726)
);

NOR2x1_ASAP7_75t_SL g1727 ( 
.A(n_1518),
.B(n_156),
.Y(n_1727)
);

INVx1_ASAP7_75t_SL g1728 ( 
.A(n_1619),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1553),
.B(n_157),
.Y(n_1729)
);

BUFx6f_ASAP7_75t_L g1730 ( 
.A(n_1592),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_SL g1731 ( 
.A(n_1525),
.B(n_422),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1615),
.Y(n_1732)
);

OAI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1617),
.A2(n_158),
.B(n_159),
.Y(n_1733)
);

OAI21x1_ASAP7_75t_L g1734 ( 
.A1(n_1614),
.A2(n_428),
.B(n_426),
.Y(n_1734)
);

AOI21x1_ASAP7_75t_L g1735 ( 
.A1(n_1607),
.A2(n_433),
.B(n_430),
.Y(n_1735)
);

OAI21x1_ASAP7_75t_L g1736 ( 
.A1(n_1583),
.A2(n_436),
.B(n_434),
.Y(n_1736)
);

NAND2x1p5_ASAP7_75t_L g1737 ( 
.A(n_1605),
.B(n_437),
.Y(n_1737)
);

BUFx6f_ASAP7_75t_L g1738 ( 
.A(n_1592),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1528),
.B(n_158),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1634),
.Y(n_1740)
);

AOI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1649),
.A2(n_160),
.B(n_161),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1562),
.B(n_161),
.Y(n_1742)
);

BUFx6f_ASAP7_75t_L g1743 ( 
.A(n_1612),
.Y(n_1743)
);

AOI221xp5_ASAP7_75t_L g1744 ( 
.A1(n_1611),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.C(n_165),
.Y(n_1744)
);

OAI21x1_ASAP7_75t_L g1745 ( 
.A1(n_1537),
.A2(n_439),
.B(n_438),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1613),
.B(n_162),
.Y(n_1746)
);

AOI221xp5_ASAP7_75t_L g1747 ( 
.A1(n_1532),
.A2(n_163),
.B1(n_165),
.B2(n_166),
.C(n_167),
.Y(n_1747)
);

OAI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1540),
.A2(n_169),
.B1(n_167),
.B2(n_168),
.Y(n_1748)
);

AO32x2_ASAP7_75t_L g1749 ( 
.A1(n_1590),
.A2(n_168),
.A3(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1620),
.B(n_171),
.Y(n_1750)
);

OAI21xp5_ASAP7_75t_L g1751 ( 
.A1(n_1598),
.A2(n_172),
.B(n_173),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1597),
.B(n_173),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1581),
.B(n_174),
.Y(n_1753)
);

OAI21x1_ASAP7_75t_L g1754 ( 
.A1(n_1542),
.A2(n_1569),
.B(n_1566),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1570),
.B(n_1574),
.Y(n_1755)
);

AOI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1647),
.A2(n_174),
.B(n_175),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1584),
.B(n_1624),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1608),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.Y(n_1758)
);

OAI21x1_ASAP7_75t_L g1759 ( 
.A1(n_1628),
.A2(n_442),
.B(n_440),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1638),
.B(n_176),
.Y(n_1760)
);

NOR2xp67_ASAP7_75t_L g1761 ( 
.A(n_1596),
.B(n_443),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_SL g1762 ( 
.A(n_1636),
.B(n_178),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1652),
.B(n_179),
.Y(n_1763)
);

NOR4xp25_ASAP7_75t_L g1764 ( 
.A(n_1580),
.B(n_181),
.C(n_179),
.D(n_180),
.Y(n_1764)
);

AOI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1653),
.A2(n_182),
.B(n_183),
.Y(n_1765)
);

AO21x1_ASAP7_75t_L g1766 ( 
.A1(n_1644),
.A2(n_184),
.B(n_185),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1655),
.B(n_184),
.Y(n_1767)
);

OAI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1751),
.A2(n_1550),
.B(n_1586),
.Y(n_1768)
);

AND2x2_ASAP7_75t_SL g1769 ( 
.A(n_1685),
.B(n_1606),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1697),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1733),
.A2(n_1654),
.B1(n_1656),
.B2(n_1594),
.Y(n_1771)
);

OAI221xp5_ASAP7_75t_SL g1772 ( 
.A1(n_1747),
.A2(n_1640),
.B1(n_1633),
.B2(n_1651),
.C(n_1632),
.Y(n_1772)
);

AO21x1_ASAP7_75t_L g1773 ( 
.A1(n_1758),
.A2(n_1568),
.B(n_1572),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1755),
.B(n_1541),
.Y(n_1774)
);

BUFx4f_ASAP7_75t_L g1775 ( 
.A(n_1694),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1662),
.Y(n_1776)
);

OAI21x1_ASAP7_75t_L g1777 ( 
.A1(n_1717),
.A2(n_1671),
.B(n_1754),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_SL g1778 ( 
.A(n_1713),
.B(n_1577),
.Y(n_1778)
);

OAI21x1_ASAP7_75t_L g1779 ( 
.A1(n_1719),
.A2(n_1524),
.B(n_1628),
.Y(n_1779)
);

OAI21x1_ASAP7_75t_L g1780 ( 
.A1(n_1720),
.A2(n_1635),
.B(n_1631),
.Y(n_1780)
);

NAND3xp33_ASAP7_75t_L g1781 ( 
.A(n_1677),
.B(n_1565),
.C(n_1554),
.Y(n_1781)
);

OAI21x1_ASAP7_75t_L g1782 ( 
.A1(n_1701),
.A2(n_1635),
.B(n_1631),
.Y(n_1782)
);

AOI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1715),
.A2(n_1600),
.B1(n_1603),
.B2(n_1657),
.Y(n_1783)
);

AOI22xp33_ASAP7_75t_L g1784 ( 
.A1(n_1766),
.A2(n_1551),
.B1(n_1582),
.B2(n_1578),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1664),
.B(n_1661),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1663),
.Y(n_1786)
);

AOI21x1_ASAP7_75t_L g1787 ( 
.A1(n_1735),
.A2(n_1548),
.B(n_1545),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1668),
.B(n_1687),
.Y(n_1788)
);

NAND3xp33_ASAP7_75t_L g1789 ( 
.A(n_1744),
.B(n_1519),
.C(n_1629),
.Y(n_1789)
);

O2A1O1Ixp5_ASAP7_75t_L g1790 ( 
.A1(n_1748),
.A2(n_1587),
.B(n_1595),
.C(n_1564),
.Y(n_1790)
);

O2A1O1Ixp33_ASAP7_75t_SL g1791 ( 
.A1(n_1676),
.A2(n_1637),
.B(n_1661),
.C(n_1581),
.Y(n_1791)
);

INVx3_ASAP7_75t_L g1792 ( 
.A(n_1730),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1684),
.B(n_1636),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1712),
.B(n_1612),
.Y(n_1794)
);

OAI21x1_ASAP7_75t_L g1795 ( 
.A1(n_1700),
.A2(n_1648),
.B(n_1636),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1729),
.B(n_1621),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_L g1797 ( 
.A(n_1709),
.B(n_1621),
.Y(n_1797)
);

BUFx6f_ASAP7_75t_L g1798 ( 
.A(n_1730),
.Y(n_1798)
);

OAI21x1_ASAP7_75t_L g1799 ( 
.A1(n_1706),
.A2(n_1648),
.B(n_1641),
.Y(n_1799)
);

BUFx2_ASAP7_75t_L g1800 ( 
.A(n_1702),
.Y(n_1800)
);

INVx4_ASAP7_75t_L g1801 ( 
.A(n_1743),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1672),
.Y(n_1802)
);

OAI21x1_ASAP7_75t_L g1803 ( 
.A1(n_1695),
.A2(n_1641),
.B(n_1621),
.Y(n_1803)
);

OAI21x1_ASAP7_75t_L g1804 ( 
.A1(n_1734),
.A2(n_446),
.B(n_445),
.Y(n_1804)
);

AOI221xp5_ASAP7_75t_SL g1805 ( 
.A1(n_1718),
.A2(n_1602),
.B1(n_187),
.B2(n_188),
.C(n_190),
.Y(n_1805)
);

AOI332xp33_ASAP7_75t_L g1806 ( 
.A1(n_1752),
.A2(n_186),
.A3(n_187),
.B1(n_188),
.B2(n_190),
.B3(n_191),
.C1(n_192),
.C2(n_193),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_L g1807 ( 
.A(n_1670),
.B(n_186),
.Y(n_1807)
);

OAI21x1_ASAP7_75t_L g1808 ( 
.A1(n_1682),
.A2(n_449),
.B(n_447),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1705),
.B(n_192),
.Y(n_1809)
);

AO21x2_ASAP7_75t_L g1810 ( 
.A1(n_1666),
.A2(n_451),
.B(n_450),
.Y(n_1810)
);

OAI21x1_ASAP7_75t_L g1811 ( 
.A1(n_1714),
.A2(n_454),
.B(n_453),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1688),
.B(n_194),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1675),
.Y(n_1813)
);

OAI21x1_ASAP7_75t_L g1814 ( 
.A1(n_1716),
.A2(n_460),
.B(n_459),
.Y(n_1814)
);

OA21x2_ASAP7_75t_L g1815 ( 
.A1(n_1674),
.A2(n_464),
.B(n_463),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1686),
.Y(n_1816)
);

OR2x6_ASAP7_75t_L g1817 ( 
.A(n_1681),
.B(n_465),
.Y(n_1817)
);

OAI21x1_ASAP7_75t_L g1818 ( 
.A1(n_1711),
.A2(n_471),
.B(n_469),
.Y(n_1818)
);

OAI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1756),
.A2(n_195),
.B(n_196),
.Y(n_1819)
);

BUFx3_ASAP7_75t_L g1820 ( 
.A(n_1721),
.Y(n_1820)
);

OAI21xp5_ASAP7_75t_L g1821 ( 
.A1(n_1707),
.A2(n_195),
.B(n_196),
.Y(n_1821)
);

O2A1O1Ixp33_ASAP7_75t_L g1822 ( 
.A1(n_1691),
.A2(n_197),
.B(n_198),
.C(n_199),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1696),
.A2(n_197),
.B1(n_199),
.B2(n_200),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1693),
.B(n_201),
.Y(n_1824)
);

OAI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1741),
.A2(n_201),
.B(n_202),
.Y(n_1825)
);

NAND2x1p5_ASAP7_75t_L g1826 ( 
.A(n_1692),
.B(n_474),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1732),
.Y(n_1827)
);

OAI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1742),
.A2(n_1722),
.B1(n_1739),
.B2(n_1760),
.Y(n_1828)
);

BUFx3_ASAP7_75t_L g1829 ( 
.A(n_1743),
.Y(n_1829)
);

BUFx3_ASAP7_75t_L g1830 ( 
.A(n_1743),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1680),
.B(n_203),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1740),
.Y(n_1832)
);

AOI21xp5_ASAP7_75t_L g1833 ( 
.A1(n_1731),
.A2(n_205),
.B(n_206),
.Y(n_1833)
);

INVx3_ASAP7_75t_L g1834 ( 
.A(n_1730),
.Y(n_1834)
);

BUFx12f_ASAP7_75t_L g1835 ( 
.A(n_1723),
.Y(n_1835)
);

AOI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1791),
.A2(n_1703),
.B(n_1690),
.Y(n_1836)
);

OAI21x1_ASAP7_75t_L g1837 ( 
.A1(n_1777),
.A2(n_1699),
.B(n_1759),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1770),
.B(n_1679),
.Y(n_1838)
);

OAI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1769),
.A2(n_1764),
.B(n_1765),
.Y(n_1839)
);

OAI21x1_ASAP7_75t_L g1840 ( 
.A1(n_1777),
.A2(n_1808),
.B(n_1782),
.Y(n_1840)
);

AOI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1791),
.A2(n_1699),
.B(n_1698),
.Y(n_1841)
);

AOI21x1_ASAP7_75t_L g1842 ( 
.A1(n_1778),
.A2(n_1683),
.B(n_1689),
.Y(n_1842)
);

HB1xp67_ASAP7_75t_L g1843 ( 
.A(n_1820),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1774),
.B(n_1708),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1827),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1820),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1774),
.B(n_1726),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1769),
.B(n_1746),
.Y(n_1848)
);

INVx2_ASAP7_75t_SL g1849 ( 
.A(n_1793),
.Y(n_1849)
);

CKINVDCx8_ASAP7_75t_R g1850 ( 
.A(n_1800),
.Y(n_1850)
);

CKINVDCx20_ASAP7_75t_R g1851 ( 
.A(n_1775),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1802),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1816),
.B(n_1724),
.Y(n_1853)
);

OA21x2_ASAP7_75t_L g1854 ( 
.A1(n_1808),
.A2(n_1745),
.B(n_1704),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1832),
.Y(n_1855)
);

AOI21x1_ASAP7_75t_L g1856 ( 
.A1(n_1778),
.A2(n_1757),
.B(n_1762),
.Y(n_1856)
);

HB1xp67_ASAP7_75t_L g1857 ( 
.A(n_1776),
.Y(n_1857)
);

INVx1_ASAP7_75t_SL g1858 ( 
.A(n_1835),
.Y(n_1858)
);

OAI21x1_ASAP7_75t_L g1859 ( 
.A1(n_1782),
.A2(n_1779),
.B(n_1803),
.Y(n_1859)
);

NOR2xp33_ASAP7_75t_L g1860 ( 
.A(n_1828),
.B(n_1750),
.Y(n_1860)
);

INVx2_ASAP7_75t_SL g1861 ( 
.A(n_1786),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1813),
.B(n_1669),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1788),
.B(n_1665),
.Y(n_1863)
);

OAI21x1_ASAP7_75t_L g1864 ( 
.A1(n_1779),
.A2(n_1725),
.B(n_1736),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1824),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1812),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1795),
.Y(n_1867)
);

OAI21xp5_ASAP7_75t_L g1868 ( 
.A1(n_1781),
.A2(n_1710),
.B(n_1763),
.Y(n_1868)
);

AOI21xp5_ASAP7_75t_L g1869 ( 
.A1(n_1822),
.A2(n_1737),
.B(n_1727),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1857),
.Y(n_1870)
);

INVx2_ASAP7_75t_SL g1871 ( 
.A(n_1843),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1863),
.B(n_1831),
.Y(n_1872)
);

INVx2_ASAP7_75t_SL g1873 ( 
.A(n_1846),
.Y(n_1873)
);

BUFx12f_ASAP7_75t_L g1874 ( 
.A(n_1862),
.Y(n_1874)
);

HB1xp67_ASAP7_75t_L g1875 ( 
.A(n_1861),
.Y(n_1875)
);

INVx4_ASAP7_75t_L g1876 ( 
.A(n_1854),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1863),
.B(n_1785),
.Y(n_1877)
);

INVx1_ASAP7_75t_SL g1878 ( 
.A(n_1838),
.Y(n_1878)
);

OR2x6_ASAP7_75t_L g1879 ( 
.A(n_1841),
.B(n_1817),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1861),
.B(n_1849),
.Y(n_1880)
);

BUFx6f_ASAP7_75t_L g1881 ( 
.A(n_1859),
.Y(n_1881)
);

AO21x2_ASAP7_75t_L g1882 ( 
.A1(n_1836),
.A2(n_1810),
.B(n_1821),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1845),
.Y(n_1883)
);

INVx3_ASAP7_75t_L g1884 ( 
.A(n_1859),
.Y(n_1884)
);

HB1xp67_ASAP7_75t_L g1885 ( 
.A(n_1867),
.Y(n_1885)
);

OA21x2_ASAP7_75t_L g1886 ( 
.A1(n_1840),
.A2(n_1837),
.B(n_1864),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1852),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1855),
.Y(n_1888)
);

OA21x2_ASAP7_75t_L g1889 ( 
.A1(n_1840),
.A2(n_1780),
.B(n_1784),
.Y(n_1889)
);

OAI321xp33_ASAP7_75t_L g1890 ( 
.A1(n_1879),
.A2(n_1823),
.A3(n_1839),
.B1(n_1860),
.B2(n_1848),
.C(n_1768),
.Y(n_1890)
);

AOI22xp33_ASAP7_75t_L g1891 ( 
.A1(n_1882),
.A2(n_1773),
.B1(n_1848),
.B2(n_1860),
.Y(n_1891)
);

OAI22xp33_ASAP7_75t_L g1892 ( 
.A1(n_1879),
.A2(n_1817),
.B1(n_1844),
.B2(n_1847),
.Y(n_1892)
);

OAI33xp33_ASAP7_75t_L g1893 ( 
.A1(n_1872),
.A2(n_1866),
.A3(n_1865),
.B1(n_1806),
.B2(n_1767),
.B3(n_1789),
.Y(n_1893)
);

AND2x4_ASAP7_75t_L g1894 ( 
.A(n_1877),
.B(n_1849),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1877),
.B(n_1850),
.Y(n_1895)
);

AOI22xp33_ASAP7_75t_L g1896 ( 
.A1(n_1882),
.A2(n_1823),
.B1(n_1784),
.B2(n_1817),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1883),
.Y(n_1897)
);

INVxp67_ASAP7_75t_L g1898 ( 
.A(n_1875),
.Y(n_1898)
);

BUFx4f_ASAP7_75t_SL g1899 ( 
.A(n_1874),
.Y(n_1899)
);

AOI21xp5_ASAP7_75t_L g1900 ( 
.A1(n_1879),
.A2(n_1869),
.B(n_1833),
.Y(n_1900)
);

AOI22xp33_ASAP7_75t_L g1901 ( 
.A1(n_1882),
.A2(n_1879),
.B1(n_1872),
.B2(n_1771),
.Y(n_1901)
);

AOI22xp33_ASAP7_75t_L g1902 ( 
.A1(n_1882),
.A2(n_1771),
.B1(n_1819),
.B2(n_1825),
.Y(n_1902)
);

AOI22xp33_ASAP7_75t_SL g1903 ( 
.A1(n_1879),
.A2(n_1853),
.B1(n_1809),
.B2(n_1810),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1879),
.A2(n_1783),
.B1(n_1853),
.B2(n_1809),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1870),
.Y(n_1905)
);

INVx1_ASAP7_75t_SL g1906 ( 
.A(n_1880),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1891),
.B(n_1870),
.Y(n_1907)
);

AND2x4_ASAP7_75t_L g1908 ( 
.A(n_1895),
.B(n_1871),
.Y(n_1908)
);

BUFx3_ASAP7_75t_L g1909 ( 
.A(n_1899),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1905),
.Y(n_1910)
);

INVx1_ASAP7_75t_SL g1911 ( 
.A(n_1899),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1897),
.Y(n_1912)
);

INVxp67_ASAP7_75t_SL g1913 ( 
.A(n_1891),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1894),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1908),
.B(n_1906),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1908),
.B(n_1898),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1910),
.B(n_1902),
.Y(n_1917)
);

NOR2x1_ASAP7_75t_SL g1918 ( 
.A(n_1914),
.B(n_1874),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1914),
.Y(n_1919)
);

OA21x2_ASAP7_75t_L g1920 ( 
.A1(n_1917),
.A2(n_1913),
.B(n_1907),
.Y(n_1920)
);

AOI221xp5_ASAP7_75t_L g1921 ( 
.A1(n_1917),
.A2(n_1890),
.B1(n_1893),
.B2(n_1904),
.C(n_1896),
.Y(n_1921)
);

OAI211xp5_ASAP7_75t_L g1922 ( 
.A1(n_1916),
.A2(n_1850),
.B(n_1900),
.C(n_1903),
.Y(n_1922)
);

NOR2x1_ASAP7_75t_L g1923 ( 
.A(n_1915),
.B(n_1909),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1918),
.B(n_1908),
.Y(n_1924)
);

INVx2_ASAP7_75t_SL g1925 ( 
.A(n_1919),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1921),
.B(n_1910),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1923),
.B(n_1911),
.Y(n_1927)
);

INVx4_ASAP7_75t_L g1928 ( 
.A(n_1924),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1927),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1928),
.Y(n_1930)
);

NOR2xp67_ASAP7_75t_L g1931 ( 
.A(n_1929),
.B(n_1928),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1931),
.B(n_1930),
.Y(n_1932)
);

AOI221xp5_ASAP7_75t_L g1933 ( 
.A1(n_1932),
.A2(n_1926),
.B1(n_1920),
.B2(n_1922),
.C(n_1925),
.Y(n_1933)
);

OAI21xp5_ASAP7_75t_L g1934 ( 
.A1(n_1932),
.A2(n_1920),
.B(n_1775),
.Y(n_1934)
);

AOI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1933),
.A2(n_1911),
.B1(n_1694),
.B2(n_1728),
.Y(n_1935)
);

AOI22xp5_ASAP7_75t_L g1936 ( 
.A1(n_1934),
.A2(n_1858),
.B1(n_1909),
.B2(n_1851),
.Y(n_1936)
);

OAI221xp5_ASAP7_75t_L g1937 ( 
.A1(n_1935),
.A2(n_1805),
.B1(n_1783),
.B2(n_1868),
.C(n_1901),
.Y(n_1937)
);

HB1xp67_ASAP7_75t_L g1938 ( 
.A(n_1936),
.Y(n_1938)
);

A2O1A1Ixp33_ASAP7_75t_L g1939 ( 
.A1(n_1935),
.A2(n_1851),
.B(n_1807),
.C(n_1790),
.Y(n_1939)
);

AOI322xp5_ASAP7_75t_L g1940 ( 
.A1(n_1938),
.A2(n_1807),
.A3(n_1892),
.B1(n_1753),
.B2(n_1797),
.C1(n_1794),
.C2(n_1796),
.Y(n_1940)
);

NOR2x1_ASAP7_75t_L g1941 ( 
.A(n_1939),
.B(n_1753),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_SL g1942 ( 
.A(n_1937),
.B(n_1881),
.Y(n_1942)
);

NAND4xp75_ASAP7_75t_L g1943 ( 
.A(n_1941),
.B(n_1761),
.C(n_1702),
.D(n_1678),
.Y(n_1943)
);

AOI21xp5_ASAP7_75t_L g1944 ( 
.A1(n_1942),
.A2(n_1876),
.B(n_1892),
.Y(n_1944)
);

NAND4xp25_ASAP7_75t_SL g1945 ( 
.A(n_1940),
.B(n_1880),
.C(n_1835),
.D(n_1724),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1941),
.Y(n_1946)
);

AOI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1942),
.A2(n_1874),
.B1(n_1797),
.B2(n_1876),
.Y(n_1947)
);

OAI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1941),
.A2(n_1876),
.B1(n_1884),
.B2(n_1881),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1942),
.A2(n_1876),
.B(n_1884),
.Y(n_1949)
);

NOR2xp67_ASAP7_75t_L g1950 ( 
.A(n_1946),
.B(n_205),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1947),
.B(n_1871),
.Y(n_1951)
);

NOR2xp67_ASAP7_75t_L g1952 ( 
.A(n_1945),
.B(n_206),
.Y(n_1952)
);

A2O1A1Ixp33_ASAP7_75t_L g1953 ( 
.A1(n_1944),
.A2(n_1884),
.B(n_1772),
.C(n_1912),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1943),
.Y(n_1954)
);

NOR2x1_ASAP7_75t_L g1955 ( 
.A(n_1949),
.B(n_207),
.Y(n_1955)
);

NOR2xp33_ASAP7_75t_L g1956 ( 
.A(n_1948),
.B(n_1912),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1946),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1946),
.Y(n_1958)
);

INVxp33_ASAP7_75t_SL g1959 ( 
.A(n_1946),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1950),
.Y(n_1960)
);

OR2x2_ASAP7_75t_L g1961 ( 
.A(n_1957),
.B(n_1871),
.Y(n_1961)
);

NAND4xp75_ASAP7_75t_L g1962 ( 
.A(n_1958),
.B(n_209),
.C(n_207),
.D(n_208),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1959),
.Y(n_1963)
);

NAND4xp75_ASAP7_75t_L g1964 ( 
.A(n_1955),
.B(n_210),
.C(n_208),
.D(n_209),
.Y(n_1964)
);

OAI22xp5_ASAP7_75t_L g1965 ( 
.A1(n_1953),
.A2(n_1884),
.B1(n_1873),
.B2(n_1881),
.Y(n_1965)
);

AND2x2_ASAP7_75t_SL g1966 ( 
.A(n_1954),
.B(n_1667),
.Y(n_1966)
);

NOR2x1_ASAP7_75t_L g1967 ( 
.A(n_1952),
.B(n_1951),
.Y(n_1967)
);

INVxp67_ASAP7_75t_SL g1968 ( 
.A(n_1956),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_L g1969 ( 
.A(n_1959),
.B(n_210),
.Y(n_1969)
);

AOI22xp5_ASAP7_75t_L g1970 ( 
.A1(n_1952),
.A2(n_1881),
.B1(n_1873),
.B2(n_1815),
.Y(n_1970)
);

AOI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1952),
.A2(n_1881),
.B1(n_1873),
.B2(n_1815),
.Y(n_1971)
);

NOR2x1_ASAP7_75t_L g1972 ( 
.A(n_1957),
.B(n_211),
.Y(n_1972)
);

AND2x4_ASAP7_75t_L g1973 ( 
.A(n_1957),
.B(n_1894),
.Y(n_1973)
);

NOR2xp67_ASAP7_75t_L g1974 ( 
.A(n_1957),
.B(n_211),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1957),
.Y(n_1975)
);

AOI22xp5_ASAP7_75t_L g1976 ( 
.A1(n_1952),
.A2(n_1881),
.B1(n_1815),
.B2(n_1854),
.Y(n_1976)
);

INVx1_ASAP7_75t_SL g1977 ( 
.A(n_1959),
.Y(n_1977)
);

NOR2x1_ASAP7_75t_L g1978 ( 
.A(n_1957),
.B(n_212),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1950),
.Y(n_1979)
);

OR2x2_ASAP7_75t_L g1980 ( 
.A(n_1957),
.B(n_213),
.Y(n_1980)
);

AOI22xp5_ASAP7_75t_L g1981 ( 
.A1(n_1952),
.A2(n_1881),
.B1(n_1854),
.B2(n_1826),
.Y(n_1981)
);

NOR2x1_ASAP7_75t_L g1982 ( 
.A(n_1957),
.B(n_213),
.Y(n_1982)
);

AOI22xp33_ASAP7_75t_L g1983 ( 
.A1(n_1952),
.A2(n_1889),
.B1(n_1826),
.B2(n_1885),
.Y(n_1983)
);

NOR2x1_ASAP7_75t_L g1984 ( 
.A(n_1957),
.B(n_214),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1957),
.Y(n_1985)
);

AOI22xp5_ASAP7_75t_L g1986 ( 
.A1(n_1975),
.A2(n_1886),
.B1(n_1889),
.B2(n_1804),
.Y(n_1986)
);

NOR3xp33_ASAP7_75t_L g1987 ( 
.A(n_1977),
.B(n_1963),
.C(n_1985),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1974),
.B(n_214),
.Y(n_1988)
);

AOI222xp33_ASAP7_75t_L g1989 ( 
.A1(n_1960),
.A2(n_1979),
.B1(n_1968),
.B2(n_1966),
.C1(n_1982),
.C2(n_1972),
.Y(n_1989)
);

AOI211xp5_ASAP7_75t_SL g1990 ( 
.A1(n_1969),
.A2(n_1961),
.B(n_1980),
.C(n_1973),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1978),
.B(n_215),
.Y(n_1991)
);

OA22x2_ASAP7_75t_L g1992 ( 
.A1(n_1973),
.A2(n_1667),
.B1(n_1801),
.B2(n_1811),
.Y(n_1992)
);

AOI22xp5_ASAP7_75t_L g1993 ( 
.A1(n_1967),
.A2(n_1886),
.B1(n_1889),
.B2(n_1811),
.Y(n_1993)
);

NAND4xp25_ASAP7_75t_L g1994 ( 
.A(n_1984),
.B(n_215),
.C(n_216),
.D(n_218),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1964),
.Y(n_1995)
);

OAI221xp5_ASAP7_75t_L g1996 ( 
.A1(n_1970),
.A2(n_1724),
.B1(n_1886),
.B2(n_220),
.C(n_221),
.Y(n_1996)
);

OA22x2_ASAP7_75t_L g1997 ( 
.A1(n_1981),
.A2(n_1801),
.B1(n_1814),
.B2(n_1792),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1962),
.B(n_218),
.Y(n_1998)
);

OAI222xp33_ASAP7_75t_L g1999 ( 
.A1(n_1971),
.A2(n_1856),
.B1(n_1842),
.B2(n_1749),
.C1(n_1787),
.C2(n_1878),
.Y(n_1999)
);

AOI221x1_ASAP7_75t_L g2000 ( 
.A1(n_1965),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.C(n_222),
.Y(n_2000)
);

AND3x1_ASAP7_75t_L g2001 ( 
.A(n_1983),
.B(n_219),
.C(n_223),
.Y(n_2001)
);

OAI221xp5_ASAP7_75t_SL g2002 ( 
.A1(n_1976),
.A2(n_1749),
.B1(n_226),
.B2(n_227),
.C(n_228),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1974),
.B(n_225),
.Y(n_2003)
);

OAI21xp33_ASAP7_75t_SL g2004 ( 
.A1(n_1977),
.A2(n_1864),
.B(n_225),
.Y(n_2004)
);

OAI211xp5_ASAP7_75t_SL g2005 ( 
.A1(n_1977),
.A2(n_229),
.B(n_230),
.C(n_231),
.Y(n_2005)
);

AOI21xp33_ASAP7_75t_SL g2006 ( 
.A1(n_1963),
.A2(n_230),
.B(n_231),
.Y(n_2006)
);

AOI211xp5_ASAP7_75t_L g2007 ( 
.A1(n_1977),
.A2(n_232),
.B(n_233),
.C(n_234),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_R g2008 ( 
.A(n_1963),
.B(n_232),
.Y(n_2008)
);

OAI221xp5_ASAP7_75t_SL g2009 ( 
.A1(n_1977),
.A2(n_1749),
.B1(n_235),
.B2(n_237),
.C(n_238),
.Y(n_2009)
);

AOI211xp5_ASAP7_75t_L g2010 ( 
.A1(n_1977),
.A2(n_234),
.B(n_235),
.C(n_237),
.Y(n_2010)
);

AO22x2_ASAP7_75t_L g2011 ( 
.A1(n_1977),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1974),
.B(n_239),
.Y(n_2012)
);

XNOR2xp5_ASAP7_75t_L g2013 ( 
.A(n_1977),
.B(n_240),
.Y(n_2013)
);

AND2x4_ASAP7_75t_L g2014 ( 
.A(n_1973),
.B(n_241),
.Y(n_2014)
);

NAND4xp75_ASAP7_75t_L g2015 ( 
.A(n_1972),
.B(n_242),
.C(n_243),
.D(n_244),
.Y(n_2015)
);

OAI22xp33_ASAP7_75t_L g2016 ( 
.A1(n_1975),
.A2(n_1886),
.B1(n_1889),
.B2(n_1798),
.Y(n_2016)
);

OAI221xp5_ASAP7_75t_L g2017 ( 
.A1(n_1977),
.A2(n_1886),
.B1(n_244),
.B2(n_245),
.C(n_246),
.Y(n_2017)
);

NAND4xp25_ASAP7_75t_L g2018 ( 
.A(n_1977),
.B(n_242),
.C(n_245),
.D(n_247),
.Y(n_2018)
);

OAI22xp5_ASAP7_75t_SL g2019 ( 
.A1(n_1977),
.A2(n_247),
.B1(n_248),
.B2(n_249),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_2011),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_2011),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_2015),
.Y(n_2022)
);

NOR2x1_ASAP7_75t_L g2023 ( 
.A(n_2018),
.B(n_252),
.Y(n_2023)
);

XOR2x2_ASAP7_75t_L g2024 ( 
.A(n_1987),
.B(n_253),
.Y(n_2024)
);

BUFx3_ASAP7_75t_L g2025 ( 
.A(n_2014),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_2014),
.B(n_253),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_2013),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_1990),
.B(n_1889),
.Y(n_2028)
);

AOI22xp5_ASAP7_75t_L g2029 ( 
.A1(n_2004),
.A2(n_1814),
.B1(n_1818),
.B2(n_1792),
.Y(n_2029)
);

XOR2x1_ASAP7_75t_SL g2030 ( 
.A(n_1995),
.B(n_254),
.Y(n_2030)
);

XNOR2x1_ASAP7_75t_L g2031 ( 
.A(n_1988),
.B(n_255),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1991),
.Y(n_2032)
);

AND3x4_ASAP7_75t_L g2033 ( 
.A(n_2005),
.B(n_256),
.C(n_257),
.Y(n_2033)
);

XNOR2xp5_ASAP7_75t_L g2034 ( 
.A(n_1994),
.B(n_256),
.Y(n_2034)
);

NOR2x1_ASAP7_75t_L g2035 ( 
.A(n_1998),
.B(n_258),
.Y(n_2035)
);

XNOR2xp5_ASAP7_75t_L g2036 ( 
.A(n_2003),
.B(n_258),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1989),
.B(n_259),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_2012),
.Y(n_2038)
);

AOI22xp33_ASAP7_75t_L g2039 ( 
.A1(n_1997),
.A2(n_1885),
.B1(n_1887),
.B2(n_1888),
.Y(n_2039)
);

HB1xp67_ASAP7_75t_L g2040 ( 
.A(n_2008),
.Y(n_2040)
);

OR2x2_ASAP7_75t_L g2041 ( 
.A(n_2006),
.B(n_260),
.Y(n_2041)
);

HB1xp67_ASAP7_75t_L g2042 ( 
.A(n_2019),
.Y(n_2042)
);

XNOR2x1_ASAP7_75t_L g2043 ( 
.A(n_2001),
.B(n_260),
.Y(n_2043)
);

NOR3xp33_ASAP7_75t_L g2044 ( 
.A(n_2007),
.B(n_261),
.C(n_262),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1992),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_2017),
.Y(n_2046)
);

OR2x2_ASAP7_75t_L g2047 ( 
.A(n_2002),
.B(n_262),
.Y(n_2047)
);

XNOR2x1_ASAP7_75t_L g2048 ( 
.A(n_2010),
.B(n_263),
.Y(n_2048)
);

OR2x6_ASAP7_75t_L g2049 ( 
.A(n_2000),
.B(n_1738),
.Y(n_2049)
);

XNOR2x1_ASAP7_75t_L g2050 ( 
.A(n_1993),
.B(n_1986),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1996),
.Y(n_2051)
);

XOR2xp5_ASAP7_75t_L g2052 ( 
.A(n_2009),
.B(n_264),
.Y(n_2052)
);

AO21x2_ASAP7_75t_L g2053 ( 
.A1(n_1999),
.A2(n_264),
.B(n_265),
.Y(n_2053)
);

NAND3x1_ASAP7_75t_L g2054 ( 
.A(n_2016),
.B(n_265),
.C(n_266),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_2011),
.Y(n_2055)
);

NAND2x1p5_ASAP7_75t_L g2056 ( 
.A(n_2014),
.B(n_1798),
.Y(n_2056)
);

NAND2xp33_ASAP7_75t_L g2057 ( 
.A(n_2042),
.B(n_266),
.Y(n_2057)
);

INVx1_ASAP7_75t_SL g2058 ( 
.A(n_2025),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_2030),
.Y(n_2059)
);

AND3x2_ASAP7_75t_L g2060 ( 
.A(n_2020),
.B(n_267),
.C(n_268),
.Y(n_2060)
);

OA22x2_ASAP7_75t_L g2061 ( 
.A1(n_2033),
.A2(n_267),
.B1(n_268),
.B2(n_269),
.Y(n_2061)
);

NAND2x1p5_ASAP7_75t_L g2062 ( 
.A(n_2035),
.B(n_1798),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_2043),
.Y(n_2063)
);

BUFx2_ASAP7_75t_L g2064 ( 
.A(n_2021),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_2049),
.Y(n_2065)
);

INVxp67_ASAP7_75t_L g2066 ( 
.A(n_2040),
.Y(n_2066)
);

INVx4_ASAP7_75t_L g2067 ( 
.A(n_2038),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_2049),
.Y(n_2068)
);

INVx3_ASAP7_75t_L g2069 ( 
.A(n_2056),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2034),
.Y(n_2070)
);

BUFx3_ASAP7_75t_L g2071 ( 
.A(n_2055),
.Y(n_2071)
);

XOR2x1_ASAP7_75t_L g2072 ( 
.A(n_2024),
.B(n_269),
.Y(n_2072)
);

OAI21xp5_ASAP7_75t_L g2073 ( 
.A1(n_2023),
.A2(n_1799),
.B(n_270),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_2028),
.B(n_270),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_2041),
.Y(n_2075)
);

INVx4_ASAP7_75t_L g2076 ( 
.A(n_2022),
.Y(n_2076)
);

XNOR2xp5_ASAP7_75t_L g2077 ( 
.A(n_2031),
.B(n_2036),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_2048),
.Y(n_2078)
);

AND2x2_ASAP7_75t_SL g2079 ( 
.A(n_2037),
.B(n_271),
.Y(n_2079)
);

AND2x4_ASAP7_75t_L g2080 ( 
.A(n_2027),
.B(n_271),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_2034),
.B(n_2036),
.Y(n_2081)
);

OAI22xp5_ASAP7_75t_L g2082 ( 
.A1(n_2066),
.A2(n_2045),
.B1(n_2052),
.B2(n_2029),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2061),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_2062),
.Y(n_2084)
);

NOR2xp33_ASAP7_75t_L g2085 ( 
.A(n_2076),
.B(n_2026),
.Y(n_2085)
);

OAI21x1_ASAP7_75t_L g2086 ( 
.A1(n_2072),
.A2(n_2054),
.B(n_2046),
.Y(n_2086)
);

AOI22xp5_ASAP7_75t_L g2087 ( 
.A1(n_2071),
.A2(n_2044),
.B1(n_2051),
.B2(n_2050),
.Y(n_2087)
);

AOI22xp5_ASAP7_75t_L g2088 ( 
.A1(n_2063),
.A2(n_2053),
.B1(n_2032),
.B2(n_2047),
.Y(n_2088)
);

BUFx2_ASAP7_75t_L g2089 ( 
.A(n_2064),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2077),
.Y(n_2090)
);

OAI22xp5_ASAP7_75t_L g2091 ( 
.A1(n_2058),
.A2(n_2039),
.B1(n_1834),
.B2(n_1830),
.Y(n_2091)
);

OAI22xp5_ASAP7_75t_L g2092 ( 
.A1(n_2065),
.A2(n_1834),
.B1(n_1829),
.B2(n_1830),
.Y(n_2092)
);

AOI31xp33_ASAP7_75t_L g2093 ( 
.A1(n_2059),
.A2(n_273),
.A3(n_274),
.B(n_275),
.Y(n_2093)
);

AOI22x1_ASAP7_75t_L g2094 ( 
.A1(n_2064),
.A2(n_273),
.B1(n_274),
.B2(n_276),
.Y(n_2094)
);

HB1xp67_ASAP7_75t_L g2095 ( 
.A(n_2077),
.Y(n_2095)
);

AOI31xp33_ASAP7_75t_L g2096 ( 
.A1(n_2068),
.A2(n_277),
.A3(n_278),
.B(n_279),
.Y(n_2096)
);

NOR2x1_ASAP7_75t_L g2097 ( 
.A(n_2067),
.B(n_277),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2060),
.Y(n_2098)
);

OAI22x1_ASAP7_75t_L g2099 ( 
.A1(n_2089),
.A2(n_2080),
.B1(n_2075),
.B2(n_2069),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2095),
.B(n_2081),
.Y(n_2100)
);

OAI21xp5_ASAP7_75t_L g2101 ( 
.A1(n_2085),
.A2(n_2070),
.B(n_2079),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2097),
.Y(n_2102)
);

XNOR2x1_ASAP7_75t_L g2103 ( 
.A(n_2090),
.B(n_2070),
.Y(n_2103)
);

XNOR2x1_ASAP7_75t_L g2104 ( 
.A(n_2087),
.B(n_2078),
.Y(n_2104)
);

OAI22xp5_ASAP7_75t_L g2105 ( 
.A1(n_2083),
.A2(n_2074),
.B1(n_2073),
.B2(n_2057),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_2098),
.B(n_279),
.Y(n_2106)
);

AO22x2_ASAP7_75t_L g2107 ( 
.A1(n_2084),
.A2(n_2082),
.B1(n_2086),
.B2(n_2088),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2096),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2093),
.Y(n_2109)
);

XNOR2xp5_ASAP7_75t_L g2110 ( 
.A(n_2103),
.B(n_2094),
.Y(n_2110)
);

AOI22xp5_ASAP7_75t_L g2111 ( 
.A1(n_2100),
.A2(n_2091),
.B1(n_2092),
.B2(n_283),
.Y(n_2111)
);

OAI21xp33_ASAP7_75t_L g2112 ( 
.A1(n_2099),
.A2(n_281),
.B(n_282),
.Y(n_2112)
);

OAI22xp5_ASAP7_75t_L g2113 ( 
.A1(n_2107),
.A2(n_281),
.B1(n_282),
.B2(n_284),
.Y(n_2113)
);

OAI22xp5_ASAP7_75t_L g2114 ( 
.A1(n_2107),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_2114)
);

OAI22xp5_ASAP7_75t_L g2115 ( 
.A1(n_2104),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2102),
.B(n_287),
.Y(n_2116)
);

CKINVDCx20_ASAP7_75t_R g2117 ( 
.A(n_2101),
.Y(n_2117)
);

OAI22xp5_ASAP7_75t_L g2118 ( 
.A1(n_2117),
.A2(n_2109),
.B1(n_2108),
.B2(n_2106),
.Y(n_2118)
);

NOR2xp33_ASAP7_75t_L g2119 ( 
.A(n_2110),
.B(n_2105),
.Y(n_2119)
);

AOI21xp33_ASAP7_75t_L g2120 ( 
.A1(n_2113),
.A2(n_288),
.B(n_289),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2116),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_SL g2122 ( 
.A(n_2114),
.B(n_288),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_2112),
.B(n_483),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2115),
.Y(n_2124)
);

AOI21xp5_ASAP7_75t_L g2125 ( 
.A1(n_2118),
.A2(n_2111),
.B(n_485),
.Y(n_2125)
);

AOI22xp33_ASAP7_75t_L g2126 ( 
.A1(n_2119),
.A2(n_1798),
.B1(n_1829),
.B2(n_1738),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_2121),
.Y(n_2127)
);

AOI22xp33_ASAP7_75t_L g2128 ( 
.A1(n_2122),
.A2(n_1738),
.B1(n_1867),
.B2(n_1888),
.Y(n_2128)
);

OA21x2_ASAP7_75t_L g2129 ( 
.A1(n_2124),
.A2(n_484),
.B(n_488),
.Y(n_2129)
);

OAI22x1_ASAP7_75t_L g2130 ( 
.A1(n_2127),
.A2(n_2123),
.B1(n_2120),
.B2(n_492),
.Y(n_2130)
);

OAI22xp5_ASAP7_75t_SL g2131 ( 
.A1(n_2129),
.A2(n_489),
.B1(n_491),
.B2(n_493),
.Y(n_2131)
);

AOI22xp33_ASAP7_75t_L g2132 ( 
.A1(n_2131),
.A2(n_2125),
.B1(n_2126),
.B2(n_2128),
.Y(n_2132)
);

AOI22xp5_ASAP7_75t_L g2133 ( 
.A1(n_2130),
.A2(n_1673),
.B1(n_495),
.B2(n_496),
.Y(n_2133)
);

OR2x6_ASAP7_75t_L g2134 ( 
.A(n_2132),
.B(n_1673),
.Y(n_2134)
);

AOI221xp5_ASAP7_75t_L g2135 ( 
.A1(n_2134),
.A2(n_2133),
.B1(n_497),
.B2(n_498),
.C(n_499),
.Y(n_2135)
);

AOI211xp5_ASAP7_75t_L g2136 ( 
.A1(n_2135),
.A2(n_494),
.B(n_501),
.C(n_502),
.Y(n_2136)
);


endmodule