module fake_jpeg_19506_n_257 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_39),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_17),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_26),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_1),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_24),
.Y(n_64)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_56),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_48),
.B(n_44),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_35),
.B1(n_23),
.B2(n_33),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_50),
.A2(n_63),
.B1(n_65),
.B2(n_39),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_30),
.B1(n_34),
.B2(n_25),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_52),
.A2(n_45),
.B1(n_38),
.B2(n_42),
.Y(n_76)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_19),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_17),
.B1(n_34),
.B2(n_25),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_57),
.A2(n_58),
.B1(n_45),
.B2(n_41),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_36),
.A2(n_29),
.B1(n_22),
.B2(n_33),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_29),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_24),
.Y(n_81)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_45),
.A2(n_35),
.B1(n_31),
.B2(n_23),
.Y(n_63)
);

FAx1_ASAP7_75t_SL g72 ( 
.A(n_64),
.B(n_32),
.CI(n_63),
.CON(n_72),
.SN(n_72)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_31),
.B1(n_28),
.B2(n_21),
.Y(n_65)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_68),
.B(n_81),
.Y(n_126)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g70 ( 
.A(n_56),
.B(n_44),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_72),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_41),
.B(n_42),
.C(n_38),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_79),
.Y(n_104)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_78),
.Y(n_106)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g115 ( 
.A(n_75),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_76),
.A2(n_88),
.B1(n_102),
.B2(n_43),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_51),
.Y(n_77)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_42),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_80),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_50),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_90),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_41),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_93),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_85),
.B(n_86),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_16),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_49),
.A2(n_39),
.B(n_24),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_20),
.C(n_2),
.Y(n_120)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_94),
.Y(n_118)
);

BUFx12_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_37),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_46),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_98),
.Y(n_122)
);

NAND2x1_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_39),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_39),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_16),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_43),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_93),
.Y(n_131)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_103),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_46),
.A2(n_39),
.B1(n_27),
.B2(n_21),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_53),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_105),
.A2(n_119),
.B(n_96),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_43),
.B1(n_21),
.B2(n_20),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_108),
.B1(n_113),
.B2(n_124),
.Y(n_140)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_109),
.B(n_130),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_74),
.A2(n_20),
.B1(n_19),
.B2(n_27),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_71),
.B(n_27),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_4),
.Y(n_149)
);

AND2x6_ASAP7_75t_L g121 ( 
.A(n_70),
.B(n_15),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_121),
.B(n_128),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_74),
.B(n_1),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_123),
.B(n_3),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_79),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_124)
);

AND2x6_ASAP7_75t_L g128 ( 
.A(n_72),
.B(n_15),
.Y(n_128)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_87),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_131),
.A2(n_84),
.B1(n_99),
.B2(n_72),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_133),
.A2(n_154),
.B1(n_157),
.B2(n_5),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_134),
.A2(n_147),
.B(n_153),
.Y(n_159)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_144),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_111),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_137),
.B(n_139),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_89),
.C(n_101),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_152),
.C(n_10),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_118),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_149),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_100),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_106),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_145),
.B(n_156),
.Y(n_178)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_146),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_119),
.A2(n_92),
.B(n_67),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_148),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_116),
.A2(n_90),
.B1(n_77),
.B2(n_75),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_150),
.A2(n_115),
.B1(n_130),
.B2(n_109),
.Y(n_167)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_158),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_92),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_119),
.A2(n_89),
.B(n_6),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_104),
.A2(n_97),
.B1(n_101),
.B2(n_7),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_5),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_114),
.A2(n_97),
.B1(n_6),
.B2(n_8),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_5),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_151),
.A2(n_135),
.B1(n_115),
.B2(n_148),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_160),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_140),
.A2(n_128),
.B1(n_107),
.B2(n_121),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_167),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_126),
.B1(n_120),
.B2(n_122),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_164),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_136),
.A2(n_113),
.B1(n_105),
.B2(n_124),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_168),
.A2(n_138),
.B1(n_158),
.B2(n_153),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_134),
.A2(n_144),
.B(n_147),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_169),
.A2(n_172),
.B(n_175),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_137),
.A2(n_105),
.B1(n_127),
.B2(n_8),
.Y(n_171)
);

INVx13_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_142),
.A2(n_123),
.B(n_127),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_155),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_174),
.B(n_181),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_150),
.A2(n_6),
.B(n_9),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_12),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_156),
.B(n_14),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_173),
.Y(n_187)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_189),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_159),
.B(n_166),
.Y(n_189)
);

AND2x4_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_154),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_174),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_166),
.A2(n_133),
.B1(n_146),
.B2(n_157),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_196),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_152),
.C(n_143),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_179),
.C(n_165),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_149),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_161),
.Y(n_201)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_165),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_176),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_179),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_178),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_203),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_172),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_168),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_207),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_209),
.A2(n_199),
.B(n_190),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_211),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_196),
.Y(n_212)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_212),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_175),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_215),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_216),
.A2(n_225),
.B1(n_162),
.B2(n_180),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_206),
.A2(n_186),
.B1(n_190),
.B2(n_185),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_220),
.A2(n_224),
.B1(n_207),
.B2(n_204),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_190),
.B(n_193),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_203),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_191),
.B1(n_200),
.B2(n_186),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_183),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_226),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_205),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_228),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_213),
.A2(n_162),
.B(n_180),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_228),
.Y(n_231)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_231),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_235),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_220),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_182),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_234),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_225),
.B(n_198),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_236),
.B(n_237),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_217),
.B(n_201),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_233),
.A2(n_224),
.B1(n_216),
.B2(n_223),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_242),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_241),
.A2(n_230),
.B1(n_208),
.B2(n_184),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_247),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_238),
.A2(n_242),
.B(n_229),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_240),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_187),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_219),
.C(n_235),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_249),
.Y(n_252)
);

AOI322xp5_ASAP7_75t_L g251 ( 
.A1(n_250),
.A2(n_184),
.A3(n_222),
.B1(n_243),
.B2(n_232),
.C1(n_217),
.C2(n_237),
.Y(n_251)
);

XNOR2x2_ASAP7_75t_SL g254 ( 
.A(n_251),
.B(n_248),
.Y(n_254)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_252),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_253),
.B(n_254),
.C(n_194),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_167),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_14),
.Y(n_257)
);


endmodule