module real_jpeg_33457_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_11;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_9;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_0),
.Y(n_128)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_0),
.Y(n_140)
);

OAI32xp33_ASAP7_75t_L g39 ( 
.A1(n_1),
.A2(n_40),
.A3(n_42),
.B1(n_47),
.B2(n_53),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_1),
.Y(n_48)
);

OAI22x1_ASAP7_75t_SL g65 ( 
.A1(n_1),
.A2(n_48),
.B1(n_66),
.B2(n_71),
.Y(n_65)
);

AO22x1_ASAP7_75t_SL g119 ( 
.A1(n_1),
.A2(n_19),
.B1(n_48),
.B2(n_91),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_1),
.B(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_2),
.Y(n_148)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_2),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_4),
.A2(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_16)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_4),
.A2(n_20),
.B1(n_101),
.B2(n_104),
.Y(n_100)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_5),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_5),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_6),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_6),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_6),
.A2(n_35),
.B1(n_158),
.B2(n_160),
.Y(n_157)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_7),
.Y(n_82)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_7),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_131),
.Y(n_8)
);

HB1xp67_ASAP7_75t_L g9 ( 
.A(n_10),
.Y(n_9)
);

AOI21xp5_ASAP7_75t_SL g10 ( 
.A1(n_11),
.A2(n_109),
.B(n_130),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_38),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_12),
.B(n_38),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_25),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_13),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_16),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_16),
.B(n_26),
.Y(n_113)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_26),
.B(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_27),
.Y(n_115)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_32),
.B(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_62),
.B1(n_63),
.B2(n_108),
.Y(n_38)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_45),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_46),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_48),
.B(n_87),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_48),
.B(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_52),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_56),
.Y(n_145)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_62),
.B(n_108),
.Y(n_133)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_98),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_75),
.Y(n_64)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_75),
.B(n_100),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_87),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_80),
.B1(n_83),
.B2(n_85),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_79),
.Y(n_86)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_88),
.B(n_157),
.Y(n_156)
);

OAI22x1_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_91),
.B1(n_93),
.B2(n_96),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_116),
.B(n_129),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_112),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_123),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_SL g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_165),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

NOR2x1_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_134),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_141),
.Y(n_134)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_155),
.B1(n_163),
.B2(n_164),
.Y(n_141)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_149),
.B2(n_152),
.Y(n_144)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_162),
.Y(n_155)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);


endmodule