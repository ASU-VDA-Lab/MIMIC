module fake_jpeg_32178_n_541 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_541);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_541;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVxp33_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx8_ASAP7_75t_SL g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx4f_ASAP7_75t_SL g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx2_ASAP7_75t_SL g146 ( 
.A(n_53),
.Y(n_146)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_22),
.B(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_93),
.Y(n_105)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_58),
.Y(n_142)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_60),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_40),
.B(n_8),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_61),
.B(n_77),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_62),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_63),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_64),
.Y(n_145)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_22),
.B(n_8),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_92),
.Y(n_106)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_69),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_70),
.Y(n_151)
);

BUFx4f_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_72),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_76),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_23),
.B(n_20),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_78),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_32),
.B(n_11),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_79),
.B(n_102),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_82),
.Y(n_163)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_83),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_32),
.B(n_11),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_98),
.Y(n_107)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_27),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_104),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_39),
.B(n_11),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_103),
.Y(n_117)
);

AOI21xp33_ASAP7_75t_L g101 ( 
.A1(n_21),
.A2(n_18),
.B(n_7),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_101),
.B(n_0),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_42),
.B(n_7),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_26),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_95),
.A2(n_27),
.B1(n_49),
.B2(n_46),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_116),
.A2(n_130),
.B1(n_135),
.B2(n_150),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_57),
.A2(n_47),
.B1(n_43),
.B2(n_42),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_118),
.A2(n_127),
.B1(n_45),
.B2(n_38),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_123),
.A2(n_37),
.B(n_24),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_74),
.A2(n_43),
.B1(n_47),
.B2(n_19),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_125),
.B(n_37),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_58),
.A2(n_26),
.B1(n_49),
.B2(n_46),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_61),
.B(n_50),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_128),
.B(n_129),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_53),
.B(n_50),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_88),
.A2(n_50),
.B1(n_30),
.B2(n_19),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_19),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_134),
.B(n_152),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_87),
.A2(n_27),
.B1(n_49),
.B2(n_26),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_80),
.B(n_30),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_141),
.B(n_164),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_64),
.A2(n_27),
.B1(n_104),
.B2(n_65),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_98),
.B(n_30),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_55),
.A2(n_26),
.B1(n_45),
.B2(n_38),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_155),
.A2(n_158),
.B1(n_33),
.B2(n_36),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_62),
.A2(n_49),
.B1(n_45),
.B2(n_24),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_69),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_165),
.Y(n_251)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_166),
.Y(n_245)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_120),
.Y(n_168)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_168),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_146),
.Y(n_169)
);

INVx13_ASAP7_75t_L g257 ( 
.A(n_169),
.Y(n_257)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_170),
.Y(n_243)
);

INVx11_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

INVx11_ASAP7_75t_L g241 ( 
.A(n_171),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_172),
.B(n_173),
.Y(n_224)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_110),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_174),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_105),
.B(n_80),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_175),
.B(n_178),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_117),
.B(n_106),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_177),
.B(n_208),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_94),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_112),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_179),
.B(n_190),
.Y(n_227)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_180),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_148),
.A2(n_96),
.B1(n_63),
.B2(n_89),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_181),
.A2(n_191),
.B1(n_109),
.B2(n_156),
.Y(n_248)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_183),
.Y(n_247)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_184),
.Y(n_253)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_185),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_153),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_186),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_187),
.B(n_192),
.Y(n_230)
);

INVx5_ASAP7_75t_SL g188 ( 
.A(n_144),
.Y(n_188)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_188),
.Y(n_260)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_189),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_143),
.B(n_94),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_158),
.A2(n_76),
.B1(n_72),
.B2(n_84),
.Y(n_191)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_139),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_193),
.Y(n_239)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_139),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_194),
.Y(n_254)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_131),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_195),
.B(n_196),
.Y(n_232)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_147),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_137),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_197),
.B(n_198),
.Y(n_259)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_111),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_121),
.A2(n_59),
.B(n_71),
.Y(n_199)
);

NAND2x1_ASAP7_75t_L g262 ( 
.A(n_199),
.B(n_41),
.Y(n_262)
);

AO22x1_ASAP7_75t_L g200 ( 
.A1(n_127),
.A2(n_49),
.B1(n_60),
.B2(n_78),
.Y(n_200)
);

AO22x1_ASAP7_75t_SL g233 ( 
.A1(n_200),
.A2(n_144),
.B1(n_159),
.B2(n_138),
.Y(n_233)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_108),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_201),
.B(n_204),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_161),
.A2(n_86),
.B1(n_24),
.B2(n_38),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_202),
.A2(n_214),
.B1(n_215),
.B2(n_219),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_145),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g256 ( 
.A(n_203),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_121),
.B(n_41),
.Y(n_204)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_162),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_205),
.B(n_206),
.Y(n_269)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_108),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_140),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_210),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_107),
.B(n_21),
.Y(n_208)
);

AND2x2_ASAP7_75t_SL g209 ( 
.A(n_122),
.B(n_0),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_36),
.Y(n_229)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_115),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_122),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_211),
.B(n_213),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_148),
.B(n_21),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_220),
.Y(n_228)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_145),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_120),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_119),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_124),
.B(n_41),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_217),
.B(n_1),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_150),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_218),
.B(n_223),
.Y(n_234)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_153),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_151),
.B(n_33),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_142),
.A2(n_70),
.B1(n_73),
.B2(n_151),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_221),
.A2(n_157),
.B1(n_156),
.B2(n_109),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_162),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_222),
.A2(n_44),
.B1(n_14),
.B2(n_15),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_135),
.A2(n_33),
.B(n_36),
.C(n_41),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_229),
.B(n_169),
.Y(n_300)
);

OAI32xp33_ASAP7_75t_L g231 ( 
.A1(n_177),
.A2(n_116),
.A3(n_119),
.B1(n_114),
.B2(n_142),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_231),
.B(n_192),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_233),
.B(n_262),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_238),
.A2(n_248),
.B1(n_261),
.B2(n_191),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_157),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_240),
.B(n_249),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_176),
.A2(n_113),
.B1(n_159),
.B2(n_138),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_244),
.A2(n_265),
.B1(n_169),
.B2(n_171),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_167),
.B(n_114),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_113),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_255),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_212),
.B(n_160),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_173),
.A2(n_160),
.B1(n_85),
.B2(n_44),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_182),
.B(n_37),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_263),
.B(n_187),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_208),
.B(n_14),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_266),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_200),
.A2(n_44),
.B1(n_37),
.B2(n_41),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_209),
.B(n_0),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_270),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_272),
.Y(n_299)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_268),
.Y(n_273)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_273),
.Y(n_319)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_268),
.Y(n_274)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_274),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_275),
.B(n_277),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_225),
.B(n_199),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_278),
.A2(n_279),
.B1(n_296),
.B2(n_298),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_224),
.A2(n_200),
.B1(n_192),
.B2(n_221),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_247),
.Y(n_280)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_280),
.Y(n_331)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_247),
.Y(n_282)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_282),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_228),
.B(n_209),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_284),
.B(n_290),
.Y(n_322)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_243),
.Y(n_286)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_286),
.Y(n_356)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_226),
.Y(n_287)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_287),
.Y(n_349)
);

OA22x2_ASAP7_75t_L g348 ( 
.A1(n_288),
.A2(n_314),
.B1(n_253),
.B2(n_237),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_225),
.B(n_249),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_289),
.B(n_305),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_228),
.B(n_172),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_230),
.A2(n_223),
.B1(n_213),
.B2(n_185),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_291),
.B(n_267),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_230),
.B(n_170),
.C(n_166),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_292),
.B(n_316),
.C(n_239),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_245),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_293),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_224),
.A2(n_165),
.B1(n_184),
.B2(n_188),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_294),
.A2(n_302),
.B1(n_312),
.B2(n_271),
.Y(n_321)
);

INVx5_ASAP7_75t_L g295 ( 
.A(n_235),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_313),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_224),
.A2(n_196),
.B1(n_222),
.B2(n_207),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_260),
.A2(n_203),
.B1(n_214),
.B2(n_205),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_297),
.A2(n_304),
.B1(n_315),
.B2(n_256),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_300),
.B(n_229),
.Y(n_338)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_226),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_301),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_261),
.A2(n_210),
.B1(n_193),
.B2(n_194),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_231),
.A2(n_211),
.B1(n_206),
.B2(n_201),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_303),
.A2(n_264),
.B1(n_242),
.B2(n_246),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_260),
.A2(n_168),
.B1(n_195),
.B2(n_215),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_242),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_242),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_306),
.B(n_245),
.Y(n_353)
);

NOR2x1p5_ASAP7_75t_L g307 ( 
.A(n_262),
.B(n_1),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_307),
.B(n_309),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_234),
.A2(n_12),
.B(n_17),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_308),
.A2(n_263),
.B(n_266),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_240),
.B(n_12),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_252),
.B(n_1),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_311),
.B(n_269),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_234),
.A2(n_12),
.B1(n_17),
.B2(n_16),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_243),
.Y(n_313)
);

OA21x2_ASAP7_75t_L g314 ( 
.A1(n_233),
.A2(n_1),
.B(n_2),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_237),
.A2(n_14),
.B1(n_17),
.B2(n_16),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_230),
.B(n_5),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_318),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_288),
.A2(n_255),
.B1(n_258),
.B2(n_233),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_320),
.A2(n_321),
.B1(n_325),
.B2(n_326),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_323),
.A2(n_337),
.B(n_343),
.Y(n_363)
);

OAI22xp33_ASAP7_75t_L g325 ( 
.A1(n_285),
.A2(n_233),
.B1(n_248),
.B2(n_262),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_290),
.A2(n_238),
.B1(n_250),
.B2(n_227),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_328),
.A2(n_340),
.B1(n_346),
.B2(n_305),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_289),
.B(n_236),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_332),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_278),
.A2(n_250),
.B1(n_236),
.B2(n_235),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_333),
.B(n_339),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_310),
.A2(n_272),
.B(n_246),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_334),
.A2(n_308),
.B(n_277),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_307),
.A2(n_246),
.B(n_232),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_338),
.B(n_283),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_279),
.A2(n_259),
.B1(n_271),
.B2(n_254),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_341),
.B(n_300),
.Y(n_369)
);

AND2x4_ASAP7_75t_L g343 ( 
.A(n_307),
.B(n_257),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_314),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_345),
.B(n_352),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_310),
.A2(n_239),
.B1(n_254),
.B2(n_245),
.Y(n_346)
);

AND2x4_ASAP7_75t_L g347 ( 
.A(n_310),
.B(n_257),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_347),
.A2(n_296),
.B(n_280),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_348),
.A2(n_354),
.B1(n_324),
.B2(n_340),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_350),
.Y(n_385)
);

AO22x1_ASAP7_75t_SL g351 ( 
.A1(n_314),
.A2(n_243),
.B1(n_251),
.B2(n_253),
.Y(n_351)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_351),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_299),
.B(n_256),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_353),
.B(n_293),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_291),
.A2(n_281),
.B1(n_294),
.B2(n_276),
.Y(n_354)
);

BUFx24_ASAP7_75t_SL g355 ( 
.A(n_275),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_355),
.Y(n_364)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_319),
.Y(n_359)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_359),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_329),
.B(n_301),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_360),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_361),
.A2(n_362),
.B1(n_379),
.B2(n_384),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_341),
.B(n_284),
.C(n_292),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_365),
.B(n_369),
.C(n_372),
.Y(n_407)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_319),
.Y(n_366)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_366),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_329),
.B(n_287),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_367),
.Y(n_409)
);

AO21x1_ASAP7_75t_L g404 ( 
.A1(n_368),
.A2(n_337),
.B(n_380),
.Y(n_404)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_330),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_370),
.B(n_373),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_338),
.B(n_322),
.C(n_354),
.Y(n_372)
);

INVx8_ASAP7_75t_L g374 ( 
.A(n_348),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_374),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_322),
.B(n_276),
.C(n_281),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_375),
.B(n_376),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_323),
.B(n_316),
.C(n_283),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_324),
.A2(n_314),
.B1(n_302),
.B2(n_312),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_323),
.A2(n_306),
.B(n_309),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_380),
.A2(n_327),
.B(n_318),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_339),
.B(n_311),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_381),
.B(n_382),
.Y(n_406)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_330),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_383),
.B(n_369),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_345),
.A2(n_348),
.B1(n_320),
.B2(n_328),
.Y(n_384)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_331),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_386),
.B(n_389),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_336),
.B(n_282),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_387),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_388),
.A2(n_391),
.B(n_353),
.Y(n_396)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_331),
.Y(n_389)
);

XOR2x2_ASAP7_75t_L g391 ( 
.A(n_343),
.B(n_298),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_378),
.A2(n_342),
.B1(n_335),
.B2(n_326),
.Y(n_393)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_393),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_390),
.A2(n_335),
.B1(n_327),
.B2(n_336),
.Y(n_395)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_395),
.Y(n_444)
);

AO22x1_ASAP7_75t_L g445 ( 
.A1(n_396),
.A2(n_366),
.B1(n_359),
.B2(n_385),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_398),
.B(n_402),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g400 ( 
.A(n_372),
.B(n_333),
.Y(n_400)
);

XNOR2x1_ASAP7_75t_L g441 ( 
.A(n_400),
.B(n_360),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_365),
.B(n_334),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_401),
.B(n_376),
.C(n_377),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_362),
.A2(n_348),
.B1(n_321),
.B2(n_351),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_403),
.A2(n_414),
.B1(n_415),
.B2(n_418),
.Y(n_434)
);

OAI21xp33_ASAP7_75t_SL g428 ( 
.A1(n_404),
.A2(n_388),
.B(n_391),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_357),
.A2(n_346),
.B1(n_351),
.B2(n_347),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_408),
.A2(n_313),
.B1(n_241),
.B2(n_256),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_383),
.B(n_347),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_410),
.B(n_398),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_363),
.A2(n_347),
.B(n_343),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_413),
.A2(n_417),
.B(n_423),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_384),
.A2(n_357),
.B1(n_374),
.B2(n_379),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_374),
.A2(n_351),
.B1(n_347),
.B2(n_343),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_377),
.Y(n_416)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_416),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_363),
.A2(n_343),
.B(n_349),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_371),
.A2(n_349),
.B1(n_344),
.B2(n_273),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_361),
.A2(n_344),
.B1(n_274),
.B2(n_356),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_421),
.A2(n_389),
.B1(n_386),
.B2(n_382),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_387),
.B(n_317),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_422),
.B(n_373),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_358),
.A2(n_356),
.B(n_256),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_405),
.B(n_375),
.Y(n_424)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_424),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_426),
.B(n_433),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_405),
.B(n_364),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_427),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_428),
.A2(n_429),
.B1(n_408),
.B2(n_415),
.Y(n_451)
);

OAI22xp33_ASAP7_75t_L g429 ( 
.A1(n_412),
.A2(n_391),
.B1(n_358),
.B2(n_390),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_422),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_430),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_431),
.B(n_447),
.Y(n_462)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_412),
.Y(n_435)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_435),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_409),
.B(n_364),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_436),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_420),
.B(n_367),
.Y(n_437)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_437),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_409),
.B(n_420),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_438),
.Y(n_469)
);

MAJx2_ASAP7_75t_L g439 ( 
.A(n_407),
.B(n_368),
.C(n_381),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_439),
.B(n_441),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_440),
.A2(n_411),
.B1(n_394),
.B2(n_413),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_399),
.B(n_370),
.Y(n_442)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_442),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_445),
.A2(n_418),
.B(n_423),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_407),
.B(n_251),
.C(n_286),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_446),
.B(n_392),
.C(n_401),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_406),
.B(n_295),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_399),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_448),
.B(n_419),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_450),
.A2(n_403),
.B1(n_421),
.B2(n_414),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_451),
.A2(n_463),
.B1(n_472),
.B2(n_444),
.Y(n_478)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_454),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_458),
.C(n_433),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_457),
.A2(n_429),
.B1(n_434),
.B2(n_445),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_446),
.B(n_426),
.C(n_439),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_443),
.A2(n_397),
.B1(n_410),
.B2(n_396),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_445),
.A2(n_417),
.B(n_397),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_464),
.B(n_467),
.Y(n_484)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_465),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_441),
.B(n_392),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_425),
.B(n_400),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_470),
.B(n_404),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_474),
.B(n_453),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_475),
.A2(n_486),
.B1(n_489),
.B2(n_472),
.Y(n_491)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_460),
.Y(n_477)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_477),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_478),
.A2(n_464),
.B1(n_454),
.B2(n_463),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_459),
.B(n_437),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_479),
.B(n_480),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g480 ( 
.A(n_465),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_462),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_481),
.B(n_482),
.Y(n_505)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_460),
.Y(n_482)
);

XNOR2x1_ASAP7_75t_L g483 ( 
.A(n_466),
.B(n_458),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_483),
.B(n_485),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_470),
.B(n_425),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_457),
.A2(n_434),
.B1(n_448),
.B2(n_440),
.Y(n_486)
);

NAND3xp33_ASAP7_75t_L g487 ( 
.A(n_455),
.B(n_469),
.C(n_468),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_487),
.B(n_431),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_488),
.B(n_484),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_461),
.A2(n_435),
.B1(n_471),
.B2(n_449),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_473),
.A2(n_461),
.B1(n_471),
.B2(n_451),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_490),
.A2(n_241),
.B1(n_257),
.B2(n_14),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_491),
.B(n_496),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_474),
.B(n_456),
.C(n_453),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_492),
.B(n_504),
.C(n_485),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_493),
.B(n_442),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_494),
.A2(n_499),
.B(n_419),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_479),
.B(n_488),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_497),
.B(n_501),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_484),
.A2(n_452),
.B(n_432),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_489),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_475),
.A2(n_450),
.B1(n_462),
.B2(n_452),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_502),
.A2(n_411),
.B1(n_394),
.B2(n_404),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_503),
.B(n_478),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_483),
.B(n_466),
.C(n_467),
.Y(n_504)
);

A2O1A1Ixp33_ASAP7_75t_SL g507 ( 
.A1(n_490),
.A2(n_432),
.B(n_486),
.C(n_476),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_507),
.B(n_511),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_509),
.B(n_510),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_500),
.B(n_406),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_512),
.A2(n_516),
.B1(n_501),
.B2(n_491),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_513),
.B(n_514),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_492),
.B(n_402),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_515),
.A2(n_498),
.B1(n_5),
.B2(n_16),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_503),
.B(n_2),
.C(n_3),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_517),
.B(n_495),
.C(n_505),
.Y(n_520)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_520),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_521),
.B(n_522),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_512),
.A2(n_493),
.B1(n_498),
.B2(n_504),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_523),
.B(n_507),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_509),
.B(n_2),
.C(n_3),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_517),
.C(n_508),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_526),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_518),
.A2(n_506),
.B(n_507),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_527),
.A2(n_522),
.B(n_524),
.Y(n_533)
);

NOR2x1_ASAP7_75t_L g532 ( 
.A(n_529),
.B(n_521),
.Y(n_532)
);

OAI321xp33_ASAP7_75t_L g534 ( 
.A1(n_532),
.A2(n_533),
.A3(n_530),
.B1(n_519),
.B2(n_528),
.C(n_507),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_534),
.B(n_535),
.C(n_530),
.Y(n_536)
);

BUFx24_ASAP7_75t_SL g535 ( 
.A(n_531),
.Y(n_535)
);

AOI322xp5_ASAP7_75t_L g537 ( 
.A1(n_536),
.A2(n_519),
.A3(n_525),
.B1(n_520),
.B2(n_5),
.C1(n_18),
.C2(n_4),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_18),
.C(n_3),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_538),
.B(n_2),
.C(n_3),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_SL g540 ( 
.A1(n_539),
.A2(n_4),
.B(n_500),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_540),
.B(n_4),
.C(n_455),
.Y(n_541)
);


endmodule