module fake_jpeg_25466_n_170 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_170);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_45),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_19),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_6),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_2),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_27),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_53),
.Y(n_90)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_0),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_66),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

BUFx4f_ASAP7_75t_SL g89 ( 
.A(n_82),
.Y(n_89)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_83),
.A2(n_72),
.B1(n_54),
.B2(n_69),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_78),
.B1(n_56),
.B2(n_70),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_91),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_55),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_76),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_92),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_93),
.B(n_60),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_82),
.A2(n_49),
.B1(n_74),
.B2(n_50),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_94),
.A2(n_61),
.B1(n_52),
.B2(n_58),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_82),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_95),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_97),
.A2(n_87),
.B1(n_96),
.B2(n_59),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_103),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_93),
.A2(n_51),
.B1(n_64),
.B2(n_70),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_107),
.B(n_75),
.Y(n_121)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_108),
.Y(n_111)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_56),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_89),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_101),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_117),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_96),
.Y(n_131)
);

AOI21xp33_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_94),
.B(n_79),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_119),
.C(n_116),
.Y(n_127)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_73),
.Y(n_119)
);

OAI32xp33_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_75),
.A3(n_73),
.B1(n_59),
.B2(n_57),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_121),
.B1(n_71),
.B2(n_2),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_122),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_130),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_132),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_123),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_129),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_97),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_131),
.B(n_134),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_116),
.A2(n_108),
.B1(n_71),
.B2(n_3),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_133),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_139)
);

AO22x1_ASAP7_75t_SL g134 ( 
.A1(n_122),
.A2(n_23),
.B1(n_46),
.B2(n_42),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_135),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_125),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_136),
.A2(n_139),
.B1(n_147),
.B2(n_15),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_79),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_144),
.Y(n_154)
);

OA21x2_ASAP7_75t_L g141 ( 
.A1(n_134),
.A2(n_7),
.B(n_8),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_141),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_131),
.B(n_9),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_138),
.C(n_141),
.Y(n_156)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_124),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_146),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_129),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_150),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_17),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_151),
.A2(n_156),
.B(n_138),
.Y(n_158)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_155),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_158),
.A2(n_145),
.B1(n_153),
.B2(n_152),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_157),
.C(n_145),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_154),
.C(n_151),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_162),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_159),
.B(n_21),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_20),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_24),
.C(n_25),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_166),
.B(n_26),
.Y(n_167)
);

O2A1O1Ixp33_ASAP7_75t_SL g168 ( 
.A1(n_167),
.A2(n_29),
.B(n_30),
.C(n_32),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_168),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_38),
.Y(n_170)
);


endmodule