module real_aes_4794_n_7 (n_4, n_0, n_3, n_5, n_2, n_6, n_1, n_7);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_6;
input n_1;
output n_7;
wire n_17;
wire n_22;
wire n_13;
wire n_12;
wire n_19;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_23;
wire n_9;
wire n_20;
wire n_18;
wire n_21;
wire n_8;
wire n_10;
AOI32xp33_ASAP7_75t_L g7 ( .A1(n_0), .A2(n_8), .A3(n_10), .B1(n_13), .B2(n_15), .Y(n_7) );
OAI321xp33_ASAP7_75t_L g15 ( .A1(n_0), .A2(n_10), .A3(n_11), .B1(n_14), .B2(n_16), .C(n_23), .Y(n_15) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_1), .Y(n_14) );
BUFx6f_ASAP7_75t_L g20 ( .A(n_2), .Y(n_20) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_3), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_4), .Y(n_21) );
HB1xp67_ASAP7_75t_L g9 ( .A(n_5), .Y(n_9) );
INVx1_ASAP7_75t_L g12 ( .A(n_6), .Y(n_12) );
NOR2xp33_ASAP7_75t_L g8 ( .A(n_9), .B(n_10), .Y(n_8) );
CKINVDCx20_ASAP7_75t_R g23 ( .A(n_9), .Y(n_23) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_11), .Y(n_10) );
HB1xp67_ASAP7_75t_L g11 ( .A(n_12), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_14), .Y(n_13) );
AOI22xp5_ASAP7_75t_L g16 ( .A1(n_17), .A2(n_18), .B1(n_21), .B2(n_22), .Y(n_16) );
INVx2_ASAP7_75t_SL g17 ( .A(n_18), .Y(n_17) );
BUFx2_ASAP7_75t_L g18 ( .A(n_19), .Y(n_18) );
HB1xp67_ASAP7_75t_L g19 ( .A(n_20), .Y(n_19) );
endmodule