module real_jpeg_12757_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_230, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_230;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_205;
wire n_110;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_202;
wire n_213;
wire n_128;
wire n_179;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_43),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_2),
.A2(n_43),
.B1(n_51),
.B2(n_52),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_2),
.A2(n_43),
.B1(n_61),
.B2(n_62),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_2),
.A2(n_22),
.B1(n_28),
.B2(n_43),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_2),
.A2(n_8),
.B(n_51),
.C(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_2),
.B(n_71),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_2),
.B(n_22),
.C(n_38),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_2),
.B(n_48),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_2),
.B(n_52),
.C(n_67),
.Y(n_190)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_5),
.A2(n_22),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_5),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_7),
.A2(n_22),
.B1(n_28),
.B2(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_7),
.A2(n_31),
.B1(n_35),
.B2(n_36),
.Y(n_117)
);

AO22x1_ASAP7_75t_L g48 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_9),
.Y(n_67)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_11),
.A2(n_35),
.B1(n_36),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_11),
.A2(n_41),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_11),
.A2(n_41),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_11),
.A2(n_22),
.B1(n_28),
.B2(n_41),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_123),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_122),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_100),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_16),
.B(n_100),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_74),
.C(n_84),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_17),
.B(n_74),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_44),
.B2(n_45),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_18),
.B(n_46),
.C(n_73),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_32),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_20),
.A2(n_32),
.B1(n_148),
.B2(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_20),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_25),
.B1(n_27),
.B2(n_30),
.Y(n_20)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_21),
.A2(n_25),
.B1(n_90),
.B2(n_142),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

INVx3_ASAP7_75t_SL g28 ( 
.A(n_22),
.Y(n_28)
);

AO22x1_ASAP7_75t_L g39 ( 
.A1(n_22),
.A2(n_28),
.B1(n_37),
.B2(n_38),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_25),
.A2(n_27),
.B(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_25),
.A2(n_88),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_25),
.B(n_43),
.Y(n_169)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_26),
.B(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_28),
.B(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_30),
.B(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_32),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_32),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_32),
.A2(n_148),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_32),
.B(n_158),
.C(n_160),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_32),
.B(n_135),
.C(n_147),
.Y(n_183)
);

AO22x1_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_33),
.B(n_42),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_33),
.A2(n_39),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_33),
.Y(n_196)
);

NOR2x1_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_39),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_35),
.B(n_154),
.Y(n_153)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_SL g132 ( 
.A1(n_36),
.A2(n_43),
.B(n_49),
.Y(n_132)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_42),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_43),
.B(n_80),
.Y(n_171)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_58),
.B1(n_72),
.B2(n_73),
.Y(n_45)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_46),
.A2(n_72),
.B1(n_91),
.B2(n_92),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_46),
.A2(n_72),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_46),
.B(n_97),
.C(n_195),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B(n_54),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_47),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_47),
.A2(n_50),
.B1(n_95),
.B2(n_96),
.Y(n_119)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

O2A1O1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_49),
.B(n_52),
.C(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_52),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_51),
.A2(n_52),
.B1(n_67),
.B2(n_68),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_58),
.A2(n_73),
.B1(n_118),
.B2(n_119),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_58),
.B(n_118),
.C(n_202),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_65),
.B1(n_70),
.B2(n_71),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OA21x2_ASAP7_75t_L g98 ( 
.A1(n_60),
.A2(n_69),
.B(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_61),
.A2(n_62),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_62),
.B(n_190),
.Y(n_189)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_70),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_65),
.B(n_71),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

INVxp33_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_72),
.B(n_92),
.C(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_78),
.B1(n_79),
.B2(n_83),
.Y(n_74)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_79),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_75),
.A2(n_83),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_76),
.B(n_90),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B(n_82),
.Y(n_79)
);

OA21x2_ASAP7_75t_L g92 ( 
.A1(n_80),
.A2(n_82),
.B(n_93),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_80),
.A2(n_196),
.B(n_197),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_84),
.B(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_94),
.C(n_97),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_85),
.A2(n_86),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_87),
.A2(n_91),
.B1(n_92),
.B2(n_205),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_87),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_91),
.A2(n_92),
.B1(n_153),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_92),
.B(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_94),
.A2(n_97),
.B1(n_98),
.B2(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_94),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_97),
.A2(n_98),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_121),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_112),
.B2(n_113),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_118),
.B(n_120),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_114),
.B(n_118),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_119),
.B1(n_137),
.B2(n_143),
.Y(n_136)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_119),
.B(n_138),
.C(n_141),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_223),
.B(n_227),
.Y(n_123)
);

OAI321xp33_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_199),
.A3(n_218),
.B1(n_221),
.B2(n_222),
.C(n_230),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_182),
.B(n_198),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_149),
.B(n_181),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_134),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_128),
.B(n_134),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_129),
.A2(n_130),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_133),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_144),
.B2(n_145),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_140),
.B(n_164),
.Y(n_173)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_141),
.B(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_146),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_175),
.B(n_180),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_162),
.B(n_174),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_152),
.B(n_155),
.Y(n_174)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_155)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_156),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_157),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_159),
.A2(n_160),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_160),
.B(n_171),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_188),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_166),
.B(n_173),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_170),
.B(n_172),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_176),
.B(n_177),
.Y(n_180)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_183),
.B(n_184),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_191),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_187),
.C(n_191),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_207),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_207),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.C(n_206),
.Y(n_200)
);

FAx1_ASAP7_75t_SL g220 ( 
.A(n_201),
.B(n_204),
.CI(n_206),
.CON(n_220),
.SN(n_220)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_217),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_214),
.B2(n_215),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_215),
.C(n_217),
.Y(n_226)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_219),
.B(n_220),
.Y(n_221)
);

BUFx24_ASAP7_75t_SL g229 ( 
.A(n_220),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_224),
.B(n_226),
.Y(n_227)
);


endmodule