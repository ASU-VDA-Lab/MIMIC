module fake_jpeg_3303_n_150 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_150);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx11_ASAP7_75t_SL g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_7),
.B(n_34),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_19),
.B(n_23),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_58),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_60),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_1),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_60),
.B(n_41),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_45),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_56),
.A2(n_44),
.B1(n_50),
.B2(n_49),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_42),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_44),
.B1(n_40),
.B2(n_50),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_71),
.B1(n_59),
.B2(n_58),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_54),
.A2(n_49),
.B1(n_42),
.B2(n_37),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_41),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_75),
.Y(n_86)
);

NAND2xp33_ASAP7_75t_SL g74 ( 
.A(n_62),
.B(n_59),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_61),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_48),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_77),
.A2(n_81),
.B1(n_68),
.B2(n_58),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_67),
.Y(n_79)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_57),
.Y(n_98)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

OAI32xp33_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_37),
.A3(n_48),
.B1(n_52),
.B2(n_59),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_61),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_93),
.B1(n_95),
.B2(n_74),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_83),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_79),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_57),
.B1(n_56),
.B2(n_68),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_46),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_97),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_38),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_104),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_81),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_31),
.C(n_29),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_97),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_105),
.A2(n_21),
.B1(n_5),
.B2(n_6),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_113),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_76),
.B(n_84),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_109),
.A2(n_26),
.B(n_24),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_91),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_110),
.B(n_111),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_86),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_112),
.Y(n_126)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_2),
.Y(n_120)
);

AOI322xp5_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_38),
.A3(n_51),
.B1(n_17),
.B2(n_22),
.C1(n_33),
.C2(n_32),
.Y(n_115)
);

AOI221xp5_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_123),
.B1(n_107),
.B2(n_9),
.C(n_10),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_106),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_121),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_122),
.C(n_11),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_8),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_106),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_108),
.B(n_27),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_127),
.B1(n_123),
.B2(n_119),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_103),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_SL g134 ( 
.A1(n_129),
.A2(n_105),
.B(n_10),
.C(n_11),
.Y(n_134)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_131),
.B(n_132),
.Y(n_140)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

NOR4xp25_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_134),
.C(n_129),
.D(n_13),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_137),
.Y(n_138)
);

NOR3xp33_ASAP7_75t_SL g141 ( 
.A(n_136),
.B(n_125),
.C(n_118),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_139),
.A2(n_141),
.B1(n_134),
.B2(n_124),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_138),
.B(n_122),
.C(n_130),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_142),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_128),
.C(n_116),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_144),
.B(n_134),
.Y(n_146)
);

NOR2xp67_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_143),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_12),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_12),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_13),
.Y(n_150)
);


endmodule