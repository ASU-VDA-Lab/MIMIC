module real_aes_7501_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_746;
wire n_153;
wire n_532;
wire n_284;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_741;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g270 ( .A1(n_0), .A2(n_271), .B(n_272), .C(n_275), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_1), .B(n_259), .Y(n_276) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_2), .B(n_90), .C(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g122 ( .A(n_2), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_3), .B(n_187), .Y(n_186) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_4), .A2(n_148), .B(n_151), .C(n_531), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_5), .A2(n_143), .B(n_555), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_6), .A2(n_143), .B(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_7), .B(n_259), .Y(n_561) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_8), .A2(n_178), .B(n_215), .Y(n_214) );
AND2x6_ASAP7_75t_L g148 ( .A(n_9), .B(n_149), .Y(n_148) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_10), .A2(n_148), .B(n_151), .C(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g499 ( .A(n_11), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_12), .B(n_107), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_12), .B(n_40), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_13), .B(n_235), .Y(n_533) );
INVx1_ASAP7_75t_L g169 ( .A(n_14), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_15), .B(n_187), .Y(n_221) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_16), .A2(n_188), .B(n_517), .C(n_519), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_17), .B(n_259), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_18), .B(n_163), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g150 ( .A1(n_19), .A2(n_151), .B(n_154), .C(n_162), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_20), .A2(n_223), .B(n_274), .C(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_21), .B(n_235), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_22), .A2(n_55), .B1(n_754), .B2(n_755), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_22), .Y(n_754) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_23), .B(n_235), .Y(n_472) );
CKINVDCx16_ASAP7_75t_R g546 ( .A(n_24), .Y(n_546) );
INVx1_ASAP7_75t_L g471 ( .A(n_25), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_26), .A2(n_151), .B(n_162), .C(n_218), .Y(n_217) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_27), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_28), .Y(n_529) );
INVx1_ASAP7_75t_L g487 ( .A(n_29), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_30), .A2(n_143), .B(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g146 ( .A(n_31), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g199 ( .A1(n_32), .A2(n_191), .B(n_200), .C(n_202), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_33), .Y(n_536) );
A2O1A1Ixp33_ASAP7_75t_L g557 ( .A1(n_34), .A2(n_274), .B(n_558), .C(n_560), .Y(n_557) );
INVxp67_ASAP7_75t_L g488 ( .A(n_35), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_36), .B(n_220), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_37), .A2(n_151), .B(n_162), .C(n_470), .Y(n_469) );
CKINVDCx14_ASAP7_75t_R g556 ( .A(n_38), .Y(n_556) );
AOI222xp33_ASAP7_75t_SL g125 ( .A1(n_39), .A2(n_126), .B1(n_132), .B2(n_738), .C1(n_739), .C2(n_743), .Y(n_125) );
INVx1_ASAP7_75t_L g107 ( .A(n_40), .Y(n_107) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_41), .A2(n_275), .B(n_497), .C(n_498), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_42), .B(n_142), .Y(n_141) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_43), .A2(n_104), .B1(n_112), .B2(n_758), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_44), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_45), .B(n_187), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_46), .B(n_143), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_47), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_48), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_49), .A2(n_191), .B(n_200), .C(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g273 ( .A(n_50), .Y(n_273) );
OAI22xp5_ASAP7_75t_SL g751 ( .A1(n_51), .A2(n_752), .B1(n_753), .B2(n_756), .Y(n_751) );
CKINVDCx16_ASAP7_75t_R g756 ( .A(n_51), .Y(n_756) );
INVx1_ASAP7_75t_L g245 ( .A(n_52), .Y(n_245) );
INVx1_ASAP7_75t_L g505 ( .A(n_53), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_54), .B(n_143), .Y(n_242) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_55), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g171 ( .A(n_56), .Y(n_171) );
CKINVDCx14_ASAP7_75t_R g495 ( .A(n_57), .Y(n_495) );
INVx1_ASAP7_75t_L g149 ( .A(n_58), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_59), .B(n_143), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_60), .B(n_259), .Y(n_258) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_61), .A2(n_161), .B(n_184), .C(n_256), .Y(n_255) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_62), .Y(n_124) );
INVx1_ASAP7_75t_L g168 ( .A(n_63), .Y(n_168) );
OAI22xp5_ASAP7_75t_L g127 ( .A1(n_64), .A2(n_102), .B1(n_128), .B2(n_129), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_64), .Y(n_129) );
INVx1_ASAP7_75t_SL g559 ( .A(n_65), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_66), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_67), .B(n_187), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_68), .B(n_259), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_69), .B(n_188), .Y(n_233) );
INVx1_ASAP7_75t_L g549 ( .A(n_70), .Y(n_549) );
CKINVDCx16_ASAP7_75t_R g269 ( .A(n_71), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_72), .B(n_156), .Y(n_155) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_73), .A2(n_151), .B(n_182), .C(n_191), .Y(n_181) );
CKINVDCx16_ASAP7_75t_R g254 ( .A(n_74), .Y(n_254) );
INVx1_ASAP7_75t_L g111 ( .A(n_75), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_76), .A2(n_143), .B(n_494), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_77), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_78), .A2(n_143), .B(n_514), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_79), .A2(n_142), .B(n_483), .Y(n_482) );
CKINVDCx16_ASAP7_75t_R g468 ( .A(n_80), .Y(n_468) );
INVx1_ASAP7_75t_L g515 ( .A(n_81), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_82), .B(n_159), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_83), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_84), .A2(n_143), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g518 ( .A(n_85), .Y(n_518) );
INVx2_ASAP7_75t_L g166 ( .A(n_86), .Y(n_166) );
INVx1_ASAP7_75t_L g532 ( .A(n_87), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_88), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_89), .B(n_235), .Y(n_234) );
OR2x2_ASAP7_75t_L g119 ( .A(n_90), .B(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g460 ( .A(n_90), .B(n_121), .Y(n_460) );
INVx2_ASAP7_75t_L g737 ( .A(n_90), .Y(n_737) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_91), .A2(n_127), .B1(n_130), .B2(n_131), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_91), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g547 ( .A1(n_92), .A2(n_151), .B(n_191), .C(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_93), .B(n_143), .Y(n_198) );
INVx1_ASAP7_75t_L g203 ( .A(n_94), .Y(n_203) );
INVxp67_ASAP7_75t_L g257 ( .A(n_95), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_96), .B(n_178), .Y(n_500) );
INVx2_ASAP7_75t_L g508 ( .A(n_97), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_98), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g183 ( .A(n_99), .Y(n_183) );
INVx1_ASAP7_75t_L g229 ( .A(n_100), .Y(n_229) );
AND2x2_ASAP7_75t_L g247 ( .A(n_101), .B(n_165), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_102), .Y(n_128) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
CKINVDCx6p67_ASAP7_75t_R g759 ( .A(n_105), .Y(n_759) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
AOI22x1_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_125), .B1(n_746), .B2(n_748), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_114), .B(n_117), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g747 ( .A(n_116), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g748 ( .A1(n_117), .A2(n_749), .B(n_757), .Y(n_748) );
NOR2xp33_ASAP7_75t_SL g117 ( .A(n_118), .B(n_124), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g757 ( .A(n_119), .Y(n_757) );
NOR2x2_ASAP7_75t_L g745 ( .A(n_120), .B(n_737), .Y(n_745) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g736 ( .A(n_121), .B(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
INVx1_ASAP7_75t_L g738 ( .A(n_126), .Y(n_738) );
INVx1_ASAP7_75t_L g130 ( .A(n_127), .Y(n_130) );
OAI22xp5_ASAP7_75t_SL g132 ( .A1(n_133), .A2(n_458), .B1(n_461), .B2(n_734), .Y(n_132) );
OAI22xp5_ASAP7_75t_SL g749 ( .A1(n_133), .A2(n_741), .B1(n_750), .B2(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
BUFx2_ASAP7_75t_L g741 ( .A(n_134), .Y(n_741) );
AND3x1_ASAP7_75t_L g134 ( .A(n_135), .B(n_362), .C(n_419), .Y(n_134) );
NOR3xp33_ASAP7_75t_L g135 ( .A(n_136), .B(n_307), .C(n_343), .Y(n_135) );
OAI211xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_209), .B(n_261), .C(n_294), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_173), .Y(n_137) );
HB1xp67_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x4_ASAP7_75t_L g264 ( .A(n_139), .B(n_265), .Y(n_264) );
INVx5_ASAP7_75t_L g293 ( .A(n_139), .Y(n_293) );
AND2x2_ASAP7_75t_L g366 ( .A(n_139), .B(n_282), .Y(n_366) );
AND2x2_ASAP7_75t_L g404 ( .A(n_139), .B(n_310), .Y(n_404) );
AND2x2_ASAP7_75t_L g424 ( .A(n_139), .B(n_266), .Y(n_424) );
OR2x6_ASAP7_75t_L g139 ( .A(n_140), .B(n_170), .Y(n_139) );
AOI21xp5_ASAP7_75t_SL g140 ( .A1(n_141), .A2(n_150), .B(n_163), .Y(n_140) );
BUFx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_148), .Y(n_143) );
NAND2x1p5_ASAP7_75t_L g230 ( .A(n_144), .B(n_148), .Y(n_230) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
INVx1_ASAP7_75t_L g161 ( .A(n_145), .Y(n_161) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g152 ( .A(n_146), .Y(n_152) );
INVx1_ASAP7_75t_L g224 ( .A(n_146), .Y(n_224) );
INVx1_ASAP7_75t_L g153 ( .A(n_147), .Y(n_153) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_147), .Y(n_157) );
INVx3_ASAP7_75t_L g188 ( .A(n_147), .Y(n_188) );
INVx1_ASAP7_75t_L g220 ( .A(n_147), .Y(n_220) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_147), .Y(n_235) );
BUFx3_ASAP7_75t_L g162 ( .A(n_148), .Y(n_162) );
INVx4_ASAP7_75t_SL g192 ( .A(n_148), .Y(n_192) );
INVx5_ASAP7_75t_L g201 ( .A(n_151), .Y(n_201) );
AND2x6_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_152), .Y(n_190) );
BUFx3_ASAP7_75t_L g206 ( .A(n_152), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_158), .B(n_160), .Y(n_154) );
INVx2_ASAP7_75t_L g159 ( .A(n_156), .Y(n_159) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx4_ASAP7_75t_L g185 ( .A(n_157), .Y(n_185) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_159), .A2(n_203), .B(n_204), .C(n_205), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_159), .A2(n_205), .B(n_245), .C(n_246), .Y(n_244) );
O2A1O1Ixp5_ASAP7_75t_L g531 ( .A1(n_159), .A2(n_532), .B(n_533), .C(n_534), .Y(n_531) );
O2A1O1Ixp33_ASAP7_75t_L g548 ( .A1(n_159), .A2(n_534), .B(n_549), .C(n_550), .Y(n_548) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_160), .A2(n_187), .B(n_471), .C(n_472), .Y(n_470) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_161), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_164), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g172 ( .A(n_165), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_165), .A2(n_198), .B(n_199), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_165), .A2(n_242), .B(n_243), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_L g467 ( .A1(n_165), .A2(n_230), .B(n_468), .C(n_469), .Y(n_467) );
OA21x2_ASAP7_75t_L g492 ( .A1(n_165), .A2(n_493), .B(n_500), .Y(n_492) );
AND2x2_ASAP7_75t_SL g165 ( .A(n_166), .B(n_167), .Y(n_165) );
AND2x2_ASAP7_75t_L g179 ( .A(n_166), .B(n_167), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_171), .B(n_172), .Y(n_170) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_172), .A2(n_528), .B(n_535), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_173), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_196), .Y(n_173) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_174), .Y(n_305) );
AND2x2_ASAP7_75t_L g319 ( .A(n_174), .B(n_265), .Y(n_319) );
INVx1_ASAP7_75t_L g342 ( .A(n_174), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_174), .B(n_293), .Y(n_381) );
OR2x2_ASAP7_75t_L g418 ( .A(n_174), .B(n_263), .Y(n_418) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_175), .Y(n_354) );
AND2x2_ASAP7_75t_L g361 ( .A(n_175), .B(n_266), .Y(n_361) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g282 ( .A(n_176), .B(n_266), .Y(n_282) );
BUFx2_ASAP7_75t_L g310 ( .A(n_176), .Y(n_310) );
AO21x2_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_180), .B(n_194), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_177), .B(n_195), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_177), .B(n_208), .Y(n_207) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_177), .A2(n_228), .B(n_236), .Y(n_227) );
INVx3_ASAP7_75t_L g259 ( .A(n_177), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_177), .B(n_474), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_177), .B(n_536), .Y(n_535) );
AO21x2_ASAP7_75t_L g544 ( .A1(n_177), .A2(n_545), .B(n_551), .Y(n_544) );
INVx4_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_178), .A2(n_216), .B(n_217), .Y(n_215) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_178), .Y(n_251) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g238 ( .A(n_179), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_181), .B(n_193), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_186), .C(n_189), .Y(n_182) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
OAI22xp33_ASAP7_75t_L g486 ( .A1(n_185), .A2(n_187), .B1(n_487), .B2(n_488), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_185), .B(n_508), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_185), .B(n_518), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_187), .B(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g271 ( .A(n_187), .Y(n_271) );
INVx5_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_188), .B(n_499), .Y(n_498) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx3_ASAP7_75t_L g560 ( .A(n_190), .Y(n_560) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
O2A1O1Ixp33_ASAP7_75t_L g253 ( .A1(n_192), .A2(n_201), .B(n_254), .C(n_255), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_SL g268 ( .A1(n_192), .A2(n_201), .B(n_269), .C(n_270), .Y(n_268) );
O2A1O1Ixp33_ASAP7_75t_SL g483 ( .A1(n_192), .A2(n_201), .B(n_484), .C(n_485), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_SL g494 ( .A1(n_192), .A2(n_201), .B(n_495), .C(n_496), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_SL g504 ( .A1(n_192), .A2(n_201), .B(n_505), .C(n_506), .Y(n_504) );
O2A1O1Ixp33_ASAP7_75t_SL g514 ( .A1(n_192), .A2(n_201), .B(n_515), .C(n_516), .Y(n_514) );
O2A1O1Ixp33_ASAP7_75t_L g555 ( .A1(n_192), .A2(n_201), .B(n_556), .C(n_557), .Y(n_555) );
INVx5_ASAP7_75t_L g263 ( .A(n_196), .Y(n_263) );
BUFx2_ASAP7_75t_L g286 ( .A(n_196), .Y(n_286) );
AND2x2_ASAP7_75t_L g443 ( .A(n_196), .B(n_297), .Y(n_443) );
OR2x6_ASAP7_75t_L g196 ( .A(n_197), .B(n_207), .Y(n_196) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g275 ( .A(n_206), .Y(n_275) );
INVx1_ASAP7_75t_L g519 ( .A(n_206), .Y(n_519) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NAND2xp33_ASAP7_75t_L g210 ( .A(n_211), .B(n_248), .Y(n_210) );
OAI221xp5_ASAP7_75t_L g343 ( .A1(n_211), .A2(n_344), .B1(n_351), .B2(n_352), .C(n_355), .Y(n_343) );
OR2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_225), .Y(n_211) );
AND2x2_ASAP7_75t_L g249 ( .A(n_212), .B(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_212), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_SL g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g278 ( .A(n_213), .B(n_226), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_213), .B(n_227), .Y(n_288) );
OR2x2_ASAP7_75t_L g299 ( .A(n_213), .B(n_250), .Y(n_299) );
AND2x2_ASAP7_75t_L g302 ( .A(n_213), .B(n_290), .Y(n_302) );
AND2x2_ASAP7_75t_L g318 ( .A(n_213), .B(n_239), .Y(n_318) );
OR2x2_ASAP7_75t_L g334 ( .A(n_213), .B(n_227), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_213), .B(n_250), .Y(n_396) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_214), .B(n_239), .Y(n_388) );
AND2x2_ASAP7_75t_L g391 ( .A(n_214), .B(n_227), .Y(n_391) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_221), .B(n_222), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_222), .A2(n_233), .B(n_234), .Y(n_232) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx3_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
OR2x2_ASAP7_75t_L g312 ( .A(n_225), .B(n_299), .Y(n_312) );
INVx2_ASAP7_75t_L g338 ( .A(n_225), .Y(n_338) );
OR2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_239), .Y(n_225) );
AND2x2_ASAP7_75t_L g260 ( .A(n_226), .B(n_240), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_226), .B(n_250), .Y(n_317) );
OR2x2_ASAP7_75t_L g328 ( .A(n_226), .B(n_240), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_226), .B(n_290), .Y(n_387) );
OAI221xp5_ASAP7_75t_L g420 ( .A1(n_226), .A2(n_421), .B1(n_423), .B2(n_425), .C(n_428), .Y(n_420) );
INVx5_ASAP7_75t_SL g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_227), .B(n_250), .Y(n_359) );
OAI21xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_231), .Y(n_228) );
OAI21xp5_ASAP7_75t_L g528 ( .A1(n_230), .A2(n_529), .B(n_530), .Y(n_528) );
OAI21xp5_ASAP7_75t_L g545 ( .A1(n_230), .A2(n_546), .B(n_547), .Y(n_545) );
INVx4_ASAP7_75t_L g274 ( .A(n_235), .Y(n_274) );
INVx2_ASAP7_75t_L g497 ( .A(n_235), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
INVx2_ASAP7_75t_L g480 ( .A(n_238), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_239), .B(n_290), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_239), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g306 ( .A(n_239), .B(n_278), .Y(n_306) );
OR2x2_ASAP7_75t_L g350 ( .A(n_239), .B(n_250), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_239), .B(n_302), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_239), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g415 ( .A(n_239), .B(n_416), .Y(n_415) );
INVx5_ASAP7_75t_SL g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_SL g279 ( .A(n_240), .B(n_249), .Y(n_279) );
O2A1O1Ixp33_ASAP7_75t_SL g283 ( .A1(n_240), .A2(n_284), .B(n_287), .C(n_291), .Y(n_283) );
OR2x2_ASAP7_75t_L g321 ( .A(n_240), .B(n_317), .Y(n_321) );
OR2x2_ASAP7_75t_L g357 ( .A(n_240), .B(n_299), .Y(n_357) );
OAI311xp33_ASAP7_75t_L g363 ( .A1(n_240), .A2(n_302), .A3(n_364), .B1(n_367), .C1(n_374), .Y(n_363) );
AND2x2_ASAP7_75t_L g414 ( .A(n_240), .B(n_250), .Y(n_414) );
AND2x2_ASAP7_75t_L g422 ( .A(n_240), .B(n_277), .Y(n_422) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_240), .Y(n_440) );
AND2x2_ASAP7_75t_L g457 ( .A(n_240), .B(n_278), .Y(n_457) );
OR2x6_ASAP7_75t_L g240 ( .A(n_241), .B(n_247), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_249), .B(n_260), .Y(n_248) );
AND2x2_ASAP7_75t_L g285 ( .A(n_249), .B(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g441 ( .A(n_249), .Y(n_441) );
AND2x2_ASAP7_75t_L g277 ( .A(n_250), .B(n_278), .Y(n_277) );
INVx3_ASAP7_75t_L g290 ( .A(n_250), .Y(n_290) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_250), .Y(n_333) );
INVxp67_ASAP7_75t_L g372 ( .A(n_250), .Y(n_372) );
OA21x2_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_252), .B(n_258), .Y(n_250) );
OA21x2_ASAP7_75t_L g502 ( .A1(n_251), .A2(n_503), .B(n_509), .Y(n_502) );
OA21x2_ASAP7_75t_L g512 ( .A1(n_251), .A2(n_513), .B(n_520), .Y(n_512) );
OA21x2_ASAP7_75t_L g553 ( .A1(n_251), .A2(n_554), .B(n_561), .Y(n_553) );
OA21x2_ASAP7_75t_L g266 ( .A1(n_259), .A2(n_267), .B(n_276), .Y(n_266) );
AND2x2_ASAP7_75t_L g450 ( .A(n_260), .B(n_298), .Y(n_450) );
AOI221xp5_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_277), .B1(n_279), .B2(n_280), .C(n_283), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_263), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g303 ( .A(n_263), .B(n_293), .Y(n_303) );
AND2x2_ASAP7_75t_L g311 ( .A(n_263), .B(n_265), .Y(n_311) );
OR2x2_ASAP7_75t_L g323 ( .A(n_263), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g341 ( .A(n_263), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g365 ( .A(n_263), .B(n_366), .Y(n_365) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_263), .Y(n_385) );
AND2x2_ASAP7_75t_L g437 ( .A(n_263), .B(n_361), .Y(n_437) );
OAI31xp33_ASAP7_75t_L g445 ( .A1(n_263), .A2(n_314), .A3(n_413), .B(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_264), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_SL g409 ( .A(n_264), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_264), .B(n_418), .Y(n_417) );
AND2x4_ASAP7_75t_L g297 ( .A(n_265), .B(n_293), .Y(n_297) );
INVx1_ASAP7_75t_L g384 ( .A(n_265), .Y(n_384) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g434 ( .A(n_266), .B(n_293), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_274), .B(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g534 ( .A(n_275), .Y(n_534) );
INVx1_ASAP7_75t_SL g444 ( .A(n_277), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_278), .B(n_349), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_279), .A2(n_391), .B1(n_429), .B2(n_432), .Y(n_428) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g292 ( .A(n_282), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g351 ( .A(n_282), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_282), .B(n_303), .Y(n_456) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g426 ( .A(n_285), .B(n_427), .Y(n_426) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_286), .A2(n_345), .B(n_347), .Y(n_344) );
OR2x2_ASAP7_75t_L g352 ( .A(n_286), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g373 ( .A(n_286), .B(n_361), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_286), .B(n_384), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_286), .B(n_424), .Y(n_423) );
OAI221xp5_ASAP7_75t_SL g400 ( .A1(n_287), .A2(n_401), .B1(n_406), .B2(n_409), .C(n_410), .Y(n_400) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
OR2x2_ASAP7_75t_L g377 ( .A(n_288), .B(n_350), .Y(n_377) );
INVx1_ASAP7_75t_L g416 ( .A(n_288), .Y(n_416) );
INVx2_ASAP7_75t_L g392 ( .A(n_289), .Y(n_392) );
INVx1_ASAP7_75t_L g326 ( .A(n_290), .Y(n_326) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g331 ( .A(n_293), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_293), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g360 ( .A(n_293), .B(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g448 ( .A(n_293), .B(n_418), .Y(n_448) );
AOI222xp33_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_298), .B1(n_300), .B2(n_303), .C1(n_304), .C2(n_306), .Y(n_294) );
INVxp67_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g304 ( .A(n_297), .B(n_305), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_297), .A2(n_347), .B1(n_375), .B2(n_376), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_297), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
OAI21xp33_ASAP7_75t_SL g335 ( .A1(n_306), .A2(n_336), .B(n_339), .Y(n_335) );
OAI211xp5_ASAP7_75t_SL g307 ( .A1(n_308), .A2(n_312), .B(n_313), .C(n_335), .Y(n_307) );
INVxp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
AOI221xp5_ASAP7_75t_L g313 ( .A1(n_311), .A2(n_314), .B1(n_319), .B2(n_320), .C(n_322), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_311), .B(n_399), .Y(n_398) );
INVxp67_ASAP7_75t_L g405 ( .A(n_311), .Y(n_405) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
AND2x2_ASAP7_75t_L g407 ( .A(n_316), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g324 ( .A(n_319), .Y(n_324) );
AND2x2_ASAP7_75t_L g330 ( .A(n_319), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_325), .B1(n_329), .B2(n_332), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_326), .B(n_338), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_327), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g427 ( .A(n_331), .Y(n_427) );
AND2x2_ASAP7_75t_L g446 ( .A(n_331), .B(n_361), .Y(n_446) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_338), .B(n_395), .Y(n_454) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_341), .B(n_409), .Y(n_452) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g375 ( .A(n_353), .Y(n_375) );
BUFx2_ASAP7_75t_L g399 ( .A(n_354), .Y(n_399) );
OAI21xp5_ASAP7_75t_SL g355 ( .A1(n_356), .A2(n_358), .B(n_360), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NOR3xp33_ASAP7_75t_L g362 ( .A(n_363), .B(n_378), .C(n_400), .Y(n_362) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OAI21xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_370), .B(n_373), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
A2O1A1Ixp33_ASAP7_75t_SL g378 ( .A1(n_379), .A2(n_382), .B(n_386), .C(n_389), .Y(n_378) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_379), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NOR2xp67_ASAP7_75t_SL g383 ( .A(n_384), .B(n_385), .Y(n_383) );
OR2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
INVx1_ASAP7_75t_SL g408 ( .A(n_388), .Y(n_408) );
OAI21xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_393), .B(n_397), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
AND2x2_ASAP7_75t_L g413 ( .A(n_391), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_403), .B(n_405), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_413), .B1(n_415), .B2(n_417), .Y(n_410) );
INVx2_ASAP7_75t_SL g431 ( .A(n_418), .Y(n_431) );
NOR3xp33_ASAP7_75t_L g419 ( .A(n_420), .B(n_435), .C(n_447), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVxp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVxp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_431), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OAI221xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_438), .B1(n_442), .B2(n_444), .C(n_445), .Y(n_435) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_436), .A2(n_448), .B(n_449), .C(n_451), .Y(n_447) );
INVx1_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
INVxp67_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B1(n_455), .B2(n_457), .Y(n_451) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g740 ( .A(n_459), .Y(n_740) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_SL g742 ( .A(n_461), .Y(n_742) );
OR5x1_ASAP7_75t_L g461 ( .A(n_462), .B(n_628), .C(n_692), .D(n_708), .E(n_723), .Y(n_461) );
NAND4xp25_ASAP7_75t_L g462 ( .A(n_463), .B(n_562), .C(n_589), .D(n_612), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_510), .B(n_521), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_475), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx3_ASAP7_75t_SL g541 ( .A(n_466), .Y(n_541) );
AND2x4_ASAP7_75t_L g575 ( .A(n_466), .B(n_564), .Y(n_575) );
OR2x2_ASAP7_75t_L g585 ( .A(n_466), .B(n_543), .Y(n_585) );
OR2x2_ASAP7_75t_L g631 ( .A(n_466), .B(n_478), .Y(n_631) );
AND2x2_ASAP7_75t_L g645 ( .A(n_466), .B(n_542), .Y(n_645) );
AND2x2_ASAP7_75t_L g688 ( .A(n_466), .B(n_578), .Y(n_688) );
AND2x2_ASAP7_75t_L g695 ( .A(n_466), .B(n_553), .Y(n_695) );
AND2x2_ASAP7_75t_L g714 ( .A(n_466), .B(n_604), .Y(n_714) );
AND2x2_ASAP7_75t_L g732 ( .A(n_466), .B(n_574), .Y(n_732) );
OR2x6_ASAP7_75t_L g466 ( .A(n_467), .B(n_473), .Y(n_466) );
INVx1_ASAP7_75t_L g697 ( .A(n_475), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_491), .Y(n_475) );
AND2x2_ASAP7_75t_L g607 ( .A(n_476), .B(n_542), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_476), .B(n_627), .Y(n_626) );
AOI32xp33_ASAP7_75t_L g640 ( .A1(n_476), .A2(n_641), .A3(n_644), .B1(n_646), .B2(n_650), .Y(n_640) );
AND2x2_ASAP7_75t_L g710 ( .A(n_476), .B(n_604), .Y(n_710) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g574 ( .A(n_478), .B(n_543), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_478), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g616 ( .A(n_478), .B(n_563), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_478), .B(n_695), .Y(n_694) );
AO21x2_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_481), .B(n_489), .Y(n_478) );
INVx1_ASAP7_75t_L g579 ( .A(n_479), .Y(n_579) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OA21x2_ASAP7_75t_L g578 ( .A1(n_482), .A2(n_490), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g581 ( .A(n_491), .B(n_525), .Y(n_581) );
AND2x2_ASAP7_75t_L g657 ( .A(n_491), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_SL g729 ( .A(n_491), .Y(n_729) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_501), .Y(n_491) );
OR2x2_ASAP7_75t_L g524 ( .A(n_492), .B(n_502), .Y(n_524) );
AND2x2_ASAP7_75t_L g538 ( .A(n_492), .B(n_539), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_492), .B(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g588 ( .A(n_492), .Y(n_588) );
AND2x2_ASAP7_75t_L g615 ( .A(n_492), .B(n_502), .Y(n_615) );
BUFx3_ASAP7_75t_L g618 ( .A(n_492), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_492), .B(n_593), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_492), .B(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g569 ( .A(n_501), .Y(n_569) );
AND2x2_ASAP7_75t_L g587 ( .A(n_501), .B(n_567), .Y(n_587) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g598 ( .A(n_502), .B(n_512), .Y(n_598) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_502), .Y(n_611) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_511), .B(n_618), .Y(n_668) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_SL g539 ( .A(n_512), .Y(n_539) );
NAND3xp33_ASAP7_75t_L g586 ( .A(n_512), .B(n_587), .C(n_588), .Y(n_586) );
OR2x2_ASAP7_75t_L g594 ( .A(n_512), .B(n_567), .Y(n_594) );
AND2x2_ASAP7_75t_L g614 ( .A(n_512), .B(n_567), .Y(n_614) );
AND2x2_ASAP7_75t_L g658 ( .A(n_512), .B(n_527), .Y(n_658) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_537), .B(n_540), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_523), .B(n_525), .Y(n_522) );
AND2x2_ASAP7_75t_L g733 ( .A(n_523), .B(n_658), .Y(n_733) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_524), .A2(n_631), .B1(n_673), .B2(n_675), .Y(n_672) );
OR2x2_ASAP7_75t_L g679 ( .A(n_524), .B(n_594), .Y(n_679) );
OR2x2_ASAP7_75t_L g703 ( .A(n_524), .B(n_704), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_524), .B(n_623), .Y(n_716) );
AND2x2_ASAP7_75t_L g609 ( .A(n_525), .B(n_610), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g696 ( .A1(n_525), .A2(n_682), .B(n_697), .Y(n_696) );
AOI32xp33_ASAP7_75t_L g717 ( .A1(n_525), .A2(n_607), .A3(n_718), .B1(n_720), .B2(n_721), .Y(n_717) );
OR2x2_ASAP7_75t_L g728 ( .A(n_525), .B(n_729), .Y(n_728) );
CKINVDCx16_ASAP7_75t_R g525 ( .A(n_526), .Y(n_525) );
OR2x2_ASAP7_75t_L g596 ( .A(n_526), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_526), .B(n_610), .Y(n_675) );
BUFx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx4_ASAP7_75t_L g567 ( .A(n_527), .Y(n_567) );
AND2x2_ASAP7_75t_L g633 ( .A(n_527), .B(n_598), .Y(n_633) );
AND3x2_ASAP7_75t_L g642 ( .A(n_527), .B(n_538), .C(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g568 ( .A(n_539), .B(n_569), .Y(n_568) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_539), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_539), .B(n_567), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
AND2x2_ASAP7_75t_L g563 ( .A(n_541), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g603 ( .A(n_541), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g621 ( .A(n_541), .B(n_553), .Y(n_621) );
AND2x2_ASAP7_75t_L g639 ( .A(n_541), .B(n_543), .Y(n_639) );
OR2x2_ASAP7_75t_L g653 ( .A(n_541), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g699 ( .A(n_541), .B(n_627), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_542), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_553), .Y(n_542) );
AND2x2_ASAP7_75t_L g600 ( .A(n_543), .B(n_578), .Y(n_600) );
OR2x2_ASAP7_75t_L g654 ( .A(n_543), .B(n_578), .Y(n_654) );
AND2x2_ASAP7_75t_L g707 ( .A(n_543), .B(n_564), .Y(n_707) );
INVx2_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
BUFx2_ASAP7_75t_L g605 ( .A(n_544), .Y(n_605) );
AND2x2_ASAP7_75t_L g627 ( .A(n_544), .B(n_553), .Y(n_627) );
INVx2_ASAP7_75t_L g564 ( .A(n_553), .Y(n_564) );
INVx1_ASAP7_75t_L g584 ( .A(n_553), .Y(n_584) );
AOI211xp5_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_565), .B(n_570), .C(n_582), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_563), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g726 ( .A(n_563), .Y(n_726) );
AND2x2_ASAP7_75t_L g604 ( .A(n_564), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_567), .B(n_568), .Y(n_576) );
INVx1_ASAP7_75t_L g661 ( .A(n_567), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_567), .B(n_588), .Y(n_685) );
AND2x2_ASAP7_75t_L g701 ( .A(n_567), .B(n_615), .Y(n_701) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_568), .B(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g592 ( .A(n_569), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_576), .B1(n_577), .B2(n_580), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_573), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_574), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g599 ( .A(n_575), .B(n_600), .Y(n_599) );
AOI221xp5_ASAP7_75t_SL g664 ( .A1(n_575), .A2(n_617), .B1(n_665), .B2(n_670), .C(n_672), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_575), .B(n_638), .Y(n_671) );
INVx1_ASAP7_75t_L g731 ( .A(n_577), .Y(n_731) );
BUFx3_ASAP7_75t_L g638 ( .A(n_578), .Y(n_638) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AOI21xp33_ASAP7_75t_SL g582 ( .A1(n_583), .A2(n_585), .B(n_586), .Y(n_582) );
INVx1_ASAP7_75t_L g647 ( .A(n_584), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_584), .B(n_638), .Y(n_691) );
INVx1_ASAP7_75t_L g648 ( .A(n_585), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_585), .B(n_638), .Y(n_649) );
INVxp67_ASAP7_75t_L g669 ( .A(n_587), .Y(n_669) );
AND2x2_ASAP7_75t_L g610 ( .A(n_588), .B(n_611), .Y(n_610) );
O2A1O1Ixp33_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_595), .B(n_599), .C(n_601), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVx1_ASAP7_75t_SL g624 ( .A(n_592), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_593), .B(n_624), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_593), .B(n_615), .Y(n_666) );
INVx2_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_596), .A2(n_602), .B1(n_606), .B2(n_608), .Y(n_601) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g617 ( .A(n_598), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g662 ( .A(n_598), .B(n_663), .Y(n_662) );
OAI21xp33_ASAP7_75t_L g665 ( .A1(n_600), .A2(n_666), .B(n_667), .Y(n_665) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g612 ( .A1(n_604), .A2(n_613), .B1(n_616), .B2(n_617), .C(n_619), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_604), .B(n_638), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_604), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g720 ( .A(n_610), .Y(n_720) );
INVxp67_ASAP7_75t_L g643 ( .A(n_611), .Y(n_643) );
INVx1_ASAP7_75t_L g650 ( .A(n_613), .Y(n_650) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
AND2x2_ASAP7_75t_L g689 ( .A(n_614), .B(n_618), .Y(n_689) );
INVx1_ASAP7_75t_L g663 ( .A(n_618), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_618), .B(n_633), .Y(n_693) );
OAI32xp33_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_622), .A3(n_624), .B1(n_625), .B2(n_626), .Y(n_619) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_SL g632 ( .A(n_627), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_627), .B(n_659), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_627), .B(n_688), .Y(n_719) );
NAND2x1p5_ASAP7_75t_L g727 ( .A(n_627), .B(n_638), .Y(n_727) );
NAND5xp2_ASAP7_75t_L g628 ( .A(n_629), .B(n_651), .C(n_664), .D(n_676), .E(n_677), .Y(n_628) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_633), .B1(n_634), .B2(n_636), .C(n_640), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NAND2xp33_ASAP7_75t_SL g655 ( .A(n_635), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_638), .B(n_707), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_639), .A2(n_652), .B1(n_655), .B2(n_659), .Y(n_651) );
INVx2_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
OAI211xp5_ASAP7_75t_SL g646 ( .A1(n_642), .A2(n_647), .B(n_648), .C(n_649), .Y(n_646) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_SL g674 ( .A(n_654), .Y(n_674) );
INVx1_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_663), .B(n_712), .Y(n_722) );
OR2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AOI222xp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_680), .B1(n_682), .B2(n_686), .C1(n_689), .C2(n_690), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
OAI221xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_694), .B1(n_696), .B2(n_698), .C(n_700), .Y(n_692) );
INVx1_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
OAI21xp33_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_702), .B(n_705), .Y(n_700) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g712 ( .A(n_704), .Y(n_712) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
OAI221xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_711), .B1(n_713), .B2(n_715), .C(n_717), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
INVxp67_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
A2O1A1Ixp33_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_727), .B(n_728), .C(n_730), .Y(n_723) );
INVxp67_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
OAI21xp33_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_732), .B(n_733), .Y(n_730) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_736), .A2(n_740), .B1(n_741), .B2(n_742), .Y(n_739) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
endmodule