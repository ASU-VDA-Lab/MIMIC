module fake_jpeg_14445_n_530 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_530);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_530;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_54),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_55),
.Y(n_133)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_17),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_57),
.B(n_61),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_58),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_59),
.Y(n_146)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_32),
.B(n_15),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_62),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_64),
.Y(n_127)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_65),
.Y(n_157)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_44),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_67),
.A2(n_38),
.B1(n_29),
.B2(n_45),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_15),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_68),
.B(n_75),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_70),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g131 ( 
.A(n_71),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_49),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_80),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_81),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_50),
.Y(n_82)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_14),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_84),
.B(n_12),
.Y(n_160)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_38),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_92),
.Y(n_118)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_88),
.Y(n_138)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_24),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_93),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

BUFx8_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_97),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_50),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_96),
.Y(n_120)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_43),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_50),
.Y(n_105)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_101),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_38),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_25),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_104),
.A2(n_114),
.B1(n_149),
.B2(n_161),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_105),
.B(n_89),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_98),
.A2(n_43),
.B1(n_44),
.B2(n_36),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_110),
.A2(n_111),
.B1(n_124),
.B2(n_99),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_82),
.A2(n_44),
.B1(n_36),
.B2(n_47),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_67),
.A2(n_38),
.B1(n_42),
.B2(n_49),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_96),
.A2(n_77),
.B1(n_64),
.B2(n_73),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_53),
.B(n_31),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_128),
.B(n_136),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_66),
.A2(n_47),
.B1(n_40),
.B2(n_37),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_135),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_70),
.B(n_31),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_141),
.B(n_144),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_74),
.B(n_40),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_76),
.B(n_22),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_79),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_86),
.A2(n_22),
.B1(n_25),
.B2(n_37),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_101),
.B(n_47),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_159),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_59),
.A2(n_45),
.B1(n_39),
.B2(n_19),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_155),
.B(n_62),
.C(n_63),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_93),
.B(n_45),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_160),
.B(n_0),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_52),
.A2(n_33),
.B1(n_30),
.B2(n_39),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_162),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_102),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_163),
.B(n_176),
.Y(n_233)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_103),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_164),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_125),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_166),
.B(n_170),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_135),
.A2(n_104),
.B1(n_29),
.B2(n_39),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_167),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_110),
.A2(n_94),
.B1(n_95),
.B2(n_58),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_168),
.A2(n_173),
.B1(n_189),
.B2(n_210),
.Y(n_264)
);

BUFx12f_ASAP7_75t_L g169 ( 
.A(n_116),
.Y(n_169)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_169),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_112),
.B(n_88),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_171),
.B(n_183),
.Y(n_226)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_172),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_124),
.A2(n_71),
.B1(n_69),
.B2(n_54),
.Y(n_173)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_174),
.Y(n_239)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_121),
.Y(n_175)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_175),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_177),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_178),
.Y(n_238)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_179),
.Y(n_242)
);

AND2x2_ASAP7_75t_SL g180 ( 
.A(n_115),
.B(n_97),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_180),
.B(n_200),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_113),
.A2(n_65),
.B1(n_90),
.B2(n_72),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_L g235 ( 
.A1(n_181),
.A2(n_190),
.B1(n_201),
.B2(n_220),
.Y(n_235)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_117),
.Y(n_182)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_182),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_107),
.B(n_91),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_131),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_184),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_33),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_186),
.B(n_209),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_123),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_187),
.B(n_192),
.Y(n_248)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_188),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_111),
.A2(n_81),
.B1(n_80),
.B2(n_83),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_132),
.A2(n_30),
.B1(n_26),
.B2(n_27),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_129),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_126),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_193),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_106),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_194),
.Y(n_240)
);

AOI32xp33_ASAP7_75t_L g195 ( 
.A1(n_142),
.A2(n_55),
.A3(n_51),
.B1(n_81),
.B2(n_80),
.Y(n_195)
);

AOI31xp33_ASAP7_75t_L g256 ( 
.A1(n_195),
.A2(n_156),
.A3(n_126),
.B(n_9),
.Y(n_256)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_196),
.Y(n_246)
);

AO21x1_ASAP7_75t_L g257 ( 
.A1(n_197),
.A2(n_213),
.B(n_215),
.Y(n_257)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_148),
.Y(n_199)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_199),
.Y(n_266)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_145),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_108),
.A2(n_27),
.B1(n_26),
.B2(n_19),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_121),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_202),
.B(n_203),
.Y(n_262)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_145),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_131),
.A2(n_19),
.B1(n_55),
.B2(n_51),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_204),
.A2(n_140),
.B1(n_189),
.B2(n_206),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_205),
.B(n_106),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_123),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_206),
.B(n_207),
.Y(n_253)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_122),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_208),
.A2(n_133),
.B(n_116),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_155),
.B(n_0),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_L g210 ( 
.A1(n_152),
.A2(n_63),
.B1(n_1),
.B2(n_2),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_118),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_211),
.B(n_214),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_152),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_212),
.A2(n_140),
.B1(n_134),
.B2(n_151),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_119),
.A2(n_13),
.B1(n_12),
.B2(n_5),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_130),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_122),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_216),
.B(n_217),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_129),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_143),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_218),
.B(n_219),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_120),
.B(n_5),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_171),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_221),
.B(n_224),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_185),
.A2(n_130),
.B1(n_137),
.B2(n_109),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_223),
.A2(n_225),
.B1(n_227),
.B2(n_234),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_170),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_185),
.A2(n_137),
.B1(n_109),
.B2(n_157),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_209),
.A2(n_157),
.B1(n_108),
.B2(n_127),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_198),
.A2(n_127),
.B1(n_143),
.B2(n_150),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_220),
.A2(n_150),
.B1(n_134),
.B2(n_151),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_237),
.A2(n_241),
.B1(n_267),
.B2(n_212),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_208),
.A2(n_183),
.B1(n_176),
.B2(n_166),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_247),
.A2(n_268),
.B1(n_252),
.B2(n_264),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_249),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_180),
.B(n_146),
.C(n_133),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_250),
.B(n_265),
.C(n_196),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_251),
.B(n_252),
.Y(n_313)
);

A2O1A1Ixp33_ASAP7_75t_SL g310 ( 
.A1(n_256),
.A2(n_261),
.B(n_271),
.C(n_257),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_186),
.A2(n_156),
.B(n_126),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_259),
.A2(n_271),
.B(n_193),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_180),
.B(n_7),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_261),
.Y(n_274)
);

NAND2xp33_ASAP7_75t_L g261 ( 
.A(n_191),
.B(n_156),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_211),
.B(n_8),
.C(n_9),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_188),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_205),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_268),
.B(n_229),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_205),
.A2(n_8),
.B(n_10),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_222),
.A2(n_182),
.B(n_162),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_273),
.A2(n_276),
.B(n_291),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_222),
.A2(n_202),
.B(n_179),
.Y(n_276)
);

NAND2xp33_ASAP7_75t_SL g361 ( 
.A(n_277),
.B(n_304),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_263),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_278),
.B(n_306),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_262),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_279),
.B(n_283),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_224),
.B(n_164),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_280),
.B(n_286),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_281),
.B(n_282),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_262),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_284),
.B(n_255),
.Y(n_337)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_243),
.Y(n_285)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_285),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_226),
.B(n_172),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_226),
.B(n_199),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_287),
.B(n_296),
.Y(n_354)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_243),
.Y(n_288)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_288),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_233),
.B(n_165),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_289),
.B(n_292),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_257),
.A2(n_210),
.B1(n_178),
.B2(n_203),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_290),
.Y(n_339)
);

AOI22x1_ASAP7_75t_L g291 ( 
.A1(n_225),
.A2(n_218),
.B1(n_200),
.B2(n_175),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_254),
.B(n_194),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_231),
.Y(n_294)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_294),
.Y(n_360)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_231),
.Y(n_295)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_295),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_221),
.B(n_11),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_11),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_298),
.B(n_301),
.Y(n_326)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_245),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_299),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_223),
.A2(n_174),
.B1(n_177),
.B2(n_169),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_300),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_270),
.B(n_169),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_258),
.Y(n_302)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_302),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_257),
.A2(n_169),
.B1(n_264),
.B2(n_236),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_303),
.B(n_230),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_228),
.A2(n_241),
.B(n_251),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_245),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_307),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_262),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_246),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_246),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_308),
.B(n_309),
.Y(n_334)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_242),
.Y(n_309)
);

OR2x2_ASAP7_75t_SL g321 ( 
.A(n_310),
.B(n_293),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_235),
.A2(n_227),
.B1(n_228),
.B2(n_236),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_311),
.A2(n_316),
.B1(n_240),
.B2(n_238),
.Y(n_340)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_242),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_312),
.B(n_318),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_269),
.B(n_265),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_314),
.B(n_319),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_229),
.A2(n_250),
.B(n_260),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_315),
.B(n_266),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_234),
.A2(n_237),
.B1(n_229),
.B2(n_259),
.Y(n_316)
);

BUFx24_ASAP7_75t_L g317 ( 
.A(n_244),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_317),
.Y(n_333)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_232),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_248),
.B(n_253),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_320),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_321),
.A2(n_331),
.B(n_316),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_313),
.A2(n_256),
.B(n_244),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_323),
.A2(n_325),
.B(n_273),
.Y(n_364)
);

AND2x6_ASAP7_75t_L g324 ( 
.A(n_304),
.B(n_258),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_324),
.B(n_353),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_313),
.A2(n_244),
.B(n_240),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_232),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_327),
.B(n_329),
.C(n_337),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_266),
.C(n_255),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_277),
.Y(n_336)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_336),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_340),
.A2(n_291),
.B1(n_317),
.B2(n_310),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_297),
.B(n_238),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_341),
.B(n_357),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_298),
.B(n_230),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_346),
.B(n_350),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_349),
.A2(n_275),
.B1(n_311),
.B2(n_281),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_280),
.B(n_230),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_296),
.B(n_239),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_301),
.Y(n_356)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_356),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_284),
.B(n_239),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_285),
.B(n_272),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_358),
.B(n_333),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_286),
.B(n_272),
.C(n_287),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_359),
.B(n_299),
.C(n_305),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_364),
.A2(n_368),
.B(n_396),
.Y(n_418)
);

OAI21xp33_ASAP7_75t_L g367 ( 
.A1(n_326),
.A2(n_274),
.B(n_279),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_367),
.A2(n_374),
.B1(n_394),
.B2(n_352),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_361),
.A2(n_293),
.B(n_276),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_369),
.A2(n_388),
.B(n_323),
.Y(n_419)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_370),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_361),
.A2(n_274),
.B(n_295),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_371),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_342),
.A2(n_294),
.B(n_288),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_372),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_354),
.B(n_308),
.Y(n_375)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_375),
.Y(n_402)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_328),
.Y(n_376)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_376),
.Y(n_404)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_328),
.Y(n_377)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_377),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_337),
.B(n_307),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_378),
.B(n_380),
.C(n_383),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_339),
.A2(n_355),
.B1(n_275),
.B2(n_349),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_379),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_354),
.B(n_318),
.Y(n_381)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_381),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_347),
.B(n_309),
.Y(n_382)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_382),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_357),
.B(n_310),
.C(n_312),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_339),
.A2(n_310),
.B1(n_291),
.B2(n_302),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_395),
.Y(n_398)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_334),
.Y(n_386)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_386),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_387),
.A2(n_390),
.B1(n_393),
.B2(n_373),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_342),
.A2(n_310),
.B(n_317),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_327),
.B(n_317),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_389),
.B(n_392),
.C(n_344),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_332),
.A2(n_340),
.B1(n_335),
.B2(n_347),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_341),
.B(n_331),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_332),
.A2(n_359),
.B1(n_345),
.B2(n_329),
.Y(n_393)
);

OAI21xp33_ASAP7_75t_L g394 ( 
.A1(n_326),
.A2(n_321),
.B(n_332),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_334),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_322),
.A2(n_331),
.B(n_325),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_350),
.B(n_353),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_397),
.B(n_338),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_380),
.B(n_352),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_400),
.B(n_406),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_376),
.B(n_330),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_409),
.A2(n_412),
.B(n_419),
.Y(n_439)
);

AND2x6_ASAP7_75t_L g412 ( 
.A(n_365),
.B(n_324),
.Y(n_412)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_413),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_397),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_414),
.B(n_423),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_375),
.B(n_338),
.Y(n_415)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_415),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_391),
.B(n_330),
.Y(n_416)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_416),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_366),
.B(n_322),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_417),
.B(n_422),
.Y(n_433)
);

AO21x2_ASAP7_75t_L g420 ( 
.A1(n_372),
.A2(n_345),
.B(n_344),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_420),
.B(n_387),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_377),
.B(n_346),
.Y(n_421)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_421),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_382),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_386),
.B(n_343),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_424),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_366),
.B(n_348),
.C(n_360),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_426),
.B(n_383),
.C(n_385),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_427),
.A2(n_395),
.B1(n_365),
.B2(n_390),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_413),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_428),
.B(n_445),
.Y(n_456)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_399),
.Y(n_429)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_429),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_430),
.B(n_431),
.C(n_434),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_426),
.B(n_378),
.C(n_389),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_432),
.A2(n_405),
.B(n_420),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_408),
.B(n_385),
.C(n_392),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_408),
.B(n_393),
.C(n_371),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_435),
.B(n_451),
.C(n_452),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_415),
.B(n_381),
.Y(n_437)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_437),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_440),
.A2(n_420),
.B1(n_399),
.B2(n_404),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_417),
.B(n_396),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_441),
.B(n_449),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_422),
.B(n_368),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_442),
.B(n_427),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_398),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_409),
.B(n_364),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_404),
.Y(n_450)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_450),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_418),
.B(n_388),
.C(n_370),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_418),
.B(n_369),
.C(n_358),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_410),
.A2(n_363),
.B(n_343),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_453),
.A2(n_410),
.B(n_403),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_454),
.A2(n_473),
.B(n_453),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_443),
.A2(n_425),
.B1(n_398),
.B2(n_407),
.Y(n_455)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_455),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_446),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_457),
.B(n_465),
.Y(n_475)
);

BUFx24_ASAP7_75t_SL g458 ( 
.A(n_447),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_458),
.B(n_433),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_440),
.A2(n_448),
.B1(n_436),
.B2(n_438),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_461),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g484 ( 
.A(n_463),
.B(n_467),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_452),
.A2(n_403),
.B1(n_401),
.B2(n_402),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_464),
.B(n_469),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_444),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_431),
.B(n_419),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_433),
.B(n_401),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_471),
.B(n_472),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_441),
.B(n_405),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_435),
.B(n_402),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_474),
.B(n_470),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_476),
.B(n_483),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_454),
.A2(n_451),
.B(n_439),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_477),
.A2(n_481),
.B(n_467),
.Y(n_494)
);

NOR2xp67_ASAP7_75t_L g481 ( 
.A(n_470),
.B(n_442),
.Y(n_481)
);

AO22x2_ASAP7_75t_L g482 ( 
.A1(n_473),
.A2(n_432),
.B1(n_407),
.B2(n_411),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_482),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_471),
.B(n_430),
.C(n_434),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_485),
.B(n_486),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_456),
.B(n_439),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_488),
.B(n_489),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_468),
.B(n_449),
.C(n_429),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_468),
.B(n_437),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_490),
.B(n_420),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_489),
.B(n_463),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_491),
.B(n_496),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_494),
.A2(n_495),
.B(n_486),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_477),
.A2(n_464),
.B(n_466),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_479),
.B(n_466),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_484),
.B(n_469),
.C(n_459),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_497),
.B(n_498),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_484),
.B(n_460),
.C(n_411),
.Y(n_498)
);

OAI321xp33_ASAP7_75t_L g499 ( 
.A1(n_478),
.A2(n_462),
.A3(n_412),
.B1(n_420),
.B2(n_362),
.C(n_360),
.Y(n_499)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_499),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_475),
.B(n_348),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_501),
.B(n_351),
.Y(n_506)
);

AOI31xp67_ASAP7_75t_SL g513 ( 
.A1(n_502),
.A2(n_503),
.A3(n_482),
.B(n_487),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_480),
.B(n_362),
.Y(n_503)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_505),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_506),
.B(n_507),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_500),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_492),
.B(n_485),
.C(n_487),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_511),
.B(n_512),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_493),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_513),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_496),
.B(n_351),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_514),
.B(n_498),
.Y(n_515)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_515),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_508),
.B(n_491),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_516),
.B(n_497),
.Y(n_522)
);

NAND3xp33_ASAP7_75t_L g521 ( 
.A(n_519),
.B(n_509),
.C(n_510),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_521),
.A2(n_524),
.B(n_520),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_522),
.B(n_517),
.C(n_518),
.Y(n_525)
);

AOI21xp33_ASAP7_75t_L g524 ( 
.A1(n_518),
.A2(n_506),
.B(n_504),
.Y(n_524)
);

CKINVDCx16_ASAP7_75t_R g527 ( 
.A(n_525),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_526),
.B(n_523),
.C(n_482),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_528),
.A2(n_482),
.B(n_351),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_529),
.B(n_527),
.Y(n_530)
);


endmodule