module real_jpeg_3789_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_1),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_1),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_1),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_1),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_1),
.B(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_1),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_1),
.B(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_1),
.B(n_353),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_2),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_2),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_2),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_2),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_2),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_2),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_2),
.B(n_374),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_3),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_4),
.B(n_133),
.Y(n_227)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_4),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_4),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_4),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_4),
.B(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_4),
.B(n_390),
.Y(n_389)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_6),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_6),
.Y(n_209)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_6),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_6),
.Y(n_374)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_7),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_7),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_7),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_7),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_8),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_8),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_8),
.B(n_49),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_8),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_8),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_8),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_8),
.B(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_8),
.Y(n_179)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_10),
.Y(n_91)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_10),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_10),
.Y(n_158)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_10),
.Y(n_178)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_10),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_11),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_11),
.B(n_110),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_11),
.B(n_147),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_11),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_11),
.B(n_49),
.Y(n_167)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_12),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_12),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_12),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_12),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_12),
.B(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_12),
.Y(n_245)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_13),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_14),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_14),
.B(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_14),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_14),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_14),
.B(n_407),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_15),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_15),
.B(n_49),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_15),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_15),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_15),
.B(n_133),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_15),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_15),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_192),
.B1(n_448),
.B2(n_449),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g448 ( 
.A(n_18),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_191),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_160),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_21),
.B(n_160),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_98),
.C(n_135),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_22),
.B(n_335),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_68),
.C(n_79),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_23),
.B(n_330),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_41),
.C(n_57),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_24),
.B(n_289),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_35),
.B2(n_36),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_31),
.B2(n_34),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_27),
.A2(n_28),
.B1(n_105),
.B2(n_106),
.Y(n_306)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_28),
.B(n_31),
.C(n_36),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_28),
.B(n_106),
.C(n_215),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_29),
.Y(n_346)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_30),
.Y(n_111)
);

BUFx8_ASAP7_75t_L g408 ( 
.A(n_30),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_31),
.A2(n_34),
.B1(n_109),
.B2(n_112),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_31),
.B(n_109),
.C(n_146),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_31),
.A2(n_34),
.B1(n_359),
.B2(n_360),
.Y(n_377)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

OR2x2_ASAP7_75t_SL g59 ( 
.A(n_32),
.B(n_60),
.Y(n_59)
);

OR2x2_ASAP7_75t_SL g86 ( 
.A(n_32),
.B(n_87),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_32),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_34),
.B(n_359),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_35),
.A2(n_36),
.B1(n_182),
.B2(n_186),
.Y(n_181)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_38),
.Y(n_129)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_39),
.Y(n_257)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_41),
.B(n_57),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_48),
.C(n_53),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_42),
.B(n_283),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g185 ( 
.A(n_47),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_47),
.Y(n_213)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_47),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_48),
.A2(n_128),
.B1(n_130),
.B2(n_131),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_48),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_48),
.B(n_53),
.Y(n_283)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_52),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_52),
.Y(n_219)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_56),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_62),
.B2(n_67),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_77),
.C(n_78),
.Y(n_76)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_64),
.Y(n_78)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_66),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_68),
.B(n_79),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_76),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_69)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_72),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_72),
.B(n_74),
.C(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_72),
.A2(n_75),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_75),
.B(n_154),
.C(n_157),
.Y(n_175)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_76),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_92),
.C(n_95),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_81),
.B(n_295),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.C(n_90),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_82),
.A2(n_90),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_82),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_82),
.A2(n_233),
.B1(n_265),
.B2(n_266),
.Y(n_368)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_86),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_86),
.Y(n_229)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_87),
.Y(n_314)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_89),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_90),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_92),
.B(n_95),
.Y(n_295)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_98),
.B(n_135),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_113),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_99),
.B(n_114),
.C(n_125),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_100),
.B(n_106),
.C(n_109),
.Y(n_171)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_109),
.B2(n_112),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_105),
.A2(n_106),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_109),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_109),
.B(n_308),
.C(n_312),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_109),
.A2(n_112),
.B1(n_355),
.B2(n_356),
.Y(n_354)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_125),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_119),
.C(n_121),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_115),
.A2(n_140),
.B1(n_255),
.B2(n_258),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_115),
.B(n_167),
.C(n_255),
.Y(n_281)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_119),
.B(n_121),
.Y(n_141)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx5_ASAP7_75t_L g350 ( 
.A(n_124),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_124),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_124),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_132),
.B2(n_134),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_131),
.C(n_132),
.Y(n_172)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_129),
.Y(n_273)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_132),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_150),
.B2(n_159),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_151),
.C(n_153),
.Y(n_161)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_143),
.C(n_144),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_138),
.A2(n_139),
.B1(n_143),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_143),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_144),
.B(n_327),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_148),
.B2(n_149),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_153),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx24_ASAP7_75t_SL g451 ( 
.A(n_160),
.Y(n_451)
);

FAx1_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_162),
.CI(n_173),
.CON(n_160),
.SN(n_160)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_169),
.B2(n_170),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_167),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_167),
.A2(n_168),
.B1(n_254),
.B2(n_259),
.Y(n_253)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_173)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_180),
.B1(n_181),
.B2(n_187),
.Y(n_176)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_177),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_182),
.Y(n_186)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_188),
.Y(n_190)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_192),
.Y(n_449)
);

AO21x2_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_333),
.B(n_336),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_322),
.B(n_332),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_298),
.B(n_321),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_195),
.B(n_446),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_285),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_196),
.B(n_285),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_252),
.C(n_279),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_197),
.B(n_320),
.Y(n_319)
);

BUFx24_ASAP7_75t_SL g450 ( 
.A(n_197),
.Y(n_450)
);

FAx1_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_228),
.CI(n_234),
.CON(n_197),
.SN(n_197)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_198),
.B(n_228),
.C(n_234),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_214),
.C(n_220),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_199),
.B(n_317),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_210),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_206),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_201),
.B(n_206),
.C(n_210),
.Y(n_284)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_202),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_204),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_205),
.Y(n_383)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_213),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_214),
.A2(n_220),
.B1(n_221),
.B2(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_214),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_215),
.B(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_226),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_222),
.A2(n_223),
.B1(n_226),
.B2(n_227),
.Y(n_315)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_225),
.Y(n_400)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_265),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_243),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_235),
.A2(n_236),
.B(n_238),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_235),
.B(n_244),
.C(n_247),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_242),
.Y(n_238)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_242),
.B(n_383),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_247),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_248),
.B(n_352),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_248),
.B(n_365),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_248),
.B(n_398),
.Y(n_397)
);

INVx8_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_252),
.B(n_279),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_260),
.C(n_262),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_253),
.A2(n_260),
.B1(n_261),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_253),
.Y(n_303)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_254),
.Y(n_259)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_255),
.Y(n_258)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_262),
.B(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_270),
.C(n_274),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_263),
.A2(n_264),
.B1(n_435),
.B2(n_436),
.Y(n_434)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_270),
.A2(n_271),
.B1(n_274),
.B2(n_275),
.Y(n_436)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_284),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_282),
.C(n_284),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_286),
.B(n_288),
.C(n_297),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_290),
.B1(n_296),
.B2(n_297),
.Y(n_287)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_288),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_290),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_291),
.B(n_293),
.C(n_294),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_319),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_299),
.B(n_319),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_304),
.C(n_316),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_300),
.A2(n_301),
.B1(n_441),
.B2(n_442),
.Y(n_440)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_304),
.B(n_316),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_307),
.C(n_315),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_305),
.B(n_428),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_307),
.B(n_315),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_308),
.A2(n_309),
.B1(n_312),
.B2(n_313),
.Y(n_356)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_311),
.Y(n_353)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_323),
.B(n_333),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_325),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_334),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g447 ( 
.A(n_325),
.B(n_334),
.Y(n_447)
);

FAx1_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_329),
.CI(n_331),
.CON(n_325),
.SN(n_325)
);

OAI31xp33_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_444),
.A3(n_445),
.B(n_447),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_438),
.B(n_443),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_339),
.A2(n_423),
.B(n_437),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_378),
.B(n_422),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_341),
.B(n_369),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_341),
.B(n_369),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_357),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_354),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_343),
.B(n_354),
.C(n_357),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_347),
.C(n_351),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_344),
.A2(n_345),
.B1(n_347),
.B2(n_348),
.Y(n_371)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_351),
.B(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_358),
.B(n_363),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_358),
.B(n_432),
.C(n_433),
.Y(n_431)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_368),
.Y(n_363)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_364),
.Y(n_432)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_368),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_372),
.C(n_377),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_370),
.B(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_372),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_372),
.A2(n_377),
.B1(n_414),
.B2(n_420),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_373),
.B(n_375),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_373),
.Y(n_412)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_374),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_375),
.Y(n_413)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_377),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_379),
.A2(n_416),
.B(n_421),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_380),
.A2(n_402),
.B(n_415),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_387),
.B(n_401),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_384),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_386),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_388),
.B(n_397),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_388),
.B(n_397),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_389),
.A2(n_392),
.B(n_396),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_389),
.B(n_392),
.Y(n_396)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_396),
.A2(n_404),
.B1(n_409),
.B2(n_410),
.Y(n_403)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_396),
.Y(n_409)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx8_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_403),
.B(n_411),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_403),
.B(n_411),
.Y(n_415)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_404),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_405),
.B(n_406),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_405),
.A2(n_406),
.B(n_409),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_412),
.A2(n_413),
.B(n_414),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_417),
.B(n_418),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_425),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_424),
.B(n_425),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_426),
.A2(n_427),
.B1(n_429),
.B2(n_430),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_426),
.B(n_431),
.C(n_434),
.Y(n_439)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_434),
.Y(n_430)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_440),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_439),
.B(n_440),
.Y(n_443)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_441),
.Y(n_442)
);


endmodule