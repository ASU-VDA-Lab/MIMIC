module fake_jpeg_13789_n_190 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_190);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_190;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_4),
.B(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_11),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_46),
.Y(n_58)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_24),
.B(n_19),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_45),
.B(n_50),
.Y(n_57)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_49),
.Y(n_60)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

NOR2x1_ASAP7_75t_R g76 ( 
.A(n_48),
.B(n_30),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_21),
.B(n_10),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_52),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_22),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_21),
.B(n_10),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_54),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_24),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_62),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_48),
.A2(n_28),
.B1(n_16),
.B2(n_31),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_59),
.A2(n_7),
.B(n_65),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_31),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_16),
.B1(n_29),
.B2(n_23),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_63),
.A2(n_75),
.B1(n_1),
.B2(n_6),
.Y(n_95)
);

AOI21xp33_ASAP7_75t_L g66 ( 
.A1(n_35),
.A2(n_33),
.B(n_25),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_51),
.C(n_34),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_37),
.A2(n_33),
.B1(n_25),
.B2(n_20),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_67),
.A2(n_78),
.B1(n_81),
.B2(n_7),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_20),
.B1(n_17),
.B2(n_26),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_73),
.B1(n_82),
.B2(n_59),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_36),
.A2(n_17),
.B1(n_27),
.B2(n_26),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_27),
.B1(n_30),
.B2(n_2),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_38),
.A2(n_30),
.B1(n_1),
.B2(n_2),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_42),
.B(n_0),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_80),
.B(n_55),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_47),
.A2(n_30),
.B1(n_3),
.B2(n_5),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_39),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_85),
.Y(n_118)
);

BUFx2_ASAP7_75t_SL g87 ( 
.A(n_56),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_88),
.B(n_90),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_58),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_92),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_64),
.B(n_9),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_51),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

BUFx12_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_97),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_99),
.B1(n_102),
.B2(n_107),
.Y(n_120)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_6),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_66),
.A2(n_62),
.B1(n_57),
.B2(n_80),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_61),
.B1(n_83),
.B2(n_92),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_57),
.B(n_70),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_72),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_70),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_61),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

INVx3_ASAP7_75t_SL g106 ( 
.A(n_77),
.Y(n_106)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_77),
.A2(n_72),
.B1(n_81),
.B2(n_78),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_119),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_74),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_124),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_85),
.A2(n_61),
.B1(n_74),
.B2(n_102),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_118),
.B1(n_120),
.B2(n_109),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_117),
.B(n_125),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_103),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_89),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_127),
.Y(n_129)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_101),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_132),
.B(n_134),
.Y(n_154)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_133),
.B(n_137),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_116),
.B(n_83),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_91),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_139),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_98),
.C(n_96),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_138),
.A2(n_113),
.B1(n_118),
.B2(n_115),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_100),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_84),
.C(n_106),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_141),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_105),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_123),
.Y(n_145)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_146),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_140),
.A2(n_116),
.B1(n_123),
.B2(n_111),
.Y(n_151)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_138),
.A2(n_106),
.B1(n_122),
.B2(n_108),
.Y(n_153)
);

AO221x1_ASAP7_75t_L g164 ( 
.A1(n_153),
.A2(n_136),
.B1(n_129),
.B2(n_133),
.C(n_143),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_108),
.B(n_114),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_142),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_130),
.A2(n_94),
.B1(n_126),
.B2(n_128),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_156),
.B(n_157),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_128),
.A2(n_94),
.B1(n_126),
.B2(n_130),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_157),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_158),
.B(n_165),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_154),
.B(n_134),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_166),
.Y(n_168)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

BUFx24_ASAP7_75t_SL g166 ( 
.A(n_154),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_149),
.B(n_137),
.Y(n_167)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_156),
.Y(n_171)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_171),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_161),
.A2(n_151),
.B(n_155),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_172),
.A2(n_161),
.B(n_163),
.Y(n_175)
);

AO21x1_ASAP7_75t_L g182 ( 
.A1(n_175),
.A2(n_171),
.B(n_173),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_160),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_176),
.B(n_179),
.Y(n_181)
);

OAI322xp33_ASAP7_75t_L g177 ( 
.A1(n_168),
.A2(n_150),
.A3(n_147),
.B1(n_160),
.B2(n_165),
.C1(n_146),
.C2(n_148),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_147),
.Y(n_180)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_182),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_172),
.C(n_170),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_183),
.A2(n_178),
.B1(n_152),
.B2(n_144),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_152),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_184),
.B(n_181),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_186),
.B(n_187),
.C(n_182),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_185),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_94),
.Y(n_190)
);


endmodule