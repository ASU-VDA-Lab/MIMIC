module real_jpeg_2188_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_273, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_273;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_173;
wire n_243;
wire n_105;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_18;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_187;
wire n_75;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_213;
wire n_167;
wire n_202;
wire n_179;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_89;

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_2),
.A2(n_37),
.B1(n_59),
.B2(n_60),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_2),
.A2(n_37),
.B1(n_70),
.B2(n_71),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_2),
.A2(n_37),
.B1(n_43),
.B2(n_44),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_3),
.A2(n_70),
.B1(n_71),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_3),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_3),
.A2(n_59),
.B1(n_60),
.B2(n_77),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_77),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_3),
.A2(n_43),
.B1(n_44),
.B2(n_77),
.Y(n_213)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_5),
.A2(n_70),
.B1(n_71),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_5),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_156),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_156),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_5),
.A2(n_59),
.B1(n_60),
.B2(n_156),
.Y(n_216)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_6),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_7),
.A2(n_33),
.B1(n_70),
.B2(n_71),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_7),
.A2(n_33),
.B1(n_43),
.B2(n_44),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_7),
.A2(n_33),
.B1(n_59),
.B2(n_60),
.Y(n_128)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_10),
.A2(n_43),
.B1(n_44),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_10),
.A2(n_52),
.B1(n_59),
.B2(n_60),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_52),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_11),
.A2(n_43),
.B1(n_44),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_11),
.A2(n_50),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_50),
.Y(n_149)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_12),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_13),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_13),
.B(n_32),
.C(n_46),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_145),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_13),
.B(n_29),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_13),
.B(n_97),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_13),
.B(n_59),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_13),
.A2(n_59),
.B(n_207),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_13),
.B(n_79),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_13),
.A2(n_70),
.B(n_243),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_14),
.A2(n_70),
.B1(n_71),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_14),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_14),
.A2(n_43),
.B1(n_44),
.B2(n_126),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_126),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_14),
.A2(n_59),
.B1(n_60),
.B2(n_126),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_132),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_130),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_109),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_20),
.B(n_109),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_81),
.B2(n_82),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_53),
.C(n_67),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_23),
.A2(n_24),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_39),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_25),
.A2(n_26),
.B1(n_39),
.B2(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_34),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_27),
.A2(n_38),
.B(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_32),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_28),
.A2(n_30),
.B(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_28),
.A2(n_87),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_28),
.A2(n_35),
.B(n_149),
.Y(n_233)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_29),
.B(n_36),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_29),
.A2(n_38),
.B1(n_121),
.B2(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_29),
.A2(n_38),
.B1(n_145),
.B2(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_29),
.A2(n_38),
.B1(n_187),
.B2(n_190),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_30),
.A2(n_87),
.B(n_122),
.Y(n_209)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_31),
.A2(n_32),
.B1(n_46),
.B2(n_47),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_32),
.B(n_185),
.Y(n_184)
);

INVxp33_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_38),
.Y(n_87)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_39),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_40),
.A2(n_51),
.B(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_40),
.A2(n_48),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_40),
.A2(n_95),
.B(n_101),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_41),
.B(n_96),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_41),
.A2(n_97),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_41),
.A2(n_97),
.B1(n_172),
.B2(n_180),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_41),
.A2(n_100),
.B(n_222),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_48),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_42)
);

OA22x2_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_44),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_43),
.B(n_55),
.Y(n_208)
);

CKINVDCx6p67_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_44),
.B(n_177),
.Y(n_176)
);

OAI32xp33_ASAP7_75t_L g205 ( 
.A1(n_44),
.A2(n_56),
.A3(n_59),
.B1(n_206),
.B2(n_208),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_48),
.B(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_48),
.A2(n_49),
.B(n_103),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_53),
.B(n_67),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_58),
.B(n_62),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_54),
.B(n_145),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_54),
.A2(n_65),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_54),
.A2(n_65),
.B1(n_151),
.B2(n_228),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_66)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_60),
.B1(n_73),
.B2(n_74),
.Y(n_75)
);

NAND3xp33_ASAP7_75t_L g146 ( 
.A(n_59),
.B(n_71),
.C(n_74),
.Y(n_146)
);

CKINVDCx6p67_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_60),
.A2(n_73),
.B(n_144),
.C(n_146),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_63),
.B(n_106),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_64),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_64),
.A2(n_106),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_65),
.A2(n_128),
.B(n_129),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_65),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_76),
.B(n_78),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_68),
.A2(n_90),
.B(n_91),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_68),
.A2(n_75),
.B1(n_76),
.B2(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_68),
.A2(n_75),
.B1(n_125),
.B2(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_68),
.A2(n_75),
.B1(n_155),
.B2(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_75),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_71),
.B(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_73),
.Y(n_74)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_92),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_80),
.Y(n_90)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_98),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_93),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_88),
.B2(n_89),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_85),
.A2(n_86),
.B1(n_94),
.B2(n_114),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_87),
.A2(n_120),
.B(n_122),
.Y(n_119)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_94),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_104),
.B(n_108),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_104),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_102),
.Y(n_99)
);

INVxp33_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_106),
.B(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.C(n_115),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_110),
.B(n_113),
.Y(n_159)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_115),
.A2(n_116),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_124),
.C(n_127),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_118),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_119),
.B(n_123),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_127),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_160),
.B(n_270),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_157),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_134),
.B(n_157),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.C(n_140),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_135),
.B(n_138),
.Y(n_255)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_140),
.B(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_150),
.C(n_154),
.Y(n_140)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_141),
.B(n_150),
.CI(n_154),
.CON(n_258),
.SN(n_258)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_147),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_142),
.A2(n_143),
.B1(n_147),
.B2(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_144),
.Y(n_243)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_147),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

AOI321xp33_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_253),
.A3(n_262),
.B1(n_268),
.B2(n_269),
.C(n_273),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_236),
.B(n_252),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_218),
.B(n_235),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_200),
.B(n_217),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_181),
.B(n_199),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_174),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_174),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_171),
.C(n_202),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_168),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_173),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_175),
.A2(n_176),
.B1(n_178),
.B2(n_179),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_193),
.B(n_198),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_188),
.B(n_192),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_191),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_190),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_197),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_203),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_203),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_210),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_211),
.C(n_214),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_209),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_209),
.Y(n_223)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_213),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_216),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_234),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_234),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_224),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_223),
.C(n_224),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_229),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_231),
.C(n_232),
.Y(n_249)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_238),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_247),
.B2(n_248),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_249),
.C(n_250),
.Y(n_263)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_244),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_245),
.C(n_246),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_256),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_259),
.C(n_261),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_257),
.A2(n_258),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx24_ASAP7_75t_SL g272 ( 
.A(n_258),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_259),
.A2(n_260),
.B1(n_261),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_261),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_264),
.Y(n_268)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);


endmodule