module fake_jpeg_4700_n_185 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_185);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_6),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_10),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_33),
.B(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g36 ( 
.A1(n_16),
.A2(n_1),
.B(n_2),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_36),
.B(n_39),
.Y(n_69)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_38),
.A2(n_46),
.B1(n_25),
.B2(n_8),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_2),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_20),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_41),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_20),
.B(n_3),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_23),
.B(n_3),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_29),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_51),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_29),
.B1(n_26),
.B2(n_21),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_52),
.A2(n_56),
.B1(n_67),
.B2(n_68),
.Y(n_99)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_55),
.B(n_58),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_26),
.B1(n_21),
.B2(n_24),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_31),
.A2(n_21),
.B1(n_26),
.B2(n_18),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_59),
.A2(n_63),
.B(n_64),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_62),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_33),
.A2(n_24),
.B1(n_27),
.B2(n_19),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_41),
.A2(n_24),
.B1(n_27),
.B2(n_19),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_15),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_65),
.B(n_66),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_15),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_41),
.A2(n_15),
.B1(n_27),
.B2(n_19),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_35),
.A2(n_14),
.B1(n_17),
.B2(n_28),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_14),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_70),
.B(n_71),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_35),
.B(n_17),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_28),
.Y(n_73)
);

FAx1_ASAP7_75t_SL g96 ( 
.A(n_73),
.B(n_16),
.CI(n_10),
.CON(n_96),
.SN(n_96)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_47),
.A2(n_25),
.B1(n_16),
.B2(n_9),
.Y(n_74)
);

BUFx4f_ASAP7_75t_SL g102 ( 
.A(n_74),
.Y(n_102)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_75),
.B(n_77),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_76),
.A2(n_75),
.B1(n_57),
.B2(n_55),
.Y(n_101)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_41),
.B(n_25),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_7),
.Y(n_90)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_79),
.Y(n_83)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_78),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_82),
.B(n_87),
.Y(n_128)
);

AND2x6_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_22),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_90),
.B(n_96),
.Y(n_107)
);

AND2x6_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_22),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_92),
.B(n_94),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_7),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_69),
.A2(n_16),
.B(n_22),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_61),
.B(n_81),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_57),
.B(n_9),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_103),
.B(n_104),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_12),
.Y(n_104)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_54),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_73),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_108),
.B(n_109),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_72),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_102),
.A2(n_80),
.B1(n_79),
.B2(n_49),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_83),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_114),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_72),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_88),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_92),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_117),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_50),
.Y(n_116)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_51),
.Y(n_120)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_60),
.B1(n_58),
.B2(n_77),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_94),
.B(n_48),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_81),
.B1(n_54),
.B2(n_12),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_99),
.A2(n_81),
.B1(n_11),
.B2(n_10),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_127),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_125),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_140),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_82),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_142),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_97),
.B1(n_102),
.B2(n_95),
.Y(n_135)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_112),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_119),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_85),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_85),
.Y(n_141)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_81),
.C(n_91),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_123),
.A2(n_91),
.B1(n_100),
.B2(n_93),
.Y(n_143)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_142),
.A2(n_118),
.B(n_136),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_147),
.A2(n_148),
.B(n_156),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_140),
.A2(n_115),
.B(n_113),
.Y(n_148)
);

AOI221xp5_ASAP7_75t_L g150 ( 
.A1(n_135),
.A2(n_123),
.B1(n_124),
.B2(n_107),
.C(n_122),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_150),
.B(n_133),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_137),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_117),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_144),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_154),
.B(n_139),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_121),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_147),
.A2(n_132),
.B(n_138),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_157),
.A2(n_162),
.B(n_165),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_146),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_160),
.B(n_164),
.Y(n_172)
);

NAND3xp33_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_163),
.C(n_156),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_139),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_119),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_148),
.A2(n_149),
.B(n_156),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_145),
.C(n_155),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_169),
.C(n_171),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_170),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_165),
.A2(n_149),
.B1(n_153),
.B2(n_144),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_145),
.C(n_155),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_172),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_173),
.B(n_174),
.Y(n_178)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_157),
.C(n_158),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_177),
.A2(n_171),
.B1(n_152),
.B2(n_114),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_179),
.B(n_180),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_175),
.A2(n_110),
.B1(n_129),
.B2(n_143),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_178),
.A2(n_176),
.B1(n_154),
.B2(n_131),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_180),
.B1(n_127),
.B2(n_134),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_181),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_184),
.Y(n_185)
);


endmodule