module fake_jpeg_3024_n_143 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_143);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_0),
.B(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_30),
.A2(n_28),
.B1(n_16),
.B2(n_22),
.Y(n_52)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_40),
.Y(n_48)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_42),
.Y(n_62)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_SL g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

NAND2xp33_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_18),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_7),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_25),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_21),
.B1(n_27),
.B2(n_20),
.Y(n_45)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_43),
.B(n_18),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_45),
.B(n_51),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_22),
.C(n_19),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_29),
.C(n_3),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_21),
.B1(n_27),
.B2(n_28),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_50),
.A2(n_52),
.B1(n_57),
.B2(n_11),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_36),
.B(n_19),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_14),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_14),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_59),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_29),
.B(n_8),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_16),
.B1(n_29),
.B2(n_2),
.Y(n_57)
);

NOR2x1_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_38),
.B(n_5),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_5),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_74),
.Y(n_84)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

AO22x1_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_81),
.B1(n_57),
.B2(n_45),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_70),
.B(n_78),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_80),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_48),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_76),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_63),
.Y(n_76)
);

NAND2x1_ASAP7_75t_SL g77 ( 
.A(n_44),
.B(n_8),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_79),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_62),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_82),
.B(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_64),
.B(n_60),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_69),
.B(n_49),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_88),
.B(n_96),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_52),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_94),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_80),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_59),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_61),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_SL g96 ( 
.A(n_68),
.B(n_62),
.C(n_56),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_79),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_99),
.B(n_104),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

AO22x1_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_67),
.B1(n_72),
.B2(n_75),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_103),
.A2(n_109),
.B1(n_92),
.B2(n_84),
.Y(n_110)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

AOI21x1_ASAP7_75t_SL g105 ( 
.A1(n_94),
.A2(n_77),
.B(n_76),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_105),
.A2(n_87),
.B(n_90),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_107),
.Y(n_113)
);

OA21x2_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_61),
.B(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_110),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_107),
.A2(n_93),
.B1(n_82),
.B2(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_97),
.B(n_107),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

AO21x1_ASAP7_75t_L g126 ( 
.A1(n_117),
.A2(n_119),
.B(n_105),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_90),
.B(n_71),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_102),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_126),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_112),
.B(n_102),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_125),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_131),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_120),
.A2(n_115),
.B1(n_113),
.B2(n_103),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_SL g133 ( 
.A1(n_130),
.A2(n_113),
.B(n_114),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_121),
.C(n_106),
.Y(n_131)
);

AOI21xp33_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_121),
.B(n_128),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_132),
.A2(n_135),
.B(n_103),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_128),
.Y(n_136)
);

AO21x1_ASAP7_75t_L g135 ( 
.A1(n_131),
.A2(n_114),
.B(n_116),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_136),
.A2(n_12),
.B(n_47),
.Y(n_139)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_138),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_47),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_140),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_47),
.Y(n_143)
);


endmodule