module real_jpeg_14629_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_3),
.A2(n_69),
.B1(n_72),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_3),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_3),
.A2(n_60),
.B1(n_61),
.B2(n_113),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_113),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_113),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_6),
.A2(n_69),
.B1(n_72),
.B2(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_6),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_6),
.A2(n_60),
.B1(n_61),
.B2(n_79),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_6),
.A2(n_44),
.B1(n_45),
.B2(n_79),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_79),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_7),
.A2(n_38),
.B1(n_44),
.B2(n_45),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_7),
.A2(n_38),
.B1(n_60),
.B2(n_61),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_9),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_47),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_9),
.A2(n_47),
.B1(n_60),
.B2(n_61),
.Y(n_130)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_11),
.A2(n_72),
.B(n_75),
.C(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_11),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_11),
.A2(n_69),
.B1(n_72),
.B2(n_102),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_11),
.B(n_80),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_11),
.A2(n_44),
.B1(n_45),
.B2(n_102),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_11),
.A2(n_24),
.B1(n_36),
.B2(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_11),
.B(n_108),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_12),
.A2(n_68),
.B1(n_69),
.B2(n_72),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_12),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_12),
.A2(n_60),
.B1(n_61),
.B2(n_68),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_12),
.A2(n_44),
.B1(n_45),
.B2(n_68),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_68),
.Y(n_209)
);

BUFx8_ASAP7_75t_L g75 ( 
.A(n_13),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_14),
.A2(n_60),
.B1(n_61),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_14),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_63),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_14),
.A2(n_63),
.B1(n_69),
.B2(n_72),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_63),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_15),
.A2(n_33),
.B1(n_44),
.B2(n_45),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_141),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_140),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_115),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_20),
.B(n_115),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_81),
.C(n_93),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_21),
.B(n_81),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_53),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_22),
.B(n_54),
.C(n_66),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_23),
.B(n_39),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_31),
.B(n_34),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_24),
.A2(n_36),
.B(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_24),
.A2(n_36),
.B1(n_209),
.B2(n_217),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_24),
.A2(n_84),
.B(n_211),
.Y(n_226)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_25),
.B(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_25),
.A2(n_30),
.B1(n_32),
.B2(n_98),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_25),
.A2(n_35),
.B(n_85),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_25),
.A2(n_30),
.B1(n_208),
.B2(n_210),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g40 ( 
.A1(n_26),
.A2(n_27),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_26),
.B(n_41),
.C(n_102),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_26),
.B(n_215),
.Y(n_214)
);

CKINVDCx6p67_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_30),
.B(n_85),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_36),
.A2(n_86),
.B(n_99),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_36),
.B(n_102),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_43),
.B(n_48),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_40),
.B(n_50),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_40),
.B(n_102),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_52)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

OA22x2_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_45),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_SL g177 ( 
.A1(n_44),
.A2(n_57),
.B(n_178),
.C(n_180),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_44),
.B(n_201),
.Y(n_200)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

NOR3xp33_ASAP7_75t_L g180 ( 
.A(n_45),
.B(n_58),
.C(n_60),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_51),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_51),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_51),
.A2(n_91),
.B(n_123),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_51),
.A2(n_123),
.B(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_51),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_51),
.A2(n_90),
.B1(n_185),
.B2(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_51),
.A2(n_90),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_51),
.A2(n_90),
.B1(n_194),
.B2(n_204),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_66),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_62),
.B(n_64),
.Y(n_54)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_55),
.B(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_55),
.A2(n_105),
.B1(n_108),
.B2(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_55),
.A2(n_108),
.B1(n_160),
.B2(n_179),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_56),
.A2(n_130),
.B(n_131),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_56),
.A2(n_106),
.B1(n_159),
.B2(n_161),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_60),
.A2(n_61),
.B1(n_75),
.B2(n_76),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_L g101 ( 
.A1(n_60),
.A2(n_76),
.B(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

HAxp5_ASAP7_75t_SL g179 ( 
.A(n_61),
.B(n_102),
.CON(n_179),
.SN(n_179)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_62),
.B(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_73),
.B1(n_78),
.B2(n_80),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_67),
.Y(n_114)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_72),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_73),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_73),
.A2(n_80),
.B1(n_112),
.B2(n_146),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_77),
.A2(n_110),
.B1(n_111),
.B2(n_114),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_78),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_80),
.B(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_88),
.B2(n_92),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_92),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_88),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_90),
.B(n_151),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_93),
.B(n_246),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_103),
.C(n_109),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_94),
.A2(n_95),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_96),
.A2(n_97),
.B1(n_100),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_100),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_103),
.B(n_109),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_106),
.B(n_107),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_110),
.A2(n_134),
.B(n_135),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_139),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_124),
.B1(n_137),
.B2(n_138),
.Y(n_116)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_133),
.Y(n_128)
);

O2A1O1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_169),
.B(n_244),
.C(n_248),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_162),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_143),
.B(n_162),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_152),
.C(n_154),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_144),
.B(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_148),
.C(n_150),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_149),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_152),
.B(n_154),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.C(n_158),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_158),
.B(n_188),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_163),
.B(n_167),
.C(n_168),
.Y(n_247)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_239),
.B(n_243),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_195),
.B(n_238),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_190),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_174),
.B(n_190),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_187),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_182),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_176),
.B(n_182),
.C(n_187),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_177),
.B(n_181),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_184),
.B(n_186),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.C(n_193),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_191),
.B(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_192),
.B(n_193),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_233),
.B(n_237),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_223),
.B(n_232),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_212),
.B(n_222),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_207),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_207),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_202),
.B1(n_205),
.B2(n_206),
.Y(n_199)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_200),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_202),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_205),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_218),
.B(n_221),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_220),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_225),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_228),
.C(n_231),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_230),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_236),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_242),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_247),
.Y(n_248)
);


endmodule