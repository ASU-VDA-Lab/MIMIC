module fake_netlist_6_4540_n_1414 (n_52, n_1, n_91, n_326, n_256, n_209, n_63, n_223, n_278, n_341, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_338, n_56, n_119, n_235, n_147, n_191, n_340, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_334, n_53, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_231, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_317, n_149, n_90, n_24, n_54, n_328, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1414);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_341;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_338;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_334;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_231;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_317;
input n_149;
input n_90;
input n_24;
input n_54;
input n_328;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1414;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1370;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1393;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_606;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_1368;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1382;
wire n_1372;
wire n_505;
wire n_1339;
wire n_537;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_351;
wire n_385;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_828;
wire n_607;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1316;
wire n_1287;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1177;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_1311;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_177),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_271),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_285),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_194),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_287),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_332),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_4),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_191),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_39),
.Y(n_350)
);

BUFx10_ASAP7_75t_L g351 ( 
.A(n_32),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_51),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_172),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_79),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_299),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_171),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_89),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_173),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_180),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_313),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_138),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_129),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_224),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_201),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_240),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_320),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_170),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_126),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_60),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_65),
.Y(n_370)
);

BUFx10_ASAP7_75t_L g371 ( 
.A(n_133),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_288),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_82),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_28),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_161),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_30),
.Y(n_376)
);

BUFx8_ASAP7_75t_SL g377 ( 
.A(n_157),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_265),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_17),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_69),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_336),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_251),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_279),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_211),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_216),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_75),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_338),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_237),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_122),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_319),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_228),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_88),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_227),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_147),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_114),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_325),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_124),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_199),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_167),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_131),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_25),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_3),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_14),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_286),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_92),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_337),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_209),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_309),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_31),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_59),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_72),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_7),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_6),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_329),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_137),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_294),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_58),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_29),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_328),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_66),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_64),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_80),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_73),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_304),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_64),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_195),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_142),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_9),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_108),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_289),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_90),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_306),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_30),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_109),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_217),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_66),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_67),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_53),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_84),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_35),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_2),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_322),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_232),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_295),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_7),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_65),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_107),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_231),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_193),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_277),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_99),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_5),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_339),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_149),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_15),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_110),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_140),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_283),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_307),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_242),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_74),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_290),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_234),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_247),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_221),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_61),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_233),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_5),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_91),
.Y(n_469)
);

BUFx10_ASAP7_75t_L g470 ( 
.A(n_19),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_85),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_267),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_113),
.Y(n_473)
);

INVxp33_ASAP7_75t_SL g474 ( 
.A(n_278),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_117),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_192),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_127),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_327),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_215),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_128),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_77),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_93),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_69),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_248),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_229),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_204),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_87),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_324),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_61),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_280),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_15),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_6),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_31),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_183),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_206),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_303),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_218),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_56),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g499 ( 
.A(n_50),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_321),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_202),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_21),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_186),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_315),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_41),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_17),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_22),
.Y(n_507)
);

CKINVDCx14_ASAP7_75t_R g508 ( 
.A(n_62),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_102),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_260),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_68),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_253),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_104),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_62),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_0),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_219),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_333),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_10),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_264),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_123),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_81),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_293),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_120),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_145),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_301),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_36),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_323),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_116),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_26),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_163),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_335),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_43),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_26),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_438),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_508),
.B(n_0),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_343),
.B(n_1),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_438),
.Y(n_537)
);

INVx5_ASAP7_75t_L g538 ( 
.A(n_439),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_439),
.Y(n_539)
);

BUFx12f_ASAP7_75t_L g540 ( 
.A(n_351),
.Y(n_540)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_439),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_508),
.B(n_1),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_438),
.B(n_2),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_375),
.B(n_3),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_375),
.B(n_4),
.Y(n_545)
);

CKINVDCx16_ASAP7_75t_R g546 ( 
.A(n_432),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_438),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_379),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_439),
.Y(n_549)
);

INVx4_ASAP7_75t_L g550 ( 
.A(n_458),
.Y(n_550)
);

INVx5_ASAP7_75t_L g551 ( 
.A(n_458),
.Y(n_551)
);

INVx5_ASAP7_75t_L g552 ( 
.A(n_458),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_403),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_410),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_412),
.Y(n_555)
);

BUFx12f_ASAP7_75t_L g556 ( 
.A(n_351),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_382),
.B(n_8),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_370),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_370),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_392),
.B(n_8),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_437),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_446),
.Y(n_562)
);

INVx5_ASAP7_75t_L g563 ( 
.A(n_458),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_343),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_474),
.B(n_9),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_408),
.B(n_10),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_362),
.B(n_11),
.Y(n_567)
);

CKINVDCx16_ASAP7_75t_R g568 ( 
.A(n_349),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_362),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_407),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_407),
.B(n_11),
.Y(n_571)
);

NOR2x1_ASAP7_75t_L g572 ( 
.A(n_427),
.B(n_76),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_408),
.B(n_12),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_427),
.B(n_12),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_413),
.B(n_13),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_487),
.B(n_13),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_452),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_462),
.B(n_14),
.Y(n_578)
);

INVx5_ASAP7_75t_L g579 ( 
.A(n_371),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_462),
.B(n_16),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_444),
.Y(n_581)
);

INVx5_ASAP7_75t_L g582 ( 
.A(n_371),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_348),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_444),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_461),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_494),
.B(n_16),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_461),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_452),
.Y(n_588)
);

INVxp67_ASAP7_75t_L g589 ( 
.A(n_445),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_497),
.B(n_18),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_497),
.B(n_18),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_371),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_498),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_513),
.B(n_19),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_377),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_474),
.B(n_20),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_361),
.B(n_20),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_342),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_501),
.B(n_21),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_498),
.Y(n_600)
);

NOR2x1_ASAP7_75t_L g601 ( 
.A(n_513),
.B(n_78),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_455),
.Y(n_602)
);

INVx5_ASAP7_75t_L g603 ( 
.A(n_377),
.Y(n_603)
);

BUFx8_ASAP7_75t_SL g604 ( 
.A(n_413),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_351),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_470),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_345),
.B(n_22),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_468),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_489),
.B(n_502),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_511),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_470),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_526),
.B(n_23),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_355),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_358),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_350),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_365),
.B(n_23),
.Y(n_616)
);

INVx5_ASAP7_75t_L g617 ( 
.A(n_470),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_383),
.B(n_24),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_528),
.B(n_24),
.Y(n_619)
);

BUFx8_ASAP7_75t_SL g620 ( 
.A(n_417),
.Y(n_620)
);

INVx5_ASAP7_75t_L g621 ( 
.A(n_344),
.Y(n_621)
);

AND2x6_ASAP7_75t_L g622 ( 
.A(n_385),
.B(n_83),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_349),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_389),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_391),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_492),
.B(n_25),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_394),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_346),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_352),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_395),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_397),
.B(n_27),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_347),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_398),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_406),
.B(n_27),
.Y(n_634)
);

OAI22xp33_ASAP7_75t_SL g635 ( 
.A1(n_575),
.A2(n_535),
.B1(n_592),
.B2(n_560),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_565),
.A2(n_386),
.B1(n_396),
.B2(n_360),
.Y(n_636)
);

AO22x2_ASAP7_75t_L g637 ( 
.A1(n_536),
.A2(n_506),
.B1(n_499),
.B2(n_424),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_583),
.B(n_353),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_547),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_534),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_SL g641 ( 
.A1(n_568),
.A2(n_441),
.B1(n_483),
.B2(n_417),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_537),
.Y(n_642)
);

OAI22xp33_ASAP7_75t_SL g643 ( 
.A1(n_575),
.A2(n_374),
.B1(n_376),
.B2(n_369),
.Y(n_643)
);

OAI22xp33_ASAP7_75t_SL g644 ( 
.A1(n_535),
.A2(n_533),
.B1(n_401),
.B2(n_402),
.Y(n_644)
);

AO22x2_ASAP7_75t_L g645 ( 
.A1(n_536),
.A2(n_426),
.B1(n_430),
.B2(n_414),
.Y(n_645)
);

OAI22xp33_ASAP7_75t_SL g646 ( 
.A1(n_592),
.A2(n_532),
.B1(n_409),
.B2(n_411),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_596),
.A2(n_386),
.B1(n_396),
.B2(n_360),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_615),
.B(n_354),
.Y(n_648)
);

OAI22xp33_ASAP7_75t_SL g649 ( 
.A1(n_557),
.A2(n_418),
.B1(n_420),
.B2(n_380),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_547),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_SL g651 ( 
.A1(n_623),
.A2(n_441),
.B1(n_483),
.B2(n_443),
.Y(n_651)
);

AOI22xp5_ASAP7_75t_L g652 ( 
.A1(n_546),
.A2(n_443),
.B1(n_510),
.B2(n_435),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_603),
.B(n_356),
.Y(n_653)
);

AO22x2_ASAP7_75t_L g654 ( 
.A1(n_590),
.A2(n_442),
.B1(n_453),
.B2(n_434),
.Y(n_654)
);

AO22x2_ASAP7_75t_L g655 ( 
.A1(n_590),
.A2(n_456),
.B1(n_459),
.B2(n_454),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_603),
.B(n_357),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_628),
.B(n_460),
.Y(n_657)
);

OAI22xp33_ASAP7_75t_L g658 ( 
.A1(n_605),
.A2(n_423),
.B1(n_425),
.B2(n_421),
.Y(n_658)
);

OAI22xp33_ASAP7_75t_SL g659 ( 
.A1(n_557),
.A2(n_433),
.B1(n_436),
.B2(n_428),
.Y(n_659)
);

OAI22xp33_ASAP7_75t_L g660 ( 
.A1(n_605),
.A2(n_440),
.B1(n_491),
.B2(n_466),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_SL g661 ( 
.A1(n_597),
.A2(n_510),
.B1(n_435),
.B2(n_505),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_549),
.Y(n_662)
);

OAI22xp33_ASAP7_75t_L g663 ( 
.A1(n_606),
.A2(n_616),
.B1(n_545),
.B2(n_566),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_SL g664 ( 
.A1(n_597),
.A2(n_507),
.B1(n_514),
.B2(n_493),
.Y(n_664)
);

OAI22xp33_ASAP7_75t_L g665 ( 
.A1(n_606),
.A2(n_518),
.B1(n_529),
.B2(n_515),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_549),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_542),
.B(n_463),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_598),
.B(n_465),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_549),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_603),
.B(n_359),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_569),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_603),
.B(n_363),
.Y(n_672)
);

OA22x2_ASAP7_75t_L g673 ( 
.A1(n_611),
.A2(n_476),
.B1(n_477),
.B2(n_467),
.Y(n_673)
);

OAI22xp33_ASAP7_75t_SL g674 ( 
.A1(n_579),
.A2(n_488),
.B1(n_495),
.B2(n_480),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_617),
.B(n_579),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_629),
.B(n_364),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_587),
.B(n_366),
.Y(n_677)
);

OAI22xp33_ASAP7_75t_SL g678 ( 
.A1(n_579),
.A2(n_516),
.B1(n_517),
.B2(n_496),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_617),
.B(n_367),
.Y(n_679)
);

OAI22xp33_ASAP7_75t_L g680 ( 
.A1(n_616),
.A2(n_524),
.B1(n_525),
.B2(n_519),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_628),
.B(n_530),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_569),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_569),
.Y(n_683)
);

OR2x6_ASAP7_75t_L g684 ( 
.A(n_595),
.B(n_531),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_570),
.Y(n_685)
);

NOR2x1p5_ASAP7_75t_L g686 ( 
.A(n_540),
.B(n_368),
.Y(n_686)
);

OAI22xp33_ASAP7_75t_SL g687 ( 
.A1(n_579),
.A2(n_373),
.B1(n_378),
.B2(n_372),
.Y(n_687)
);

OAI22xp33_ASAP7_75t_L g688 ( 
.A1(n_544),
.A2(n_384),
.B1(n_387),
.B2(n_381),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_564),
.B(n_584),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_570),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_570),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_599),
.A2(n_390),
.B1(n_393),
.B2(n_388),
.Y(n_692)
);

AO22x2_ASAP7_75t_L g693 ( 
.A1(n_591),
.A2(n_32),
.B1(n_28),
.B2(n_29),
.Y(n_693)
);

OAI22xp33_ASAP7_75t_L g694 ( 
.A1(n_544),
.A2(n_400),
.B1(n_404),
.B2(n_399),
.Y(n_694)
);

OAI22xp33_ASAP7_75t_L g695 ( 
.A1(n_545),
.A2(n_415),
.B1(n_416),
.B2(n_405),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_581),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_581),
.Y(n_697)
);

BUFx2_ASAP7_75t_L g698 ( 
.A(n_556),
.Y(n_698)
);

NOR2x1p5_ASAP7_75t_L g699 ( 
.A(n_566),
.B(n_419),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_599),
.A2(n_429),
.B1(n_431),
.B2(n_422),
.Y(n_700)
);

OR2x6_ASAP7_75t_L g701 ( 
.A(n_612),
.B(n_33),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_561),
.Y(n_702)
);

OAI22xp5_ASAP7_75t_SL g703 ( 
.A1(n_619),
.A2(n_448),
.B1(n_449),
.B2(n_447),
.Y(n_703)
);

OAI22xp33_ASAP7_75t_L g704 ( 
.A1(n_573),
.A2(n_451),
.B1(n_457),
.B2(n_450),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_562),
.Y(n_705)
);

XOR2xp5_ASAP7_75t_L g706 ( 
.A(n_626),
.B(n_464),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_632),
.B(n_469),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_619),
.A2(n_472),
.B1(n_473),
.B2(n_471),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_576),
.A2(n_478),
.B1(n_479),
.B2(n_475),
.Y(n_709)
);

AND2x4_ASAP7_75t_L g710 ( 
.A(n_617),
.B(n_481),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_602),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_617),
.B(n_482),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_610),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_581),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_585),
.Y(n_715)
);

OAI22xp33_ASAP7_75t_L g716 ( 
.A1(n_573),
.A2(n_527),
.B1(n_523),
.B2(n_522),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_582),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_582),
.Y(n_718)
);

OAI22xp33_ASAP7_75t_L g719 ( 
.A1(n_578),
.A2(n_521),
.B1(n_520),
.B2(n_512),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_668),
.B(n_564),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_685),
.Y(n_721)
);

AND2x2_ASAP7_75t_SL g722 ( 
.A(n_636),
.B(n_591),
.Y(n_722)
);

NAND2xp33_ASAP7_75t_SL g723 ( 
.A(n_664),
.B(n_567),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_685),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_666),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_666),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_662),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_669),
.Y(n_728)
);

BUFx2_ASAP7_75t_L g729 ( 
.A(n_706),
.Y(n_729)
);

XOR2xp5_ASAP7_75t_L g730 ( 
.A(n_652),
.B(n_484),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_671),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_690),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_703),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_696),
.Y(n_734)
);

NAND2x1p5_ASAP7_75t_L g735 ( 
.A(n_699),
.B(n_572),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_663),
.B(n_689),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_640),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_677),
.B(n_582),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_697),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_667),
.B(n_621),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_642),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_714),
.Y(n_742)
);

INVx4_ASAP7_75t_L g743 ( 
.A(n_707),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_715),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_682),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_700),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_683),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_691),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_650),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_639),
.Y(n_750)
);

NOR2x1_ASAP7_75t_L g751 ( 
.A(n_675),
.B(n_539),
.Y(n_751)
);

BUFx8_ASAP7_75t_L g752 ( 
.A(n_698),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_638),
.B(n_582),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_639),
.Y(n_754)
);

AND2x6_ASAP7_75t_L g755 ( 
.A(n_676),
.B(n_594),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_702),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_702),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_648),
.B(n_584),
.Y(n_758)
);

AOI21x1_ASAP7_75t_L g759 ( 
.A1(n_667),
.A2(n_624),
.B(n_601),
.Y(n_759)
);

NOR2xp67_ASAP7_75t_L g760 ( 
.A(n_692),
.B(n_621),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_705),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_717),
.B(n_585),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_718),
.B(n_585),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_653),
.Y(n_764)
);

INVxp67_ASAP7_75t_SL g765 ( 
.A(n_705),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_711),
.Y(n_766)
);

AND2x6_ASAP7_75t_L g767 ( 
.A(n_656),
.B(n_594),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_711),
.Y(n_768)
);

XOR2xp5_ASAP7_75t_L g769 ( 
.A(n_651),
.B(n_485),
.Y(n_769)
);

XNOR2x1_ASAP7_75t_L g770 ( 
.A(n_647),
.B(n_604),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_713),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_713),
.Y(n_772)
);

AND2x2_ASAP7_75t_SL g773 ( 
.A(n_707),
.B(n_571),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_673),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_710),
.B(n_589),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_710),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_658),
.B(n_621),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_657),
.B(n_621),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_660),
.B(n_574),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_645),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_670),
.A2(n_551),
.B(n_538),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_641),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_645),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_665),
.B(n_576),
.Y(n_784)
);

INVxp67_ASAP7_75t_SL g785 ( 
.A(n_681),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_654),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_708),
.B(n_586),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_654),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_701),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_684),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_655),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_709),
.A2(n_622),
.B(n_618),
.Y(n_792)
);

AND2x4_ASAP7_75t_L g793 ( 
.A(n_684),
.B(n_607),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_655),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_672),
.Y(n_795)
);

XNOR2x2_ASAP7_75t_L g796 ( 
.A(n_693),
.B(n_586),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_701),
.Y(n_797)
);

XNOR2xp5_ASAP7_75t_L g798 ( 
.A(n_661),
.B(n_686),
.Y(n_798)
);

INVxp33_ASAP7_75t_L g799 ( 
.A(n_637),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_693),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_674),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_678),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_688),
.B(n_613),
.Y(n_803)
);

INVxp67_ASAP7_75t_SL g804 ( 
.A(n_680),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_637),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_694),
.B(n_614),
.Y(n_806)
);

INVx3_ASAP7_75t_R g807 ( 
.A(n_646),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_644),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_756),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_776),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_757),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_754),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_761),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_785),
.B(n_695),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_785),
.B(n_558),
.Y(n_815)
);

INVx1_ASAP7_75t_SL g816 ( 
.A(n_775),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_720),
.B(n_635),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_720),
.B(n_704),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_758),
.B(n_589),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_736),
.B(n_773),
.Y(n_820)
);

AND2x2_ASAP7_75t_SL g821 ( 
.A(n_722),
.B(n_607),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_773),
.B(n_716),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_776),
.B(n_719),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_736),
.B(n_765),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_776),
.B(n_792),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_766),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_795),
.B(n_622),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_808),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_768),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_754),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_765),
.B(n_558),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_746),
.B(n_643),
.Y(n_832)
);

INVx1_ASAP7_75t_SL g833 ( 
.A(n_729),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_771),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_750),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_776),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_804),
.B(n_774),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_772),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_767),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_737),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_753),
.B(n_588),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_737),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_743),
.B(n_722),
.Y(n_843)
);

AND2x2_ASAP7_75t_SL g844 ( 
.A(n_787),
.B(n_618),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_804),
.B(n_588),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_764),
.B(n_600),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_764),
.B(n_600),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_787),
.B(n_649),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_755),
.B(n_622),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_794),
.B(n_634),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_780),
.B(n_783),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_741),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_755),
.B(n_622),
.Y(n_853)
);

INVxp67_ASAP7_75t_L g854 ( 
.A(n_784),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_743),
.B(n_548),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_741),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_755),
.B(n_622),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_749),
.Y(n_858)
);

INVx4_ASAP7_75t_L g859 ( 
.A(n_767),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_762),
.B(n_553),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_767),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_784),
.B(n_659),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_767),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_767),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_803),
.B(n_634),
.Y(n_865)
);

AND2x6_ASAP7_75t_L g866 ( 
.A(n_800),
.B(n_578),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_732),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_779),
.B(n_687),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_755),
.B(n_679),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_727),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_786),
.B(n_554),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_803),
.B(n_486),
.Y(n_872)
);

BUFx24_ASAP7_75t_L g873 ( 
.A(n_796),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_733),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_779),
.B(n_712),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_777),
.B(n_620),
.Y(n_876)
);

INVxp67_ASAP7_75t_SL g877 ( 
.A(n_742),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_728),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_806),
.B(n_625),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_747),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_725),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_755),
.B(n_630),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_777),
.B(n_631),
.Y(n_883)
);

CKINVDCx14_ASAP7_75t_R g884 ( 
.A(n_723),
.Y(n_884)
);

AND2x2_ASAP7_75t_SL g885 ( 
.A(n_806),
.B(n_580),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_763),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_793),
.B(n_555),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_788),
.B(n_608),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_791),
.B(n_801),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_735),
.B(n_490),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_742),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_723),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_802),
.B(n_631),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_738),
.B(n_627),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_731),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_734),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_735),
.B(n_543),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_789),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_778),
.B(n_627),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_726),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_740),
.B(n_627),
.Y(n_901)
);

OR2x2_ASAP7_75t_L g902 ( 
.A(n_805),
.B(n_612),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_739),
.B(n_609),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_824),
.B(n_797),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_SL g905 ( 
.A(n_821),
.B(n_782),
.Y(n_905)
);

CKINVDCx16_ASAP7_75t_R g906 ( 
.A(n_884),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_812),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_812),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_854),
.B(n_799),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_830),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_824),
.B(n_885),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_816),
.B(n_799),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_830),
.Y(n_913)
);

NAND2xp33_ASAP7_75t_L g914 ( 
.A(n_810),
.B(n_861),
.Y(n_914)
);

AO21x2_ASAP7_75t_L g915 ( 
.A1(n_825),
.A2(n_759),
.B(n_760),
.Y(n_915)
);

OR2x6_ASAP7_75t_L g916 ( 
.A(n_892),
.B(n_789),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_810),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_SL g918 ( 
.A(n_821),
.B(n_782),
.Y(n_918)
);

INVxp67_ASAP7_75t_L g919 ( 
.A(n_819),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_830),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_846),
.Y(n_921)
);

NAND2x1p5_ASAP7_75t_L g922 ( 
.A(n_861),
.B(n_863),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_835),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_886),
.B(n_793),
.Y(n_924)
);

CKINVDCx16_ASAP7_75t_R g925 ( 
.A(n_884),
.Y(n_925)
);

BUFx2_ASAP7_75t_L g926 ( 
.A(n_898),
.Y(n_926)
);

BUFx2_ASAP7_75t_SL g927 ( 
.A(n_846),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_835),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_886),
.B(n_745),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_885),
.B(n_744),
.Y(n_930)
);

BUFx2_ASAP7_75t_L g931 ( 
.A(n_837),
.Y(n_931)
);

INVx5_ASAP7_75t_L g932 ( 
.A(n_861),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_867),
.Y(n_933)
);

INVxp67_ASAP7_75t_SL g934 ( 
.A(n_810),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_837),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_845),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_871),
.B(n_748),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_851),
.Y(n_938)
);

AND2x2_ASAP7_75t_SL g939 ( 
.A(n_844),
.B(n_770),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_871),
.B(n_721),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_815),
.B(n_831),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_810),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_875),
.B(n_730),
.Y(n_943)
);

OR2x6_ASAP7_75t_L g944 ( 
.A(n_843),
.B(n_724),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_847),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_820),
.B(n_807),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_815),
.B(n_769),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_840),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_831),
.B(n_847),
.Y(n_949)
);

NOR2x1_ASAP7_75t_L g950 ( 
.A(n_836),
.B(n_890),
.Y(n_950)
);

NOR2x1_ASAP7_75t_SL g951 ( 
.A(n_861),
.B(n_538),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_865),
.B(n_751),
.Y(n_952)
);

BUFx2_ASAP7_75t_L g953 ( 
.A(n_845),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_871),
.B(n_790),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_874),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_851),
.Y(n_956)
);

OR2x2_ASAP7_75t_L g957 ( 
.A(n_833),
.B(n_798),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_842),
.Y(n_958)
);

NOR2x1p5_ASAP7_75t_SL g959 ( 
.A(n_881),
.B(n_781),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_841),
.B(n_609),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_820),
.B(n_752),
.Y(n_961)
);

NOR2x1_ASAP7_75t_L g962 ( 
.A(n_836),
.B(n_580),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_865),
.B(n_543),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_817),
.B(n_633),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_867),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_852),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_879),
.B(n_633),
.Y(n_967)
);

INVx8_ASAP7_75t_L g968 ( 
.A(n_866),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_856),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_883),
.B(n_559),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_851),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_879),
.B(n_633),
.Y(n_972)
);

INVxp67_ASAP7_75t_SL g973 ( 
.A(n_825),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_818),
.B(n_500),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_809),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_926),
.Y(n_976)
);

BUFx2_ASAP7_75t_L g977 ( 
.A(n_945),
.Y(n_977)
);

BUFx2_ASAP7_75t_R g978 ( 
.A(n_955),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_971),
.B(n_811),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_954),
.Y(n_980)
);

INVx5_ASAP7_75t_L g981 ( 
.A(n_968),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_954),
.Y(n_982)
);

BUFx3_ASAP7_75t_L g983 ( 
.A(n_931),
.Y(n_983)
);

BUFx10_ASAP7_75t_L g984 ( 
.A(n_961),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_922),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_917),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_907),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_938),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_971),
.B(n_813),
.Y(n_989)
);

INVx8_ASAP7_75t_L g990 ( 
.A(n_968),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_944),
.Y(n_991)
);

AOI22xp33_ASAP7_75t_SL g992 ( 
.A1(n_943),
.A2(n_844),
.B1(n_832),
.B2(n_868),
.Y(n_992)
);

NAND2xp33_ASAP7_75t_L g993 ( 
.A(n_932),
.B(n_863),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_938),
.Y(n_994)
);

BUFx12f_ASAP7_75t_L g995 ( 
.A(n_916),
.Y(n_995)
);

INVxp67_ASAP7_75t_SL g996 ( 
.A(n_934),
.Y(n_996)
);

INVx3_ASAP7_75t_SL g997 ( 
.A(n_906),
.Y(n_997)
);

INVx2_ASAP7_75t_SL g998 ( 
.A(n_917),
.Y(n_998)
);

INVx11_ASAP7_75t_L g999 ( 
.A(n_927),
.Y(n_999)
);

INVx4_ASAP7_75t_L g1000 ( 
.A(n_917),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_941),
.B(n_814),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_956),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_908),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_942),
.Y(n_1004)
);

INVx4_ASAP7_75t_L g1005 ( 
.A(n_942),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_942),
.Y(n_1006)
);

CKINVDCx11_ASAP7_75t_R g1007 ( 
.A(n_925),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_932),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_956),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_949),
.B(n_970),
.Y(n_1010)
);

INVx6_ASAP7_75t_L g1011 ( 
.A(n_932),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_975),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_923),
.Y(n_1013)
);

BUFx12f_ASAP7_75t_L g1014 ( 
.A(n_916),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_928),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_944),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_932),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_944),
.Y(n_1018)
);

BUFx4_ASAP7_75t_SL g1019 ( 
.A(n_916),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_911),
.B(n_897),
.Y(n_1020)
);

INVx1_ASAP7_75t_SL g1021 ( 
.A(n_936),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_910),
.Y(n_1022)
);

CKINVDCx16_ASAP7_75t_R g1023 ( 
.A(n_957),
.Y(n_1023)
);

AOI22xp33_ASAP7_75t_L g1024 ( 
.A1(n_911),
.A2(n_848),
.B1(n_862),
.B2(n_822),
.Y(n_1024)
);

CKINVDCx16_ASAP7_75t_R g1025 ( 
.A(n_905),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_948),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_953),
.B(n_897),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_958),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_921),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_966),
.Y(n_1030)
);

BUFx12f_ASAP7_75t_L g1031 ( 
.A(n_924),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_968),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_960),
.B(n_963),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_935),
.B(n_848),
.Y(n_1034)
);

BUFx2_ASAP7_75t_L g1035 ( 
.A(n_976),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_1003),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1012),
.Y(n_1037)
);

CKINVDCx11_ASAP7_75t_R g1038 ( 
.A(n_997),
.Y(n_1038)
);

INVx1_ASAP7_75t_SL g1039 ( 
.A(n_1021),
.Y(n_1039)
);

CKINVDCx11_ASAP7_75t_R g1040 ( 
.A(n_997),
.Y(n_1040)
);

INVx4_ASAP7_75t_L g1041 ( 
.A(n_1011),
.Y(n_1041)
);

AOI22xp33_ASAP7_75t_SL g1042 ( 
.A1(n_1025),
.A2(n_905),
.B1(n_918),
.B2(n_939),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_992),
.A2(n_918),
.B1(n_822),
.B2(n_862),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_986),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1026),
.Y(n_1045)
);

BUFx8_ASAP7_75t_L g1046 ( 
.A(n_977),
.Y(n_1046)
);

OAI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_1033),
.A2(n_874),
.B1(n_947),
.B2(n_919),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_978),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_SL g1049 ( 
.A1(n_1024),
.A2(n_946),
.B(n_873),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_1001),
.A2(n_904),
.B1(n_963),
.B2(n_934),
.Y(n_1050)
);

BUFx2_ASAP7_75t_L g1051 ( 
.A(n_976),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_983),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_986),
.Y(n_1053)
);

CKINVDCx20_ASAP7_75t_R g1054 ( 
.A(n_1007),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1028),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_1020),
.B(n_964),
.Y(n_1056)
);

INVx6_ASAP7_75t_L g1057 ( 
.A(n_995),
.Y(n_1057)
);

AOI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_1020),
.A2(n_872),
.B1(n_909),
.B2(n_828),
.Y(n_1058)
);

INVx3_ASAP7_75t_SL g1059 ( 
.A(n_1023),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_1027),
.A2(n_872),
.B1(n_876),
.B2(n_919),
.Y(n_1060)
);

INVx6_ASAP7_75t_L g1061 ( 
.A(n_995),
.Y(n_1061)
);

INVx1_ASAP7_75t_SL g1062 ( 
.A(n_977),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1030),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_1011),
.Y(n_1064)
);

INVx2_ASAP7_75t_SL g1065 ( 
.A(n_999),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_1027),
.A2(n_924),
.B1(n_937),
.B2(n_866),
.Y(n_1066)
);

CKINVDCx11_ASAP7_75t_R g1067 ( 
.A(n_1007),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_1010),
.A2(n_904),
.B1(n_873),
.B2(n_967),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1003),
.Y(n_1069)
);

CKINVDCx11_ASAP7_75t_R g1070 ( 
.A(n_1014),
.Y(n_1070)
);

AOI22xp33_ASAP7_75t_L g1071 ( 
.A1(n_1034),
.A2(n_937),
.B1(n_866),
.B2(n_823),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1013),
.Y(n_1072)
);

AOI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_1034),
.A2(n_866),
.B1(n_823),
.B2(n_912),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_987),
.Y(n_1074)
);

OAI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_987),
.A2(n_973),
.B(n_964),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1022),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_986),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1015),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_1031),
.A2(n_866),
.B1(n_940),
.B2(n_890),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1022),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_1011),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_986),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_988),
.Y(n_1083)
);

AOI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_979),
.A2(n_950),
.B1(n_974),
.B2(n_952),
.Y(n_1084)
);

AOI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_979),
.A2(n_974),
.B1(n_952),
.B2(n_855),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_994),
.Y(n_1086)
);

OAI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_996),
.A2(n_967),
.B1(n_972),
.B2(n_893),
.Y(n_1087)
);

INVx2_ASAP7_75t_SL g1088 ( 
.A(n_999),
.Y(n_1088)
);

INVx6_ASAP7_75t_L g1089 ( 
.A(n_1014),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1002),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_1009),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_1043),
.A2(n_983),
.B1(n_984),
.B2(n_991),
.Y(n_1092)
);

NOR2xp67_ASAP7_75t_SL g1093 ( 
.A(n_1048),
.B(n_981),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_1042),
.A2(n_1047),
.B1(n_1068),
.B2(n_1060),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_1039),
.B(n_984),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_1042),
.A2(n_1016),
.B1(n_1018),
.B2(n_991),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_1068),
.A2(n_984),
.B1(n_1018),
.B2(n_1016),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1058),
.B(n_1029),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_1062),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_1039),
.B(n_980),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1056),
.B(n_889),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_1046),
.Y(n_1102)
);

BUFx4f_ASAP7_75t_SL g1103 ( 
.A(n_1054),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_1071),
.A2(n_989),
.B1(n_979),
.B2(n_1031),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1037),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_1073),
.A2(n_989),
.B1(n_930),
.B2(n_962),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_1059),
.B(n_980),
.Y(n_1107)
);

AOI22xp33_ASAP7_75t_L g1108 ( 
.A1(n_1056),
.A2(n_989),
.B1(n_930),
.B2(n_866),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_1066),
.A2(n_826),
.B1(n_834),
.B2(n_829),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1036),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_1085),
.A2(n_838),
.B1(n_969),
.B2(n_858),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1045),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1076),
.Y(n_1113)
);

AOI22xp33_ASAP7_75t_SL g1114 ( 
.A1(n_1046),
.A2(n_752),
.B1(n_973),
.B2(n_982),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1055),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1049),
.A2(n_982),
.B1(n_902),
.B2(n_971),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1050),
.B(n_972),
.Y(n_1117)
);

AOI22xp33_ASAP7_75t_SL g1118 ( 
.A1(n_1050),
.A2(n_981),
.B1(n_914),
.B2(n_887),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_SL g1119 ( 
.A1(n_1049),
.A2(n_860),
.B(n_869),
.Y(n_1119)
);

OR2x2_ASAP7_75t_L g1120 ( 
.A(n_1062),
.B(n_903),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1063),
.Y(n_1121)
);

OR2x2_ASAP7_75t_L g1122 ( 
.A(n_1086),
.B(n_1091),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_1052),
.B(n_903),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1084),
.B(n_903),
.Y(n_1124)
);

BUFx12f_ASAP7_75t_L g1125 ( 
.A(n_1038),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_1079),
.A2(n_915),
.B1(n_929),
.B2(n_878),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1035),
.A2(n_929),
.B1(n_981),
.B2(n_895),
.Y(n_1127)
);

OAI222xp33_ASAP7_75t_L g1128 ( 
.A1(n_1087),
.A2(n_933),
.B1(n_965),
.B2(n_920),
.C1(n_913),
.C2(n_981),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_1040),
.A2(n_915),
.B1(n_896),
.B2(n_940),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_1044),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1051),
.B(n_888),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_1041),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_1067),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_1044),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1072),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_1057),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_SL g1137 ( 
.A1(n_1057),
.A2(n_981),
.B1(n_993),
.B2(n_990),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1083),
.B(n_888),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1078),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_1061),
.A2(n_880),
.B1(n_870),
.B2(n_881),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_1061),
.A2(n_880),
.B1(n_870),
.B2(n_900),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1089),
.A2(n_1087),
.B1(n_1088),
.B2(n_1065),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_1075),
.Y(n_1143)
);

OAI21xp5_ASAP7_75t_SL g1144 ( 
.A1(n_1075),
.A2(n_888),
.B(n_850),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1069),
.Y(n_1145)
);

CKINVDCx20_ASAP7_75t_R g1146 ( 
.A(n_1070),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1089),
.A2(n_1090),
.B1(n_895),
.B2(n_894),
.Y(n_1147)
);

OR2x2_ASAP7_75t_L g1148 ( 
.A(n_1074),
.B(n_901),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_1080),
.Y(n_1149)
);

AOI22xp33_ASAP7_75t_L g1150 ( 
.A1(n_1064),
.A2(n_900),
.B1(n_882),
.B2(n_863),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_SL g1151 ( 
.A1(n_1041),
.A2(n_993),
.B1(n_990),
.B2(n_1011),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1044),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1094),
.A2(n_1081),
.B1(n_1064),
.B2(n_899),
.Y(n_1153)
);

AOI22xp33_ASAP7_75t_L g1154 ( 
.A1(n_1124),
.A2(n_1081),
.B1(n_827),
.B2(n_863),
.Y(n_1154)
);

OAI221xp5_ASAP7_75t_L g1155 ( 
.A1(n_1119),
.A2(n_503),
.B1(n_504),
.B2(n_509),
.C(n_559),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1097),
.A2(n_985),
.B1(n_922),
.B2(n_1032),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1101),
.B(n_1053),
.Y(n_1157)
);

NAND3xp33_ASAP7_75t_L g1158 ( 
.A(n_1129),
.B(n_593),
.C(n_577),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1116),
.A2(n_864),
.B1(n_839),
.B2(n_985),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1096),
.A2(n_864),
.B1(n_839),
.B2(n_985),
.Y(n_1160)
);

AOI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1142),
.A2(n_864),
.B1(n_839),
.B2(n_859),
.Y(n_1161)
);

AOI22xp33_ASAP7_75t_SL g1162 ( 
.A1(n_1098),
.A2(n_990),
.B1(n_1032),
.B2(n_1019),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1099),
.B(n_1053),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_1104),
.A2(n_891),
.B1(n_859),
.B2(n_1032),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1092),
.A2(n_1032),
.B1(n_1006),
.B2(n_998),
.Y(n_1165)
);

NOR3xp33_ASAP7_75t_L g1166 ( 
.A(n_1144),
.B(n_593),
.C(n_577),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1099),
.B(n_1053),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_SL g1168 ( 
.A1(n_1095),
.A2(n_990),
.B1(n_1032),
.B2(n_1077),
.Y(n_1168)
);

NAND3xp33_ASAP7_75t_L g1169 ( 
.A(n_1147),
.B(n_891),
.C(n_1077),
.Y(n_1169)
);

AOI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1111),
.A2(n_850),
.B1(n_859),
.B2(n_891),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1118),
.A2(n_1108),
.B1(n_1106),
.B2(n_1126),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1143),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1143),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1122),
.B(n_1077),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1145),
.Y(n_1175)
);

AOI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1109),
.A2(n_1138),
.B1(n_1118),
.B2(n_1114),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_1100),
.A2(n_853),
.B1(n_857),
.B2(n_849),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1110),
.B(n_1082),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1114),
.A2(n_1082),
.B1(n_998),
.B2(n_1006),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1107),
.A2(n_1082),
.B1(n_850),
.B2(n_1005),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_SL g1181 ( 
.A1(n_1127),
.A2(n_1017),
.B1(n_1008),
.B2(n_986),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1120),
.A2(n_1123),
.B1(n_1102),
.B2(n_1131),
.Y(n_1182)
);

AOI222xp33_ASAP7_75t_L g1183 ( 
.A1(n_1103),
.A2(n_959),
.B1(n_34),
.B2(n_35),
.C1(n_36),
.C2(n_37),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_L g1184 ( 
.A1(n_1136),
.A2(n_1000),
.B1(n_1005),
.B2(n_1004),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1125),
.A2(n_1000),
.B1(n_1005),
.B2(n_1004),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1117),
.A2(n_1140),
.B1(n_1141),
.B2(n_1139),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_SL g1187 ( 
.A1(n_1146),
.A2(n_1112),
.B1(n_1115),
.B2(n_1105),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1121),
.A2(n_1000),
.B1(n_1004),
.B2(n_877),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1135),
.A2(n_1004),
.B1(n_1008),
.B2(n_1017),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1113),
.B(n_1004),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1148),
.A2(n_1149),
.B1(n_1150),
.B2(n_1132),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1137),
.A2(n_1151),
.B1(n_1132),
.B2(n_1149),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1137),
.A2(n_1017),
.B1(n_1008),
.B2(n_539),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1152),
.A2(n_1017),
.B1(n_1008),
.B2(n_541),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1130),
.B(n_33),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_L g1196 ( 
.A1(n_1151),
.A2(n_541),
.B1(n_550),
.B2(n_538),
.Y(n_1196)
);

OAI222xp33_ASAP7_75t_L g1197 ( 
.A1(n_1093),
.A2(n_550),
.B1(n_37),
.B2(n_38),
.C1(n_39),
.C2(n_40),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1133),
.A2(n_538),
.B1(n_551),
.B2(n_552),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1130),
.A2(n_551),
.B1(n_552),
.B2(n_563),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_SL g1200 ( 
.A1(n_1134),
.A2(n_951),
.B1(n_38),
.B2(n_40),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1130),
.A2(n_563),
.B1(n_552),
.B2(n_551),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1130),
.A2(n_563),
.B1(n_552),
.B2(n_42),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_SL g1203 ( 
.A1(n_1134),
.A2(n_34),
.B1(n_41),
.B2(n_42),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1134),
.A2(n_563),
.B1(n_44),
.B2(n_45),
.Y(n_1204)
);

OAI222xp33_ASAP7_75t_L g1205 ( 
.A1(n_1128),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.C1(n_46),
.C2(n_47),
.Y(n_1205)
);

NAND3xp33_ASAP7_75t_SL g1206 ( 
.A(n_1128),
.B(n_46),
.C(n_47),
.Y(n_1206)
);

AOI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1134),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_1207)
);

HB1xp67_ASAP7_75t_L g1208 ( 
.A(n_1099),
.Y(n_1208)
);

OAI221xp5_ASAP7_75t_L g1209 ( 
.A1(n_1094),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.C(n_52),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1094),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1208),
.B(n_54),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1187),
.B(n_55),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1157),
.B(n_55),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1163),
.B(n_1167),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1172),
.B(n_56),
.Y(n_1215)
);

OAI211xp5_ASAP7_75t_L g1216 ( 
.A1(n_1183),
.A2(n_57),
.B(n_58),
.C(n_59),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_1176),
.B(n_86),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1172),
.B(n_57),
.Y(n_1218)
);

OA211x2_ASAP7_75t_L g1219 ( 
.A1(n_1206),
.A2(n_60),
.B(n_63),
.C(n_67),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1173),
.B(n_63),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_SL g1221 ( 
.A1(n_1207),
.A2(n_1210),
.B(n_1197),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1209),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_1176),
.B(n_1166),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1174),
.B(n_70),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1175),
.B(n_71),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1175),
.B(n_72),
.Y(n_1226)
);

NAND3xp33_ASAP7_75t_L g1227 ( 
.A(n_1207),
.B(n_73),
.C(n_94),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1155),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1173),
.B(n_98),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1179),
.A2(n_100),
.B1(n_101),
.B2(n_103),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_SL g1231 ( 
.A1(n_1158),
.A2(n_105),
.B(n_106),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1195),
.B(n_111),
.Y(n_1232)
);

NAND3xp33_ASAP7_75t_L g1233 ( 
.A(n_1203),
.B(n_112),
.C(n_115),
.Y(n_1233)
);

NOR3xp33_ASAP7_75t_L g1234 ( 
.A(n_1205),
.B(n_118),
.C(n_119),
.Y(n_1234)
);

OA21x2_ASAP7_75t_L g1235 ( 
.A1(n_1171),
.A2(n_121),
.B(n_125),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_SL g1236 ( 
.A1(n_1204),
.A2(n_130),
.B(n_132),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1182),
.B(n_134),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1195),
.B(n_135),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1191),
.B(n_136),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1192),
.B(n_341),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1186),
.B(n_139),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_1169),
.B(n_141),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1178),
.B(n_143),
.Y(n_1243)
);

OA21x2_ASAP7_75t_L g1244 ( 
.A1(n_1154),
.A2(n_144),
.B(n_146),
.Y(n_1244)
);

OAI21xp5_ASAP7_75t_SL g1245 ( 
.A1(n_1162),
.A2(n_1200),
.B(n_1202),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1170),
.B(n_148),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1190),
.B(n_150),
.Y(n_1247)
);

OAI221xp5_ASAP7_75t_SL g1248 ( 
.A1(n_1198),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.C(n_154),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1160),
.B(n_155),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1161),
.B(n_1168),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1159),
.B(n_156),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1153),
.B(n_158),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1170),
.B(n_159),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1185),
.B(n_340),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1181),
.B(n_160),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1180),
.A2(n_162),
.B1(n_164),
.B2(n_165),
.Y(n_1256)
);

OAI221xp5_ASAP7_75t_SL g1257 ( 
.A1(n_1196),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.C(n_174),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1214),
.B(n_1189),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1215),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1215),
.Y(n_1260)
);

NAND3xp33_ASAP7_75t_L g1261 ( 
.A(n_1227),
.B(n_1188),
.C(n_1194),
.Y(n_1261)
);

OAI211xp5_ASAP7_75t_SL g1262 ( 
.A1(n_1216),
.A2(n_1184),
.B(n_1164),
.C(n_1177),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1223),
.B(n_1165),
.Y(n_1263)
);

NAND3xp33_ASAP7_75t_L g1264 ( 
.A(n_1217),
.B(n_1193),
.C(n_1156),
.Y(n_1264)
);

AOI211xp5_ASAP7_75t_SL g1265 ( 
.A1(n_1248),
.A2(n_1201),
.B(n_1199),
.C(n_178),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1218),
.B(n_175),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1218),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1220),
.B(n_176),
.Y(n_1268)
);

OAI211xp5_ASAP7_75t_L g1269 ( 
.A1(n_1221),
.A2(n_179),
.B(n_181),
.C(n_182),
.Y(n_1269)
);

NAND4xp75_ASAP7_75t_L g1270 ( 
.A(n_1219),
.B(n_184),
.C(n_185),
.D(n_187),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1223),
.B(n_188),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1220),
.B(n_1213),
.Y(n_1272)
);

NOR2x1_ASAP7_75t_L g1273 ( 
.A(n_1211),
.B(n_189),
.Y(n_1273)
);

AOI211xp5_ASAP7_75t_L g1274 ( 
.A1(n_1217),
.A2(n_190),
.B(n_196),
.C(n_197),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1250),
.B(n_198),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1234),
.A2(n_200),
.B1(n_203),
.B2(n_205),
.Y(n_1276)
);

OR2x2_ASAP7_75t_L g1277 ( 
.A(n_1224),
.B(n_1225),
.Y(n_1277)
);

NAND3xp33_ASAP7_75t_L g1278 ( 
.A(n_1233),
.B(n_207),
.C(n_208),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1226),
.B(n_210),
.Y(n_1279)
);

NAND3xp33_ASAP7_75t_L g1280 ( 
.A(n_1228),
.B(n_212),
.C(n_213),
.Y(n_1280)
);

NAND4xp75_ASAP7_75t_L g1281 ( 
.A(n_1235),
.B(n_214),
.C(n_220),
.D(n_222),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1229),
.Y(n_1282)
);

NAND4xp75_ASAP7_75t_L g1283 ( 
.A(n_1235),
.B(n_223),
.C(n_225),
.D(n_226),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1250),
.B(n_230),
.Y(n_1284)
);

NOR3xp33_ASAP7_75t_L g1285 ( 
.A(n_1222),
.B(n_235),
.C(n_236),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1235),
.Y(n_1286)
);

XNOR2xp5_ASAP7_75t_L g1287 ( 
.A(n_1275),
.B(n_1212),
.Y(n_1287)
);

XNOR2xp5_ASAP7_75t_L g1288 ( 
.A(n_1275),
.B(n_1232),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1260),
.B(n_1244),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1282),
.B(n_1240),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1260),
.B(n_1232),
.Y(n_1291)
);

NAND4xp75_ASAP7_75t_SL g1292 ( 
.A(n_1263),
.B(n_1244),
.C(n_1255),
.D(n_1254),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_1259),
.B(n_1255),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1267),
.Y(n_1294)
);

AOI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1263),
.A2(n_1245),
.B1(n_1246),
.B2(n_1236),
.Y(n_1295)
);

NAND4xp75_ASAP7_75t_L g1296 ( 
.A(n_1271),
.B(n_1246),
.C(n_1242),
.D(n_1244),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1282),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1286),
.Y(n_1298)
);

INVx2_ASAP7_75t_SL g1299 ( 
.A(n_1277),
.Y(n_1299)
);

XNOR2xp5_ASAP7_75t_L g1300 ( 
.A(n_1284),
.B(n_1268),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1272),
.Y(n_1301)
);

NAND4xp75_ASAP7_75t_SL g1302 ( 
.A(n_1271),
.B(n_1251),
.C(n_1231),
.D(n_1257),
.Y(n_1302)
);

NAND4xp75_ASAP7_75t_L g1303 ( 
.A(n_1273),
.B(n_1242),
.C(n_1241),
.D(n_1238),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1258),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1258),
.B(n_1243),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1268),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1299),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1294),
.Y(n_1308)
);

INVxp67_ASAP7_75t_L g1309 ( 
.A(n_1299),
.Y(n_1309)
);

INVx1_ASAP7_75t_SL g1310 ( 
.A(n_1291),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1294),
.Y(n_1311)
);

XOR2x2_ASAP7_75t_L g1312 ( 
.A(n_1287),
.B(n_1270),
.Y(n_1312)
);

INVx2_ASAP7_75t_SL g1313 ( 
.A(n_1298),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1298),
.Y(n_1314)
);

OA22x2_ASAP7_75t_L g1315 ( 
.A1(n_1295),
.A2(n_1269),
.B1(n_1284),
.B2(n_1266),
.Y(n_1315)
);

INVxp33_ASAP7_75t_L g1316 ( 
.A(n_1287),
.Y(n_1316)
);

INVx1_ASAP7_75t_SL g1317 ( 
.A(n_1291),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1304),
.B(n_1281),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1316),
.A2(n_1296),
.B1(n_1264),
.B2(n_1303),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1308),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1311),
.Y(n_1321)
);

OA22x2_ASAP7_75t_L g1322 ( 
.A1(n_1318),
.A2(n_1300),
.B1(n_1288),
.B2(n_1309),
.Y(n_1322)
);

OA22x2_ASAP7_75t_L g1323 ( 
.A1(n_1318),
.A2(n_1293),
.B1(n_1301),
.B2(n_1305),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1316),
.A2(n_1305),
.B1(n_1276),
.B2(n_1293),
.Y(n_1324)
);

INVx2_ASAP7_75t_SL g1325 ( 
.A(n_1307),
.Y(n_1325)
);

OA22x2_ASAP7_75t_L g1326 ( 
.A1(n_1310),
.A2(n_1293),
.B1(n_1305),
.B2(n_1306),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1314),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1315),
.A2(n_1276),
.B1(n_1283),
.B2(n_1290),
.Y(n_1328)
);

OA22x2_ASAP7_75t_L g1329 ( 
.A1(n_1317),
.A2(n_1306),
.B1(n_1291),
.B2(n_1289),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1313),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1313),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1315),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1325),
.Y(n_1333)
);

INVxp67_ASAP7_75t_L g1334 ( 
.A(n_1322),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1320),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1331),
.Y(n_1336)
);

INVx1_ASAP7_75t_SL g1337 ( 
.A(n_1323),
.Y(n_1337)
);

INVxp67_ASAP7_75t_SL g1338 ( 
.A(n_1332),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1321),
.Y(n_1339)
);

INVxp67_ASAP7_75t_L g1340 ( 
.A(n_1332),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1327),
.Y(n_1341)
);

AOI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1334),
.A2(n_1319),
.B1(n_1328),
.B2(n_1312),
.Y(n_1342)
);

AOI221xp5_ASAP7_75t_L g1343 ( 
.A1(n_1338),
.A2(n_1324),
.B1(n_1330),
.B2(n_1285),
.C(n_1312),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1335),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1335),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1337),
.A2(n_1326),
.B1(n_1329),
.B2(n_1280),
.Y(n_1346)
);

OA22x2_ASAP7_75t_L g1347 ( 
.A1(n_1340),
.A2(n_1289),
.B1(n_1297),
.B2(n_1279),
.Y(n_1347)
);

AND4x1_ASAP7_75t_L g1348 ( 
.A(n_1342),
.B(n_1274),
.C(n_1265),
.D(n_1339),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1344),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1345),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1343),
.A2(n_1333),
.B1(n_1336),
.B2(n_1341),
.Y(n_1351)
);

AOI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1346),
.A2(n_1333),
.B1(n_1336),
.B2(n_1261),
.Y(n_1352)
);

AOI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1347),
.A2(n_1278),
.B1(n_1262),
.B2(n_1230),
.Y(n_1353)
);

NOR4xp25_ASAP7_75t_L g1354 ( 
.A(n_1351),
.B(n_1239),
.C(n_1237),
.D(n_1253),
.Y(n_1354)
);

OA22x2_ASAP7_75t_L g1355 ( 
.A1(n_1352),
.A2(n_1302),
.B1(n_1292),
.B2(n_1256),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1350),
.B(n_1251),
.Y(n_1356)
);

AO22x2_ASAP7_75t_L g1357 ( 
.A1(n_1349),
.A2(n_1252),
.B1(n_1249),
.B2(n_1247),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1353),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1348),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1350),
.Y(n_1360)
);

AOI211x1_ASAP7_75t_L g1361 ( 
.A1(n_1348),
.A2(n_238),
.B(n_239),
.C(n_241),
.Y(n_1361)
);

NOR2x1_ASAP7_75t_L g1362 ( 
.A(n_1360),
.B(n_1359),
.Y(n_1362)
);

OAI22x1_ASAP7_75t_L g1363 ( 
.A1(n_1358),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1356),
.Y(n_1364)
);

INVx2_ASAP7_75t_SL g1365 ( 
.A(n_1355),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1357),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1357),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1361),
.Y(n_1368)
);

AND4x1_ASAP7_75t_L g1369 ( 
.A(n_1362),
.B(n_1354),
.C(n_249),
.D(n_250),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1368),
.A2(n_246),
.B1(n_252),
.B2(n_254),
.Y(n_1370)
);

AOI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1365),
.A2(n_255),
.B1(n_256),
.B2(n_257),
.Y(n_1371)
);

NAND4xp25_ASAP7_75t_L g1372 ( 
.A(n_1367),
.B(n_258),
.C(n_259),
.D(n_261),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1364),
.Y(n_1373)
);

AOI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1363),
.A2(n_262),
.B1(n_263),
.B2(n_266),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1367),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1373),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1375),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1374),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1371),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1369),
.Y(n_1380)
);

INVx3_ASAP7_75t_L g1381 ( 
.A(n_1372),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1370),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1375),
.Y(n_1383)
);

AOI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1373),
.A2(n_1366),
.B1(n_269),
.B2(n_270),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1375),
.Y(n_1385)
);

AOI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1380),
.A2(n_268),
.B1(n_272),
.B2(n_273),
.Y(n_1386)
);

OAI22x1_ASAP7_75t_L g1387 ( 
.A1(n_1376),
.A2(n_274),
.B1(n_275),
.B2(n_276),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1385),
.Y(n_1388)
);

OAI22x1_ASAP7_75t_L g1389 ( 
.A1(n_1378),
.A2(n_281),
.B1(n_282),
.B2(n_284),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1377),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1385),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1383),
.Y(n_1392)
);

AO22x2_ASAP7_75t_SL g1393 ( 
.A1(n_1381),
.A2(n_291),
.B1(n_292),
.B2(n_296),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1381),
.Y(n_1394)
);

AOI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1382),
.A2(n_297),
.B1(n_298),
.B2(n_300),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1379),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1391),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1388),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1390),
.B(n_1384),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1396),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1392),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1394),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_SL g1403 ( 
.A1(n_1402),
.A2(n_1393),
.B1(n_1389),
.B2(n_1387),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1400),
.A2(n_1395),
.B1(n_1386),
.B2(n_308),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1399),
.A2(n_1397),
.B1(n_1401),
.B2(n_1398),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1405),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1403),
.Y(n_1407)
);

OAI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1406),
.A2(n_1404),
.B1(n_305),
.B2(n_310),
.Y(n_1408)
);

AO22x2_ASAP7_75t_L g1409 ( 
.A1(n_1407),
.A2(n_302),
.B1(n_311),
.B2(n_312),
.Y(n_1409)
);

AOI22xp5_ASAP7_75t_SL g1410 ( 
.A1(n_1406),
.A2(n_314),
.B1(n_316),
.B2(n_317),
.Y(n_1410)
);

INVxp67_ASAP7_75t_SL g1411 ( 
.A(n_1410),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1409),
.Y(n_1412)
);

AOI221x1_ASAP7_75t_L g1413 ( 
.A1(n_1412),
.A2(n_1408),
.B1(n_318),
.B2(n_326),
.C(n_330),
.Y(n_1413)
);

AOI211xp5_ASAP7_75t_L g1414 ( 
.A1(n_1413),
.A2(n_1411),
.B(n_331),
.C(n_334),
.Y(n_1414)
);


endmodule