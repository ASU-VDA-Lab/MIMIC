module fake_aes_1611_n_37 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_37);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_30;
wire n_16;
wire n_26;
wire n_13;
wire n_25;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g9 ( .A(n_0), .Y(n_9) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_2), .Y(n_10) );
BUFx10_ASAP7_75t_L g11 ( .A(n_6), .Y(n_11) );
NOR2xp33_ASAP7_75t_R g12 ( .A(n_8), .B(n_3), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_6), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_7), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_7), .Y(n_15) );
OR2x4_ASAP7_75t_L g16 ( .A(n_15), .B(n_0), .Y(n_16) );
AOI21xp5_ASAP7_75t_L g17 ( .A1(n_9), .A2(n_1), .B(n_2), .Y(n_17) );
OR2x6_ASAP7_75t_L g18 ( .A(n_11), .B(n_1), .Y(n_18) );
INVx1_ASAP7_75t_SL g19 ( .A(n_9), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_11), .B(n_3), .Y(n_20) );
AOI22xp5_ASAP7_75t_L g21 ( .A1(n_14), .A2(n_4), .B1(n_5), .B2(n_10), .Y(n_21) );
AND2x4_ASAP7_75t_L g22 ( .A(n_18), .B(n_13), .Y(n_22) );
NOR3xp33_ASAP7_75t_SL g23 ( .A(n_17), .B(n_11), .C(n_12), .Y(n_23) );
BUFx3_ASAP7_75t_L g24 ( .A(n_16), .Y(n_24) );
NOR2xp33_ASAP7_75t_R g25 ( .A(n_19), .B(n_4), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_22), .B(n_20), .Y(n_26) );
AND2x4_ASAP7_75t_L g27 ( .A(n_22), .B(n_18), .Y(n_27) );
OR2x2_ASAP7_75t_L g28 ( .A(n_22), .B(n_18), .Y(n_28) );
INVxp67_ASAP7_75t_SL g29 ( .A(n_27), .Y(n_29) );
OAI22xp33_ASAP7_75t_SL g30 ( .A1(n_28), .A2(n_21), .B1(n_22), .B2(n_24), .Y(n_30) );
AND2x2_ASAP7_75t_L g31 ( .A(n_29), .B(n_26), .Y(n_31) );
NAND4xp25_ASAP7_75t_L g32 ( .A(n_30), .B(n_21), .C(n_28), .D(n_24), .Y(n_32) );
OAI22xp5_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_27), .B1(n_26), .B2(n_23), .Y(n_33) );
BUFx6f_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
OR5x1_ASAP7_75t_L g35 ( .A(n_34), .B(n_5), .C(n_25), .D(n_23), .E(n_27), .Y(n_35) );
INVxp67_ASAP7_75t_L g36 ( .A(n_34), .Y(n_36) );
AOI22xp5_ASAP7_75t_L g37 ( .A1(n_36), .A2(n_24), .B1(n_33), .B2(n_35), .Y(n_37) );
endmodule