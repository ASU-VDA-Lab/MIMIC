module fake_jpeg_3627_n_573 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_573);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_573;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_6),
.B(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx8_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_53),
.Y(n_126)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g142 ( 
.A(n_54),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_17),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_55),
.B(n_76),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_18),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_58),
.B(n_63),
.Y(n_111)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_61),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_21),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_21),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_64),
.B(n_72),
.Y(n_112)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_65),
.Y(n_131)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g153 ( 
.A(n_67),
.Y(n_153)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_71),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_75),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_32),
.B(n_17),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_77),
.Y(n_152)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_78),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_79),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_40),
.B(n_18),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_95),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_81),
.Y(n_166)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_82),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_83),
.Y(n_167)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_84),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_85),
.Y(n_150)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_86),
.Y(n_158)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVxp67_ASAP7_75t_SL g134 ( 
.A(n_87),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_88),
.Y(n_151)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_89),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_35),
.Y(n_93)
);

INVx5_ASAP7_75t_SL g133 ( 
.A(n_93),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_19),
.B(n_18),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_94),
.B(n_16),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_42),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

BUFx12_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_97),
.Y(n_159)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

BUFx8_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_34),
.Y(n_103)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_104),
.Y(n_162)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

CKINVDCx9p33_ASAP7_75t_R g143 ( 
.A(n_105),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_49),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_106),
.B(n_41),
.Y(n_165)
);

HAxp5_ASAP7_75t_SL g109 ( 
.A(n_80),
.B(n_35),
.CON(n_109),
.SN(n_109)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_109),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_53),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_110),
.B(n_139),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_78),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_119),
.B(n_145),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_58),
.A2(n_41),
.B1(n_49),
.B2(n_52),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_120),
.A2(n_137),
.B1(n_69),
.B2(n_84),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_43),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_127),
.B(n_135),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_43),
.C(n_50),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_130),
.B(n_34),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_56),
.A2(n_52),
.B1(n_50),
.B2(n_48),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_61),
.A2(n_44),
.B(n_48),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_105),
.Y(n_145)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_74),
.Y(n_160)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_165),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_62),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_81),
.Y(n_192)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_75),
.Y(n_170)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_170),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_171),
.A2(n_198),
.B1(n_208),
.B2(n_216),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_126),
.A2(n_85),
.B1(n_88),
.B2(n_104),
.Y(n_172)
);

OAI22x1_ASAP7_75t_L g239 ( 
.A1(n_172),
.A2(n_210),
.B1(n_214),
.B2(n_159),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_163),
.Y(n_173)
);

BUFx2_ASAP7_75t_SL g259 ( 
.A(n_173),
.Y(n_259)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_174),
.Y(n_237)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_178),
.Y(n_255)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_180),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_126),
.Y(n_181)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_181),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_127),
.A2(n_100),
.B1(n_90),
.B2(n_77),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_182),
.A2(n_195),
.B1(n_167),
.B2(n_166),
.Y(n_240)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_115),
.Y(n_183)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_183),
.Y(n_246)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_115),
.Y(n_184)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_184),
.Y(n_241)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_116),
.Y(n_185)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_185),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_44),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_186),
.B(n_194),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_112),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_188),
.B(n_201),
.Y(n_236)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_150),
.Y(n_189)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_189),
.Y(n_285)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_190),
.Y(n_235)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_118),
.Y(n_191)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_191),
.Y(n_276)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_192),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_193),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_111),
.B(n_117),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_107),
.A2(n_83),
.B1(n_52),
.B2(n_60),
.Y(n_195)
);

INVx11_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_197),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_137),
.A2(n_49),
.B1(n_45),
.B2(n_38),
.Y(n_198)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_113),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_199),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_113),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_200),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_123),
.B(n_26),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_131),
.B(n_26),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_202),
.B(n_203),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_122),
.B(n_23),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_144),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_204),
.Y(n_269)
);

AO22x1_ASAP7_75t_SL g205 ( 
.A1(n_138),
.A2(n_85),
.B1(n_88),
.B2(n_91),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_219),
.Y(n_238)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_121),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_206),
.Y(n_271)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_132),
.Y(n_207)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_207),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_128),
.A2(n_19),
.B1(n_23),
.B2(n_30),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_148),
.Y(n_209)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_209),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_143),
.A2(n_101),
.B1(n_86),
.B2(n_82),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_163),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_211),
.B(n_213),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_142),
.B(n_73),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_147),
.A2(n_34),
.B1(n_46),
.B2(n_45),
.Y(n_214)
);

CKINVDCx9p33_ASAP7_75t_R g215 ( 
.A(n_129),
.Y(n_215)
);

INVx13_ASAP7_75t_L g280 ( 
.A(n_215),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_154),
.A2(n_36),
.B1(n_46),
.B2(n_31),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_132),
.Y(n_217)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_217),
.Y(n_260)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_121),
.Y(n_218)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_218),
.Y(n_263)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_162),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_220),
.Y(n_274)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_162),
.Y(n_221)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_221),
.Y(n_275)
);

BUFx12f_ASAP7_75t_L g222 ( 
.A(n_129),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_222),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_141),
.Y(n_223)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_156),
.Y(n_225)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_225),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_142),
.B(n_38),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_230),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_141),
.Y(n_227)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_227),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_129),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_228),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_136),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_154),
.A2(n_128),
.B1(n_149),
.B2(n_109),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_231),
.A2(n_108),
.B1(n_97),
.B2(n_152),
.Y(n_286)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_134),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_133),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_134),
.B(n_158),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_233),
.B(n_164),
.Y(n_268)
);

BUFx24_ASAP7_75t_SL g234 ( 
.A(n_212),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_234),
.B(n_267),
.Y(n_289)
);

INVxp67_ASAP7_75t_SL g292 ( 
.A(n_239),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_240),
.A2(n_261),
.B1(n_215),
.B2(n_238),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_140),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_250),
.B(n_266),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_216),
.A2(n_31),
.B1(n_30),
.B2(n_36),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_251),
.A2(n_214),
.B1(n_195),
.B2(n_172),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_177),
.A2(n_124),
.B1(n_136),
.B2(n_164),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_253),
.B(n_228),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_175),
.B(n_147),
.C(n_108),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_257),
.B(n_238),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_182),
.A2(n_149),
.B1(n_166),
.B2(n_167),
.Y(n_261)
);

AO22x2_ASAP7_75t_L g296 ( 
.A1(n_261),
.A2(n_205),
.B1(n_217),
.B2(n_207),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_262),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_179),
.B(n_146),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_196),
.B(n_133),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_268),
.B(n_286),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_187),
.B(n_146),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_282),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_229),
.A2(n_159),
.B(n_97),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_281),
.A2(n_35),
.B(n_222),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_233),
.Y(n_282)
);

FAx1_ASAP7_75t_SL g284 ( 
.A(n_229),
.B(n_153),
.CI(n_125),
.CON(n_284),
.SN(n_284)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_284),
.B(n_181),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_288),
.A2(n_290),
.B1(n_304),
.B2(n_315),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_294),
.B(n_299),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_269),
.Y(n_295)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_295),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_296),
.B(n_303),
.Y(n_381)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_241),
.Y(n_297)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_297),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_249),
.A2(n_152),
.B1(n_210),
.B2(n_206),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_298),
.A2(n_273),
.B1(n_237),
.B2(n_259),
.Y(n_339)
);

AND2x6_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_205),
.Y(n_299)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_246),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_300),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_245),
.B(n_176),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_301),
.B(n_308),
.Y(n_357)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_246),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_302),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_238),
.A2(n_199),
.B1(n_218),
.B2(n_223),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_274),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_305),
.B(n_317),
.Y(n_347)
);

MAJx2_ASAP7_75t_L g306 ( 
.A(n_250),
.B(n_224),
.C(n_197),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_306),
.B(n_270),
.C(n_264),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_281),
.A2(n_221),
.B(n_220),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_SL g362 ( 
.A(n_307),
.B(n_329),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_258),
.B(n_244),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_268),
.Y(n_309)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_309),
.Y(n_340)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_275),
.Y(n_310)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_310),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_311),
.B(n_0),
.Y(n_356)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_283),
.Y(n_313)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_313),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_249),
.A2(n_227),
.B1(n_200),
.B2(n_184),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_266),
.B(n_183),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_316),
.Y(n_351)
);

A2O1A1Ixp33_ASAP7_75t_L g317 ( 
.A1(n_279),
.A2(n_35),
.B(n_222),
.C(n_125),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_284),
.B(n_190),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_318),
.B(n_319),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_236),
.B(n_189),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_320),
.A2(n_336),
.B(n_8),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_278),
.B(n_257),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_321),
.B(n_323),
.Y(n_372)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_241),
.Y(n_322)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_322),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_254),
.B(n_125),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_287),
.Y(n_324)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_324),
.Y(n_374)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_255),
.Y(n_325)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_325),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_274),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_326),
.B(n_328),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_285),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_327),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_285),
.B(n_174),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_255),
.B(n_193),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_263),
.B(n_34),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_330),
.B(n_5),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_248),
.B(n_17),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_331),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_240),
.A2(n_235),
.B1(n_239),
.B2(n_252),
.Y(n_332)
);

OAI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_332),
.A2(n_337),
.B1(n_252),
.B2(n_280),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_260),
.B(n_16),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_333),
.Y(n_370)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_243),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_334),
.Y(n_363)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_256),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_335),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_286),
.A2(n_35),
.B(n_39),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_235),
.A2(n_39),
.B1(n_1),
.B2(n_2),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g402 ( 
.A1(n_338),
.A2(n_378),
.B1(n_290),
.B2(n_341),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_339),
.A2(n_348),
.B1(n_350),
.B2(n_354),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_315),
.A2(n_243),
.B1(n_271),
.B2(n_265),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_343),
.A2(n_345),
.B1(n_346),
.B2(n_365),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_292),
.A2(n_271),
.B1(n_265),
.B2(n_237),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_298),
.A2(n_273),
.B1(n_276),
.B2(n_272),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_314),
.A2(n_242),
.B1(n_276),
.B2(n_272),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_314),
.A2(n_242),
.B1(n_256),
.B2(n_247),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_318),
.A2(n_264),
.B1(n_280),
.B2(n_270),
.Y(n_354)
);

NAND3xp33_ASAP7_75t_L g404 ( 
.A(n_355),
.B(n_323),
.C(n_329),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_356),
.B(n_358),
.C(n_309),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_311),
.B(n_1),
.C(n_2),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_312),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_359),
.A2(n_368),
.B1(n_371),
.B2(n_379),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_312),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_365)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_367),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_312),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_369),
.B(n_320),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_299),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_375),
.B(n_317),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_319),
.A2(n_291),
.B1(n_293),
.B2(n_321),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_304),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_344),
.Y(n_382)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_382),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_383),
.B(n_398),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_364),
.B(n_294),
.Y(n_384)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_384),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_385),
.A2(n_371),
.B1(n_359),
.B2(n_354),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_344),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_386),
.Y(n_440)
);

O2A1O1Ixp33_ASAP7_75t_L g389 ( 
.A1(n_347),
.A2(n_375),
.B(n_364),
.C(n_362),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_389),
.B(n_393),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_362),
.B(n_307),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_391),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_357),
.B(n_295),
.Y(n_392)
);

NAND3xp33_ASAP7_75t_L g434 ( 
.A(n_392),
.B(n_395),
.C(n_397),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_351),
.B(n_305),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_351),
.B(n_326),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_394),
.B(n_399),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_366),
.B(n_291),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_366),
.B(n_370),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_347),
.A2(n_303),
.B(n_336),
.Y(n_399)
);

CKINVDCx14_ASAP7_75t_R g400 ( 
.A(n_372),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_400),
.B(n_411),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g401 ( 
.A(n_340),
.B(n_306),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_401),
.B(n_406),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_402),
.A2(n_404),
.B1(n_408),
.B2(n_416),
.Y(n_425)
);

AND2x2_ASAP7_75t_SL g403 ( 
.A(n_340),
.B(n_328),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_403),
.B(n_381),
.Y(n_420)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_380),
.Y(n_405)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_405),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_380),
.B(n_330),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_349),
.Y(n_407)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_407),
.Y(n_441)
);

INVx11_ASAP7_75t_L g408 ( 
.A(n_376),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_372),
.B(n_313),
.C(n_310),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_409),
.B(n_377),
.C(n_352),
.Y(n_427)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_360),
.Y(n_410)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_410),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_370),
.B(n_289),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_350),
.Y(n_412)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_412),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_361),
.B(n_324),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_413),
.B(n_414),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_348),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_353),
.A2(n_296),
.B(n_327),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_415),
.B(n_417),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_381),
.A2(n_296),
.B1(n_324),
.B2(n_334),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_342),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_361),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_418),
.B(n_360),
.Y(n_436)
);

AO21x1_ASAP7_75t_L g469 ( 
.A1(n_420),
.A2(n_428),
.B(n_439),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_412),
.A2(n_405),
.B1(n_416),
.B2(n_414),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_423),
.A2(n_430),
.B1(n_431),
.B2(n_442),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_384),
.A2(n_381),
.B1(n_346),
.B2(n_339),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_424),
.A2(n_388),
.B1(n_396),
.B2(n_374),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_393),
.B(n_356),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_426),
.B(n_449),
.C(n_388),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_427),
.B(n_444),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_394),
.A2(n_390),
.B1(n_391),
.B2(n_418),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_390),
.A2(n_391),
.B1(n_399),
.B2(n_384),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g472 ( 
.A(n_436),
.Y(n_472)
);

XOR2x2_ASAP7_75t_L g437 ( 
.A(n_409),
.B(n_355),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_437),
.B(n_446),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_385),
.A2(n_374),
.B1(n_376),
.B2(n_363),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_406),
.A2(n_343),
.B1(n_345),
.B2(n_352),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_398),
.B(n_383),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_403),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_401),
.B(n_358),
.C(n_377),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_389),
.B(n_369),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_450),
.B(n_368),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_430),
.B(n_413),
.Y(n_452)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_452),
.Y(n_486)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_438),
.Y(n_455)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_455),
.Y(n_501)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_438),
.Y(n_456)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_456),
.Y(n_504)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_447),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_L g497 ( 
.A1(n_457),
.A2(n_458),
.B1(n_463),
.B2(n_476),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_434),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_419),
.A2(n_415),
.B(n_401),
.Y(n_459)
);

AO21x1_ASAP7_75t_L g483 ( 
.A1(n_459),
.A2(n_460),
.B(n_462),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_419),
.A2(n_385),
.B(n_387),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_451),
.B(n_403),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_461),
.B(n_420),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_443),
.A2(n_387),
.B(n_417),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_433),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_427),
.B(n_392),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_464),
.B(n_465),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_435),
.B(n_407),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_443),
.A2(n_403),
.B(n_410),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_466),
.A2(n_445),
.B(n_451),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_467),
.B(n_471),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_468),
.A2(n_474),
.B1(n_478),
.B2(n_479),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_421),
.A2(n_365),
.B(n_396),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_473),
.A2(n_477),
.B(n_429),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_424),
.A2(n_386),
.B1(n_382),
.B2(n_373),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_423),
.A2(n_379),
.B1(n_386),
.B2(n_382),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_475),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_440),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_421),
.A2(n_373),
.B(n_325),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_448),
.A2(n_296),
.B1(n_349),
.B2(n_322),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_425),
.A2(n_302),
.B1(n_297),
.B2(n_300),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g480 ( 
.A(n_429),
.Y(n_480)
);

INVx13_ASAP7_75t_L g496 ( 
.A(n_480),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_453),
.B(n_437),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_SL g512 ( 
.A(n_482),
.B(n_488),
.Y(n_512)
);

AO21x1_ASAP7_75t_L g515 ( 
.A1(n_484),
.A2(n_491),
.B(n_469),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_453),
.B(n_444),
.C(n_432),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_487),
.B(n_499),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_471),
.B(n_431),
.Y(n_488)
);

XOR2x2_ASAP7_75t_L g489 ( 
.A(n_459),
.B(n_450),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g505 ( 
.A(n_489),
.Y(n_505)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_490),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_452),
.B(n_440),
.Y(n_492)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_492),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_454),
.B(n_426),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_495),
.B(n_487),
.C(n_482),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_472),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_498),
.B(n_470),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_467),
.B(n_449),
.C(n_439),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_477),
.B(n_441),
.C(n_428),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_500),
.B(n_460),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_469),
.B(n_442),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_502),
.B(n_474),
.C(n_479),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_476),
.B(n_422),
.Y(n_503)
);

OAI321xp33_ASAP7_75t_L g510 ( 
.A1(n_503),
.A2(n_466),
.A3(n_461),
.B1(n_463),
.B2(n_457),
.C(n_462),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_493),
.A2(n_456),
.B1(n_455),
.B2(n_468),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_506),
.A2(n_510),
.B1(n_516),
.B2(n_484),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_485),
.B(n_458),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_509),
.B(n_519),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_481),
.A2(n_470),
.B1(n_473),
.B2(n_475),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_511),
.A2(n_521),
.B1(n_497),
.B2(n_504),
.Y(n_525)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_513),
.Y(n_524)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_514),
.Y(n_527)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_515),
.Y(n_532)
);

CKINVDCx14_ASAP7_75t_R g516 ( 
.A(n_500),
.Y(n_516)
);

MAJx2_ASAP7_75t_L g528 ( 
.A(n_518),
.B(n_499),
.C(n_502),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_488),
.B(n_478),
.C(n_422),
.Y(n_519)
);

OA22x2_ASAP7_75t_L g520 ( 
.A1(n_504),
.A2(n_296),
.B1(n_408),
.B2(n_335),
.Y(n_520)
);

OAI21xp33_ASAP7_75t_SL g531 ( 
.A1(n_520),
.A2(n_503),
.B(n_492),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_SL g521 ( 
.A1(n_481),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_494),
.B(n_14),
.C(n_15),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_522),
.B(n_491),
.C(n_501),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_523),
.B(n_495),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_525),
.B(n_528),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_526),
.B(n_529),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_530),
.B(n_531),
.Y(n_549)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_514),
.Y(n_533)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_533),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_505),
.A2(n_483),
.B(n_494),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_534),
.B(n_535),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_508),
.B(n_489),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g537 ( 
.A(n_505),
.B(n_490),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_537),
.B(n_538),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_519),
.B(n_512),
.C(n_523),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_515),
.B(n_483),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_539),
.B(n_517),
.Y(n_548)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_536),
.Y(n_542)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_542),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_538),
.B(n_512),
.C(n_511),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_543),
.B(n_544),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_526),
.B(n_506),
.C(n_518),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_535),
.B(n_507),
.Y(n_545)
);

CKINVDCx16_ASAP7_75t_R g555 ( 
.A(n_545),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_548),
.B(n_528),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_SL g550 ( 
.A(n_524),
.B(n_529),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_550),
.A2(n_539),
.B1(n_522),
.B2(n_496),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_549),
.A2(n_532),
.B1(n_527),
.B2(n_486),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_552),
.B(n_553),
.Y(n_563)
);

INVx6_ASAP7_75t_L g553 ( 
.A(n_551),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_554),
.B(n_556),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_L g559 ( 
.A1(n_549),
.A2(n_531),
.B(n_496),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_559),
.B(n_557),
.C(n_540),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_SL g565 ( 
.A1(n_560),
.A2(n_559),
.B(n_541),
.Y(n_565)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_558),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_L g566 ( 
.A1(n_561),
.A2(n_555),
.B(n_547),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_562),
.A2(n_553),
.B(n_556),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_564),
.B(n_546),
.Y(n_568)
);

AO21x2_ASAP7_75t_L g567 ( 
.A1(n_565),
.A2(n_566),
.B(n_552),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_567),
.B(n_568),
.C(n_563),
.Y(n_569)
);

AOI322xp5_ASAP7_75t_L g570 ( 
.A1(n_569),
.A2(n_520),
.A3(n_543),
.B1(n_544),
.B2(n_546),
.C1(n_563),
.C2(n_568),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_570),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_571),
.B(n_520),
.Y(n_572)
);

BUFx24_ASAP7_75t_SL g573 ( 
.A(n_572),
.Y(n_573)
);


endmodule