module real_jpeg_2946_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_150;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_1),
.A2(n_35),
.B1(n_37),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_52),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_1),
.A2(n_48),
.B1(n_50),
.B2(n_52),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_1),
.A2(n_52),
.B1(n_62),
.B2(n_64),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_2),
.A2(n_48),
.B1(n_50),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_2),
.A2(n_62),
.B1(n_64),
.B2(n_69),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_3),
.A2(n_62),
.B1(n_64),
.B2(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_3),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_4),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_5),
.A2(n_35),
.B1(n_37),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_5),
.A2(n_54),
.B1(n_62),
.B2(n_64),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_5),
.A2(n_48),
.B1(n_50),
.B2(n_54),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_6),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_6),
.A2(n_39),
.B1(n_48),
.B2(n_50),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_6),
.A2(n_39),
.B1(n_62),
.B2(n_64),
.Y(n_152)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_10),
.A2(n_25),
.B(n_27),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_10),
.B(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_10),
.B(n_59),
.C(n_62),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_10),
.A2(n_29),
.B1(n_48),
.B2(n_50),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_10),
.B(n_76),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_10),
.B(n_70),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_10),
.B(n_37),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_10),
.A2(n_37),
.B(n_172),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_12),
.A2(n_48),
.B1(n_50),
.B2(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_12),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_12),
.A2(n_35),
.B1(n_37),
.B2(n_66),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_12),
.A2(n_62),
.B1(n_64),
.B2(n_66),
.Y(n_133)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_14),
.A2(n_62),
.B1(n_64),
.B2(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_14),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_14),
.A2(n_48),
.B1(n_50),
.B2(n_79),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_124),
.B1(n_200),
.B2(n_201),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_18),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_122),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_98),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_20),
.B(n_98),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_71),
.C(n_85),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_21),
.A2(n_22),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_23),
.B(n_41),
.C(n_55),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B1(n_34),
.B2(n_38),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_29),
.Y(n_28)
);

NAND3xp33_ASAP7_75t_L g84 ( 
.A(n_26),
.B(n_33),
.C(n_37),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_28),
.A2(n_32),
.B(n_35),
.C(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_29),
.B(n_47),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_29),
.A2(n_74),
.B1(n_76),
.B2(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_30),
.A2(n_34),
.B1(n_38),
.B2(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_32),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_33),
.B1(n_35),
.B2(n_37),
.Y(n_34)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

CKINVDCx6p67_ASAP7_75t_R g37 ( 
.A(n_35),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_37),
.B1(n_44),
.B2(n_46),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI32xp33_ASAP7_75t_L g170 ( 
.A1(n_37),
.A2(n_44),
.A3(n_48),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_55),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_47),
.B1(n_51),
.B2(n_53),
.Y(n_41)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_42),
.A2(n_53),
.B(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_42),
.A2(n_47),
.B1(n_88),
.B2(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_47),
.Y(n_42)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

OA22x2_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_47)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_46),
.B(n_50),
.Y(n_173)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

CKINVDCx6p67_ASAP7_75t_R g50 ( 
.A(n_48),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_50),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_48),
.B(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_65),
.B(n_67),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_56),
.A2(n_61),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_57),
.B(n_68),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_57),
.A2(n_70),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_57),
.A2(n_70),
.B1(n_137),
.B2(n_145),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_57),
.A2(n_186),
.B(n_187),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_64),
.Y(n_61)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_61),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_61),
.B(n_65),
.Y(n_187)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_62),
.B(n_150),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_71),
.B(n_85),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_82),
.B2(n_83),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_82),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_76),
.B1(n_77),
.B2(n_80),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_74),
.B(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_74),
.A2(n_131),
.B(n_132),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_74),
.A2(n_76),
.B1(n_152),
.B2(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_78),
.B(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_75),
.B(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_75),
.A2(n_116),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_76),
.B(n_97),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_80),
.Y(n_117)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_92),
.C(n_94),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_86),
.B(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_90),
.B(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_92),
.A2(n_94),
.B1(n_95),
.B2(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_92),
.Y(n_191)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_109),
.B2(n_110),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_119),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B(n_118),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_116),
.A2(n_118),
.B(n_133),
.Y(n_174)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_124),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_194),
.B(n_199),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_182),
.B(n_193),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_165),
.B(n_181),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_146),
.B(n_164),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_139),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_139),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_134),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_136),
.C(n_167),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_131),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_140),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_158),
.B(n_163),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_153),
.B(n_157),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_156),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_155),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_162),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_168),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_175),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_176),
.C(n_179),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_174),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_174),
.Y(n_188)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_178),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_192),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_192),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_189),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_188),
.C(n_189),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_196),
.Y(n_199)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);


endmodule