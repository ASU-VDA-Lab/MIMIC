module fake_aes_207_n_16 (n_1, n_2, n_0, n_16);
input n_1;
input n_2;
input n_0;
output n_16;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
INVx1_ASAP7_75t_SL g3 ( .A(n_1), .Y(n_3) );
INVx2_ASAP7_75t_L g4 ( .A(n_0), .Y(n_4) );
AOI21x1_ASAP7_75t_L g5 ( .A1(n_4), .A2(n_0), .B(n_1), .Y(n_5) );
BUFx6f_ASAP7_75t_L g6 ( .A(n_4), .Y(n_6) );
AND2x2_ASAP7_75t_L g7 ( .A(n_6), .B(n_3), .Y(n_7) );
INVx2_ASAP7_75t_L g8 ( .A(n_6), .Y(n_8) );
OAI211xp5_ASAP7_75t_L g9 ( .A1(n_7), .A2(n_5), .B(n_6), .C(n_0), .Y(n_9) );
OR2x2_ASAP7_75t_L g10 ( .A(n_8), .B(n_1), .Y(n_10) );
NAND2xp5_ASAP7_75t_L g11 ( .A(n_9), .B(n_0), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_10), .B(n_0), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_12), .B(n_1), .Y(n_13) );
OAI211xp5_ASAP7_75t_SL g14 ( .A1(n_11), .A2(n_8), .B(n_2), .C(n_6), .Y(n_14) );
OAI22xp5_ASAP7_75t_L g15 ( .A1(n_13), .A2(n_2), .B1(n_6), .B2(n_14), .Y(n_15) );
OAI21xp5_ASAP7_75t_L g16 ( .A1(n_15), .A2(n_2), .B(n_13), .Y(n_16) );
endmodule