module fake_jpeg_8614_n_134 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_134);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_134;

wire n_117;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx2_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_12),
.B(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_19),
.Y(n_27)
);

NAND3xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_29),
.C(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_30),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_32),
.A2(n_39),
.B1(n_40),
.B2(n_17),
.Y(n_51)
);

OR2x6_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_10),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_22),
.B(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_38),
.B(n_4),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_27),
.A2(n_15),
.B1(n_18),
.B2(n_20),
.Y(n_39)
);

OA22x2_ASAP7_75t_L g40 ( 
.A1(n_26),
.A2(n_16),
.B1(n_20),
.B2(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_42),
.Y(n_65)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_36),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_48),
.Y(n_60)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_44),
.B(n_50),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_47),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_23),
.C(n_19),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_56),
.B(n_11),
.Y(n_76)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_25),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_17),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_49),
.B(n_54),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_31),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_51),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_52),
.A2(n_30),
.B(n_28),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_53),
.B(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_24),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_1),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_30),
.C(n_28),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_6),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_1),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_58),
.B(n_3),
.Y(n_75)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_59),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_71),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_16),
.B(n_3),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_21),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_26),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_67),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_21),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_46),
.B(n_4),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_72),
.Y(n_79)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_74),
.Y(n_80)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_76),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_53),
.B1(n_51),
.B2(n_59),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_78),
.Y(n_94)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_81),
.B(n_86),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_45),
.C(n_52),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_90),
.C(n_76),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_83),
.Y(n_95)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_84),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_77),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_87),
.B(n_91),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_88),
.B(n_62),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_57),
.C(n_41),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_62),
.A2(n_47),
.B1(n_42),
.B2(n_11),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_61),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_82),
.C(n_79),
.Y(n_106)
);

NOR3xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_66),
.C(n_69),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_99),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_84),
.B(n_60),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_103),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_89),
.B(n_64),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_106),
.Y(n_112)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_109),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_89),
.C(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_111),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_115),
.Y(n_122)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_113),
.A2(n_97),
.B(n_109),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_119),
.C(n_112),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_117),
.A2(n_106),
.B(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_100),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_124),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_102),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_SL g129 ( 
.A1(n_126),
.A2(n_99),
.B(n_94),
.C(n_63),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_73),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_127),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_129),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_125),
.Y(n_132)
);

OAI32xp33_ASAP7_75t_SL g133 ( 
.A1(n_132),
.A2(n_130),
.A3(n_126),
.B1(n_92),
.B2(n_9),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_131),
.Y(n_134)
);


endmodule