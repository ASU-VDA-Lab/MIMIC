module fake_netlist_1_9859_n_21 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_21);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_21;
wire n_20;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_19;
NAND2xp5_ASAP7_75t_SL g11 ( .A(n_8), .B(n_7), .Y(n_11) );
INVx6_ASAP7_75t_L g12 ( .A(n_7), .Y(n_12) );
NAND2xp5_ASAP7_75t_SL g13 ( .A(n_4), .B(n_10), .Y(n_13) );
AND2x6_ASAP7_75t_L g14 ( .A(n_5), .B(n_6), .Y(n_14) );
INVx4_ASAP7_75t_L g15 ( .A(n_2), .Y(n_15) );
OAI21x1_ASAP7_75t_L g16 ( .A1(n_11), .A2(n_9), .B(n_1), .Y(n_16) );
OAI211xp5_ASAP7_75t_SL g17 ( .A1(n_16), .A2(n_13), .B(n_15), .C(n_12), .Y(n_17) );
AOI22xp5_ASAP7_75t_L g18 ( .A1(n_17), .A2(n_14), .B1(n_12), .B2(n_16), .Y(n_18) );
AOI222xp33_ASAP7_75t_L g19 ( .A1(n_18), .A2(n_14), .B1(n_1), .B2(n_2), .C1(n_3), .C2(n_0), .Y(n_19) );
OAI22xp5_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_14), .B1(n_3), .B2(n_4), .Y(n_20) );
AOI22xp33_ASAP7_75t_SL g21 ( .A1(n_20), .A2(n_0), .B1(n_5), .B2(n_6), .Y(n_21) );
endmodule