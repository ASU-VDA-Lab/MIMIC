module real_jpeg_3679_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_38;
wire n_35;
wire n_33;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_23;
wire n_11;
wire n_14;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_0),
.B(n_9),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_0),
.B(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_0),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_0),
.B(n_36),
.Y(n_44)
);

OR2x4_ASAP7_75t_L g17 ( 
.A(n_1),
.B(n_18),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_1),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_1),
.B(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_2),
.A2(n_37),
.B(n_38),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_3),
.B(n_5),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_3),
.B(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_4),
.B(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_5),
.B(n_12),
.Y(n_11)
);

NAND2x1_ASAP7_75t_SL g13 ( 
.A(n_5),
.B(n_12),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_5),
.B(n_21),
.Y(n_20)
);

AOI221xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_16),
.B1(n_19),
.B2(n_24),
.C(n_27),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_14),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_9),
.B(n_21),
.Y(n_23)
);

OA21x2_ASAP7_75t_L g9 ( 
.A1(n_10),
.A2(n_11),
.B(n_13),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_10),
.B(n_21),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_10),
.B(n_21),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_17),
.Y(n_16)
);

AND2x2_ASAP7_75t_SL g29 ( 
.A(n_18),
.B(n_26),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_22),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_30),
.B1(n_39),
.B2(n_42),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);


endmodule