module fake_netlist_1_532_n_20 (n_1, n_2, n_0, n_20);
input n_1;
input n_2;
input n_0;
output n_20;
wire n_5;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_3;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_6;
wire n_4;
wire n_7;
NOR2xp33_ASAP7_75t_R g3 ( .A(n_0), .B(n_2), .Y(n_3) );
CKINVDCx5p33_ASAP7_75t_R g4 ( .A(n_2), .Y(n_4) );
BUFx3_ASAP7_75t_L g5 ( .A(n_0), .Y(n_5) );
A2O1A1Ixp33_ASAP7_75t_L g6 ( .A1(n_5), .A2(n_0), .B(n_1), .C(n_2), .Y(n_6) );
AOI21xp5_ASAP7_75t_L g7 ( .A1(n_5), .A2(n_0), .B(n_1), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_5), .B(n_0), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
INVxp67_ASAP7_75t_L g10 ( .A(n_8), .Y(n_10) );
AND2x2_ASAP7_75t_L g11 ( .A(n_10), .B(n_4), .Y(n_11) );
INVx6_ASAP7_75t_L g12 ( .A(n_9), .Y(n_12) );
AOI322xp5_ASAP7_75t_SL g13 ( .A1(n_11), .A2(n_3), .A3(n_2), .B1(n_6), .B2(n_1), .C1(n_4), .C2(n_9), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_12), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_14), .Y(n_15) );
AOI211xp5_ASAP7_75t_L g16 ( .A1(n_13), .A2(n_7), .B(n_3), .C(n_5), .Y(n_16) );
AO22x1_ASAP7_75t_L g17 ( .A1(n_15), .A2(n_13), .B1(n_14), .B2(n_1), .Y(n_17) );
NOR2xp33_ASAP7_75t_L g18 ( .A(n_15), .B(n_12), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_17), .Y(n_19) );
AOI222xp33_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_1), .B1(n_12), .B2(n_16), .C1(n_18), .C2(n_17), .Y(n_20) );
endmodule