module fake_jpeg_2405_n_444 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_444);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_444;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_15),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_5),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_54),
.Y(n_127)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_57),
.Y(n_136)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_58),
.Y(n_142)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_60),
.Y(n_148)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_17),
.B(n_12),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_62),
.B(n_88),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_63),
.Y(n_144)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_64),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_34),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_65),
.B(n_75),
.Y(n_139)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_67),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_68),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_69),
.Y(n_175)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_70),
.Y(n_181)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_71),
.Y(n_183)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_72),
.Y(n_156)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_73),
.Y(n_180)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_74),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_77),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_78),
.Y(n_137)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_26),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_79),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_42),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_80),
.B(n_86),
.Y(n_149)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_81),
.Y(n_140)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_83),
.Y(n_165)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_84),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_85),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_30),
.B(n_12),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_87),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_19),
.B(n_16),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_42),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_90),
.B(n_92),
.Y(n_159)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_42),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_47),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_93),
.B(n_101),
.Y(n_164)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_19),
.B(n_0),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_95),
.B(n_97),
.Y(n_160)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

AO22x1_ASAP7_75t_L g141 ( 
.A1(n_96),
.A2(n_103),
.B1(n_107),
.B2(n_110),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_20),
.B(n_0),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_98),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_99),
.Y(n_122)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_100),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_32),
.Y(n_101)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_31),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_102),
.B(n_104),
.Y(n_168)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_32),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_105),
.B(n_106),
.Y(n_178)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_22),
.Y(n_106)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_30),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_30),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_108),
.B(n_111),
.Y(n_166)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_24),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_109),
.B(n_112),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g110 ( 
.A(n_31),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_20),
.B(n_0),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_51),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_51),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_113),
.B(n_18),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_86),
.A2(n_29),
.B1(n_33),
.B2(n_24),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_114),
.A2(n_160),
.B(n_166),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_63),
.A2(n_29),
.B1(n_33),
.B2(n_28),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_116),
.A2(n_123),
.B1(n_125),
.B2(n_143),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_79),
.A2(n_31),
.B1(n_46),
.B2(n_44),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g239 ( 
.A1(n_117),
.A2(n_120),
.B1(n_135),
.B2(n_152),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_60),
.A2(n_35),
.B1(n_46),
.B2(n_44),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_76),
.A2(n_41),
.B1(n_38),
.B2(n_36),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_54),
.B(n_41),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_124),
.B(n_146),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_68),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_69),
.A2(n_18),
.B1(n_49),
.B2(n_40),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_128),
.A2(n_131),
.B1(n_173),
.B2(n_141),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_129),
.B(n_139),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_104),
.A2(n_49),
.B1(n_40),
.B2(n_39),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_59),
.A2(n_50),
.B1(n_39),
.B2(n_37),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_78),
.A2(n_50),
.B1(n_37),
.B2(n_25),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_55),
.A2(n_25),
.B1(n_23),
.B2(n_4),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_150),
.A2(n_151),
.B1(n_153),
.B2(n_154),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_87),
.A2(n_23),
.B1(n_2),
.B2(n_5),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_64),
.A2(n_1),
.B1(n_2),
.B2(n_7),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_71),
.A2(n_1),
.B1(n_7),
.B2(n_8),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_74),
.A2(n_1),
.B1(n_7),
.B2(n_8),
.Y(n_154)
);

OA22x2_ASAP7_75t_L g161 ( 
.A1(n_57),
.A2(n_1),
.B1(n_8),
.B2(n_9),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_163),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_99),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_163),
.A2(n_167),
.B1(n_152),
.B2(n_117),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_105),
.A2(n_9),
.B1(n_107),
.B2(n_83),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_81),
.B(n_91),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_96),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_L g173 ( 
.A1(n_72),
.A2(n_94),
.B1(n_98),
.B2(n_110),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_85),
.A2(n_89),
.B1(n_66),
.B2(n_84),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_176),
.A2(n_167),
.B(n_179),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_110),
.B(n_102),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_182),
.C(n_133),
.Y(n_212)
);

AND2x2_ASAP7_75t_SL g182 ( 
.A(n_85),
.B(n_89),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_134),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_103),
.C(n_77),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_185),
.B(n_193),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_186),
.B(n_218),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_146),
.A2(n_168),
.B1(n_148),
.B2(n_134),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_187),
.A2(n_229),
.B1(n_231),
.B2(n_235),
.Y(n_255)
);

BUFx4f_ASAP7_75t_SL g188 ( 
.A(n_170),
.Y(n_188)
);

INVx13_ASAP7_75t_L g246 ( 
.A(n_188),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g251 ( 
.A(n_189),
.B(n_204),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_190),
.A2(n_195),
.B1(n_203),
.B2(n_244),
.Y(n_267)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_191),
.Y(n_278)
);

AOI21xp33_ASAP7_75t_L g285 ( 
.A1(n_192),
.A2(n_208),
.B(n_214),
.Y(n_285)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_194),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_128),
.A2(n_149),
.B1(n_124),
.B2(n_119),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_184),
.A2(n_178),
.B(n_168),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_197),
.A2(n_238),
.B(n_240),
.Y(n_274)
);

INVx4_ASAP7_75t_SL g198 ( 
.A(n_170),
.Y(n_198)
);

INVx13_ASAP7_75t_L g265 ( 
.A(n_198),
.Y(n_265)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_199),
.Y(n_254)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_171),
.Y(n_200)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_200),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_201),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_142),
.A2(n_130),
.B1(n_132),
.B2(n_180),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_141),
.A2(n_147),
.B1(n_127),
.B2(n_136),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_136),
.Y(n_205)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_205),
.Y(n_273)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_144),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_206),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_164),
.B(n_159),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_207),
.B(n_211),
.Y(n_261)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_209),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_144),
.Y(n_210)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_210),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_133),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_212),
.B(n_232),
.C(n_234),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_151),
.A2(n_143),
.B1(n_167),
.B2(n_123),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_213),
.A2(n_222),
.B1(n_234),
.B2(n_202),
.Y(n_247)
);

OR2x2_ASAP7_75t_SL g214 ( 
.A(n_161),
.B(n_165),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_157),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_215),
.Y(n_283)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_171),
.Y(n_216)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_216),
.Y(n_282)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_126),
.Y(n_217)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_217),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_126),
.B(n_174),
.Y(n_218)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_170),
.Y(n_219)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_219),
.Y(n_289)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_169),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g287 ( 
.A(n_220),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_161),
.B(n_140),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_221),
.B(n_223),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_115),
.B(n_135),
.Y(n_223)
);

BUFx12_ASAP7_75t_L g224 ( 
.A(n_148),
.Y(n_224)
);

INVx13_ASAP7_75t_L g276 ( 
.A(n_224),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_120),
.B(n_156),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_226),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_156),
.B(n_177),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_177),
.B(n_183),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_228),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_118),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_118),
.Y(n_229)
);

CKINVDCx9p33_ASAP7_75t_R g230 ( 
.A(n_176),
.Y(n_230)
);

BUFx12_ASAP7_75t_L g271 ( 
.A(n_230),
.Y(n_271)
);

CKINVDCx6p67_ASAP7_75t_R g231 ( 
.A(n_122),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_183),
.B(n_162),
.C(n_175),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_121),
.B(n_137),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_236),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_L g234 ( 
.A1(n_121),
.A2(n_137),
.B1(n_138),
.B2(n_162),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_138),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_175),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_129),
.B(n_184),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_241),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_179),
.A2(n_160),
.B(n_166),
.Y(n_240)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_158),
.Y(n_241)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_144),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_243),
.Y(n_258)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_158),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_247),
.A2(n_252),
.B1(n_251),
.B2(n_288),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_212),
.Y(n_249)
);

XOR2x2_ASAP7_75t_L g313 ( 
.A(n_249),
.B(n_269),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_190),
.A2(n_213),
.B1(n_196),
.B2(n_214),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_252),
.A2(n_272),
.B1(n_277),
.B2(n_281),
.Y(n_318)
);

A2O1A1Ixp33_ASAP7_75t_L g257 ( 
.A1(n_208),
.A2(n_197),
.B(n_239),
.C(n_232),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_257),
.B(n_274),
.Y(n_306)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_203),
.A2(n_187),
.B1(n_239),
.B2(n_231),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_264),
.A2(n_286),
.B1(n_271),
.B2(n_278),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_269),
.B(n_249),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_239),
.B(n_216),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_280),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_231),
.A2(n_217),
.B1(n_236),
.B2(n_210),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_200),
.A2(n_243),
.B1(n_194),
.B2(n_241),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_191),
.B(n_199),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_206),
.A2(n_242),
.B1(n_198),
.B2(n_188),
.Y(n_281)
);

O2A1O1Ixp33_ASAP7_75t_SL g286 ( 
.A1(n_224),
.A2(n_223),
.B(n_225),
.C(n_230),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_188),
.A2(n_190),
.B1(n_221),
.B2(n_202),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_288),
.A2(n_255),
.B1(n_281),
.B2(n_284),
.Y(n_319)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_258),
.Y(n_291)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_291),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_260),
.B(n_219),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_292),
.B(n_294),
.Y(n_328)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_258),
.Y(n_293)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_293),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_261),
.B(n_256),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_270),
.A2(n_224),
.B(n_257),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_295),
.A2(n_304),
.B(n_306),
.Y(n_351)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_280),
.Y(n_296)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_296),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_297),
.B(n_313),
.C(n_273),
.Y(n_331)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_279),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_298),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_250),
.B(n_268),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_299),
.B(n_316),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_261),
.B(n_256),
.Y(n_300)
);

INVxp33_ASAP7_75t_L g343 ( 
.A(n_300),
.Y(n_343)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_266),
.Y(n_301)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_301),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_262),
.B(n_274),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_302),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_250),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_303),
.B(n_308),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_248),
.A2(n_286),
.B(n_251),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_275),
.Y(n_305)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_305),
.Y(n_345)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_275),
.Y(n_307)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_307),
.Y(n_350)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_253),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_253),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_309),
.B(n_310),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_277),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_311),
.A2(n_319),
.B1(n_266),
.B2(n_263),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_245),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_312),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_272),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_314),
.B(n_320),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_247),
.A2(n_248),
.B1(n_267),
.B2(n_286),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_315),
.A2(n_317),
.B1(n_321),
.B2(n_323),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_259),
.B(n_283),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_285),
.A2(n_284),
.B1(n_279),
.B2(n_254),
.Y(n_317)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_282),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_254),
.A2(n_283),
.B1(n_259),
.B2(n_282),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_278),
.B(n_289),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_322),
.B(n_245),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_273),
.B(n_263),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_324),
.B(n_316),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_324),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_325),
.B(n_340),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_331),
.B(n_308),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_332),
.A2(n_318),
.B1(n_314),
.B2(n_310),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_336),
.B(n_349),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_313),
.B(n_289),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_339),
.B(n_297),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_321),
.Y(n_340)
);

AOI222xp33_ASAP7_75t_L g344 ( 
.A1(n_306),
.A2(n_265),
.B1(n_271),
.B2(n_246),
.C1(n_276),
.C2(n_287),
.Y(n_344)
);

XOR2x1_ASAP7_75t_L g367 ( 
.A(n_344),
.B(n_319),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_292),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_347),
.B(n_348),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_290),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_352),
.A2(n_356),
.B1(n_332),
.B2(n_338),
.Y(n_382)
);

AOI322xp5_ASAP7_75t_L g353 ( 
.A1(n_328),
.A2(n_299),
.A3(n_300),
.B1(n_290),
.B2(n_297),
.C1(n_315),
.C2(n_311),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_353),
.B(n_363),
.Y(n_375)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_346),
.Y(n_355)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_355),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_341),
.A2(n_332),
.B1(n_348),
.B2(n_340),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_346),
.Y(n_357)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_357),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_351),
.A2(n_295),
.B(n_304),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_358),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_334),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_359),
.B(n_362),
.Y(n_385)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_345),
.Y(n_361)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_361),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_325),
.B(n_303),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_328),
.B(n_343),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_345),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_364),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_365),
.B(n_339),
.Y(n_380)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_350),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_366),
.B(n_371),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_367),
.A2(n_372),
.B1(n_373),
.B2(n_341),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_333),
.B(n_291),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_369),
.A2(n_338),
.B1(n_335),
.B2(n_326),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_370),
.B(n_339),
.C(n_331),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_333),
.B(n_293),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_350),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_337),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_377),
.B(n_382),
.Y(n_397)
);

OA21x2_ASAP7_75t_SL g378 ( 
.A1(n_362),
.A2(n_327),
.B(n_329),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_378),
.B(n_368),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_380),
.B(n_384),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_370),
.B(n_313),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_383),
.B(n_354),
.C(n_309),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_386),
.A2(n_388),
.B1(n_352),
.B2(n_356),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_365),
.B(n_331),
.C(n_329),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_387),
.B(n_391),
.C(n_357),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_356),
.A2(n_330),
.B1(n_326),
.B2(n_335),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_365),
.B(n_330),
.C(n_351),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_393),
.B(n_394),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_390),
.A2(n_358),
.B(n_360),
.Y(n_394)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_395),
.Y(n_409)
);

AO221x1_ASAP7_75t_L g396 ( 
.A1(n_388),
.A2(n_317),
.B1(n_352),
.B2(n_347),
.C(n_363),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_396),
.B(n_403),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_374),
.B(n_294),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_398),
.B(n_399),
.Y(n_414)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_389),
.Y(n_399)
);

XOR2x1_ASAP7_75t_L g400 ( 
.A(n_385),
.B(n_367),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_400),
.B(n_401),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_383),
.B(n_354),
.C(n_336),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_402),
.B(n_381),
.C(n_391),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_375),
.B(n_368),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_387),
.B(n_371),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_404),
.B(n_377),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_405),
.B(n_384),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_407),
.B(n_412),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_408),
.B(n_411),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_401),
.B(n_380),
.C(n_390),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_397),
.A2(n_386),
.B1(n_355),
.B2(n_360),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_413),
.B(n_416),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_392),
.B(n_385),
.C(n_358),
.Y(n_416)
);

MAJx2_ASAP7_75t_L g418 ( 
.A(n_416),
.B(n_392),
.C(n_402),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_418),
.B(n_422),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_410),
.B(n_394),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_419),
.B(n_400),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_410),
.A2(n_405),
.B(n_397),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_420),
.A2(n_349),
.B(n_359),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_411),
.A2(n_353),
.B(n_369),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_414),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_423),
.B(n_369),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_425),
.B(n_431),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_417),
.A2(n_415),
.B1(n_409),
.B2(n_406),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_426),
.A2(n_424),
.B1(n_393),
.B2(n_382),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_428),
.B(n_419),
.Y(n_433)
);

INVx11_ASAP7_75t_L g429 ( 
.A(n_423),
.Y(n_429)
);

INVx11_ASAP7_75t_L g434 ( 
.A(n_429),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_421),
.B(n_407),
.C(n_412),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_430),
.B(n_418),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_432),
.A2(n_433),
.B1(n_425),
.B2(n_427),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_436),
.B(n_430),
.C(n_426),
.Y(n_437)
);

AOI322xp5_ASAP7_75t_L g440 ( 
.A1(n_437),
.A2(n_438),
.A3(n_439),
.B1(n_435),
.B2(n_434),
.C1(n_376),
.C2(n_432),
.Y(n_440)
);

AOI322xp5_ASAP7_75t_L g439 ( 
.A1(n_435),
.A2(n_431),
.A3(n_429),
.B1(n_428),
.B2(n_376),
.C1(n_361),
.C2(n_364),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_440),
.A2(n_441),
.B(n_379),
.Y(n_442)
);

AOI322xp5_ASAP7_75t_L g441 ( 
.A1(n_439),
.A2(n_434),
.A3(n_366),
.B1(n_372),
.B2(n_342),
.C1(n_296),
.C2(n_367),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_442),
.B(n_373),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_443),
.B(n_334),
.Y(n_444)
);


endmodule