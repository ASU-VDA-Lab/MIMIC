module fake_jpeg_10801_n_257 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_3),
.B(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_41),
.Y(n_111)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_19),
.Y(n_42)
);

CKINVDCx9p33_ASAP7_75t_R g99 ( 
.A(n_42),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_43),
.Y(n_70)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_61),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_17),
.B(n_15),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_50),
.B(n_64),
.Y(n_78)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

NAND2xp33_ASAP7_75t_SL g53 ( 
.A(n_20),
.B(n_2),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_20),
.B(n_32),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_60),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_2),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_63),
.Y(n_76)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_33),
.B(n_14),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_66),
.Y(n_75)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_68),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_23),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_34),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_79),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_73),
.B(n_85),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_26),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_34),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_81),
.B(n_89),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_38),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_87),
.B(n_94),
.Y(n_146)
);

CKINVDCx12_ASAP7_75t_R g88 ( 
.A(n_44),
.Y(n_88)
);

BUFx8_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_26),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_22),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_93),
.B(n_100),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_35),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_41),
.A2(n_47),
.B1(n_49),
.B2(n_54),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_12),
.B1(n_100),
.B2(n_104),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_63),
.A2(n_22),
.B1(n_29),
.B2(n_23),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_96),
.A2(n_71),
.B(n_75),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_21),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_52),
.A2(n_18),
.B1(n_23),
.B2(n_29),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_102),
.A2(n_109),
.B1(n_70),
.B2(n_108),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_51),
.B(n_21),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_103),
.B(n_104),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_16),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_48),
.A2(n_18),
.B1(n_16),
.B2(n_23),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_110),
.B1(n_45),
.B2(n_9),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_56),
.B(n_3),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_107),
.B(n_70),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_43),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_42),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_81),
.A2(n_45),
.B1(n_43),
.B2(n_10),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_113),
.A2(n_125),
.B1(n_127),
.B2(n_112),
.Y(n_164)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_114),
.Y(n_169)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_116),
.A2(n_131),
.B1(n_96),
.B2(n_97),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_99),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_122),
.Y(n_152)
);

OR2x4_ASAP7_75t_L g118 ( 
.A(n_73),
.B(n_6),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_118),
.Y(n_171)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_120),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_76),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_121),
.A2(n_127),
.B(n_113),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_89),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_123),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_78),
.B(n_11),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_124),
.B(n_126),
.Y(n_168)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_128),
.Y(n_165)
);

HAxp5_ASAP7_75t_SL g130 ( 
.A(n_72),
.B(n_79),
.CON(n_130),
.SN(n_130)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_134),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_80),
.Y(n_132)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_74),
.B(n_82),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_135),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_76),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_76),
.B(n_92),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_143),
.Y(n_160)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_92),
.B(n_93),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_136),
.C(n_127),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_83),
.B(n_90),
.Y(n_143)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_101),
.A2(n_111),
.B1(n_106),
.B2(n_80),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_145),
.A2(n_101),
.B1(n_106),
.B2(n_111),
.Y(n_148)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_77),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_161),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_112),
.B(n_71),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_167),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_97),
.B(n_91),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_132),
.B(n_142),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_91),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_91),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_163),
.B(n_164),
.Y(n_181)
);

AND2x2_ASAP7_75t_SL g167 ( 
.A(n_136),
.B(n_130),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_170),
.B(n_129),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_116),
.Y(n_192)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_132),
.Y(n_174)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_174),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_142),
.Y(n_180)
);

A2O1A1O1Ixp25_ASAP7_75t_L g205 ( 
.A1(n_180),
.A2(n_185),
.B(n_151),
.C(n_157),
.D(n_166),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_182),
.A2(n_170),
.B(n_171),
.Y(n_199)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_119),
.Y(n_185)
);

AND2x6_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_118),
.Y(n_186)
);

AOI221xp5_ASAP7_75t_L g208 ( 
.A1(n_186),
.A2(n_157),
.B1(n_129),
.B2(n_166),
.C(n_162),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_187),
.B(n_158),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_152),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_190),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_150),
.A2(n_121),
.B(n_139),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_189),
.A2(n_194),
.B(n_165),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_159),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_174),
.Y(n_191)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_191),
.Y(n_210)
);

OAI21x1_ASAP7_75t_L g198 ( 
.A1(n_192),
.A2(n_150),
.B(n_160),
.Y(n_198)
);

INVx4_ASAP7_75t_SL g193 ( 
.A(n_162),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_193),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_150),
.A2(n_114),
.B(n_138),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_147),
.Y(n_195)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_195),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_168),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_185),
.Y(n_203)
);

AO32x1_ASAP7_75t_L g217 ( 
.A1(n_198),
.A2(n_199),
.A3(n_189),
.B1(n_186),
.B2(n_200),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_199),
.A2(n_200),
.B(n_182),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_177),
.A2(n_161),
.B(n_164),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_177),
.A2(n_172),
.B1(n_151),
.B2(n_148),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_201),
.A2(n_206),
.B(n_208),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_205),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_204),
.B(n_176),
.Y(n_220)
);

OAI32xp33_ASAP7_75t_L g209 ( 
.A1(n_181),
.A2(n_165),
.A3(n_128),
.B1(n_140),
.B2(n_169),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_214),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_178),
.A2(n_145),
.B1(n_149),
.B2(n_169),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_213),
.A2(n_183),
.B1(n_191),
.B2(n_179),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_195),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_212),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_226),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_216),
.A2(n_217),
.B(n_218),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_206),
.A2(n_178),
.B1(n_175),
.B2(n_180),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_218),
.A2(n_221),
.B1(n_201),
.B2(n_211),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_220),
.B(n_219),
.Y(n_232)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_210),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_224),
.Y(n_230)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_202),
.A2(n_175),
.B(n_194),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_227),
.A2(n_197),
.B1(n_184),
.B2(n_179),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_204),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_229),
.C(n_232),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_176),
.C(n_205),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_231),
.A2(n_223),
.B(n_209),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_233),
.A2(n_211),
.B1(n_207),
.B2(n_225),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_235),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_221),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_237),
.B(n_241),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_236),
.A2(n_216),
.B(n_223),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_232),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_226),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_240),
.B(n_242),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_149),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_243),
.C(n_239),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_245),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_243),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_246),
.A2(n_229),
.B1(n_228),
.B2(n_215),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_249),
.A2(n_244),
.B1(n_247),
.B2(n_173),
.Y(n_252)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_248),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_250),
.A2(n_193),
.B(n_129),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_253),
.C(n_251),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_251),
.C(n_173),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_120),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_144),
.Y(n_257)
);


endmodule