module fake_jpeg_4996_n_210 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_210);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_210;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_30),
.B(n_31),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_23),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_34),
.A2(n_28),
.B1(n_26),
.B2(n_16),
.Y(n_70)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_14),
.B(n_1),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_36),
.B(n_26),
.Y(n_76)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_39),
.B(n_45),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_40),
.Y(n_72)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_42),
.B(n_44),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_24),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_15),
.B(n_1),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_46),
.B(n_20),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_55),
.Y(n_84)
);

NOR2x1_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_25),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_51),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_16),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_76),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_58),
.Y(n_85)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_64),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_30),
.B(n_27),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_61),
.Y(n_106)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_62),
.A2(n_65),
.B1(n_70),
.B2(n_9),
.Y(n_101)
);

NOR2x1_ASAP7_75t_L g63 ( 
.A(n_32),
.B(n_28),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_63),
.B(n_68),
.Y(n_107)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_32),
.B(n_18),
.Y(n_66)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_69),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_18),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_41),
.B(n_15),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_75),
.Y(n_105)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_36),
.B(n_20),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_42),
.B(n_11),
.Y(n_81)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_42),
.B(n_4),
.Y(n_82)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_29),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_86),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_29),
.C(n_22),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_90),
.A2(n_98),
.B(n_73),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_70),
.A2(n_21),
.B1(n_22),
.B2(n_7),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_50),
.A2(n_5),
.B(n_6),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_9),
.B1(n_6),
.B2(n_8),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_47),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_71),
.A2(n_9),
.B1(n_65),
.B2(n_59),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_52),
.B1(n_72),
.B2(n_57),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_126),
.B1(n_127),
.B2(n_130),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_123),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_54),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_112),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_48),
.Y(n_111)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

BUFx4f_ASAP7_75t_SL g113 ( 
.A(n_93),
.Y(n_113)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_116),
.Y(n_141)
);

OA21x2_ASAP7_75t_L g115 ( 
.A1(n_104),
.A2(n_60),
.B(n_56),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_115),
.A2(n_97),
.B1(n_89),
.B2(n_92),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_94),
.B(n_80),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_94),
.B(n_77),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_118),
.Y(n_151)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_58),
.Y(n_119)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_120),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_86),
.B(n_71),
.Y(n_121)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_73),
.Y(n_122)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_64),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_124),
.A2(n_95),
.B1(n_99),
.B2(n_90),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_55),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_125),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_97),
.B(n_52),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_74),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g146 ( 
.A1(n_131),
.A2(n_128),
.B(n_89),
.Y(n_146)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_100),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_139),
.C(n_145),
.Y(n_154)
);

MAJx2_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_91),
.C(n_105),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_115),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_92),
.C(n_98),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_146),
.B(n_115),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_106),
.C(n_102),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_115),
.Y(n_167)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_156),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_135),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_143),
.A2(n_126),
.B(n_127),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_131),
.Y(n_158)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

NOR2xp67_ASAP7_75t_SL g159 ( 
.A(n_139),
.B(n_147),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_SL g168 ( 
.A(n_159),
.B(n_163),
.C(n_134),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_162),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_167),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_135),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_132),
.B(n_106),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_164),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_146),
.B(n_112),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_152),
.C(n_145),
.Y(n_169)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_166),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_168),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_175),
.C(n_166),
.Y(n_185)
);

OAI21x1_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_144),
.B(n_142),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_SL g189 ( 
.A(n_170),
.B(n_110),
.C(n_113),
.Y(n_189)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_137),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_158),
.C(n_167),
.Y(n_183)
);

XNOR2x1_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_138),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_174),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_183),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_173),
.A2(n_155),
.B1(n_153),
.B2(n_164),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_185),
.Y(n_193)
);

INVxp33_ASAP7_75t_SL g186 ( 
.A(n_172),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_186),
.A2(n_177),
.B(n_148),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_114),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_136),
.Y(n_195)
);

AOI31xp67_ASAP7_75t_L g196 ( 
.A1(n_189),
.A2(n_186),
.A3(n_180),
.B(n_176),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_181),
.B(n_140),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_192),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_189),
.A2(n_173),
.B(n_171),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_195),
.C(n_149),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_196),
.A2(n_120),
.B1(n_180),
.B2(n_150),
.Y(n_198)
);

NAND4xp25_ASAP7_75t_SL g197 ( 
.A(n_192),
.B(n_113),
.C(n_187),
.D(n_129),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_150),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_198),
.B(n_199),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_183),
.C(n_179),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_193),
.Y(n_202)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_202),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_200),
.Y(n_204)
);

OAI321xp33_ASAP7_75t_L g207 ( 
.A1(n_205),
.A2(n_113),
.A3(n_200),
.B1(n_118),
.B2(n_178),
.C(n_124),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_207),
.B(n_203),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_208),
.B(n_209),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_206),
.B(n_204),
.Y(n_209)
);


endmodule