module real_aes_17328_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_863, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_863;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_635;
wire n_287;
wire n_357;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_860;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_0), .Y(n_214) );
AND2x4_ASAP7_75t_L g858 ( .A(n_1), .B(n_859), .Y(n_858) );
INVx1_ASAP7_75t_SL g833 ( .A(n_2), .Y(n_833) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_3), .A2(n_5), .B1(n_161), .B2(n_565), .Y(n_564) );
AOI21xp33_ASAP7_75t_SL g837 ( .A1(n_4), .A2(n_838), .B(n_845), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_6), .A2(n_21), .B1(n_124), .B2(n_164), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_7), .A2(n_53), .B1(n_212), .B2(n_514), .Y(n_513) );
BUFx3_ASAP7_75t_L g155 ( .A(n_8), .Y(n_155) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_9), .A2(n_15), .B1(n_501), .B2(n_528), .Y(n_539) );
INVx1_ASAP7_75t_L g859 ( .A(n_10), .Y(n_859) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_11), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_12), .B(n_127), .Y(n_126) );
OR2x2_ASAP7_75t_L g819 ( .A(n_13), .B(n_31), .Y(n_819) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_14), .Y(n_125) );
AOI22xp5_ASAP7_75t_L g806 ( .A1(n_16), .A2(n_83), .B1(n_807), .B2(n_808), .Y(n_806) );
INVx1_ASAP7_75t_L g808 ( .A(n_16), .Y(n_808) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_17), .B(n_149), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_18), .B(n_174), .Y(n_173) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_19), .A2(n_84), .B1(n_124), .B2(n_149), .Y(n_223) );
OAI21x1_ASAP7_75t_L g119 ( .A1(n_20), .A2(n_48), .B(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_22), .B(n_164), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g637 ( .A(n_23), .Y(n_637) );
INVx4_ASAP7_75t_R g553 ( .A(n_24), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_25), .B(n_129), .Y(n_586) );
AO32x2_ASAP7_75t_L g220 ( .A1(n_26), .A2(n_141), .A3(n_142), .B1(n_221), .B2(n_224), .Y(n_220) );
AO32x1_ASAP7_75t_L g258 ( .A1(n_26), .A2(n_141), .A3(n_142), .B1(n_221), .B2(n_224), .Y(n_258) );
INVx1_ASAP7_75t_L g567 ( .A(n_27), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_28), .B(n_164), .Y(n_592) );
A2O1A1Ixp33_ASAP7_75t_SL g500 ( .A1(n_29), .A2(n_128), .B(n_501), .C(n_502), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_30), .A2(n_45), .B1(n_132), .B2(n_501), .Y(n_635) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_32), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_33), .A2(n_51), .B1(n_152), .B2(n_164), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_34), .A2(n_89), .B1(n_124), .B2(n_132), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_35), .B(n_131), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g834 ( .A(n_36), .Y(n_834) );
INVx1_ASAP7_75t_L g836 ( .A(n_36), .Y(n_836) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_37), .B(n_187), .Y(n_247) );
INVx1_ASAP7_75t_L g589 ( .A(n_38), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_39), .A2(n_67), .B1(n_132), .B2(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_40), .B(n_501), .Y(n_591) );
CKINVDCx5p33_ASAP7_75t_R g529 ( .A(n_41), .Y(n_529) );
INVx2_ASAP7_75t_L g814 ( .A(n_42), .Y(n_814) );
BUFx3_ASAP7_75t_L g817 ( .A(n_43), .Y(n_817) );
INVx1_ASAP7_75t_L g828 ( .A(n_43), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_44), .B(n_249), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_46), .A2(n_85), .B1(n_132), .B2(n_501), .Y(n_540) );
CKINVDCx5p33_ASAP7_75t_R g554 ( .A(n_47), .Y(n_554) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_49), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_50), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_52), .A2(n_77), .B1(n_186), .B2(n_187), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_54), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g148 ( .A1(n_55), .A2(n_81), .B1(n_124), .B2(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g120 ( .A(n_56), .Y(n_120) );
AND2x4_ASAP7_75t_L g138 ( .A(n_57), .B(n_139), .Y(n_138) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_58), .A2(n_90), .B1(n_132), .B2(n_563), .Y(n_562) );
AO22x1_ASAP7_75t_L g518 ( .A1(n_59), .A2(n_72), .B1(n_519), .B2(n_520), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_60), .B(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g139 ( .A(n_61), .Y(n_139) );
AND2x2_ASAP7_75t_L g504 ( .A(n_62), .B(n_141), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_63), .B(n_141), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_64), .A2(n_212), .B(n_213), .C(n_215), .Y(n_211) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_65), .A2(n_102), .B1(n_851), .B2(n_860), .Y(n_101) );
NAND3xp33_ASAP7_75t_L g136 ( .A(n_66), .B(n_124), .C(n_134), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g497 ( .A(n_68), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_69), .B(n_212), .Y(n_533) );
AND2x2_ASAP7_75t_L g217 ( .A(n_70), .B(n_218), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_71), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_73), .B(n_164), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_74), .A2(n_94), .B1(n_149), .B2(n_186), .Y(n_190) );
INVx2_ASAP7_75t_L g129 ( .A(n_75), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_76), .B(n_168), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_78), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_79), .B(n_141), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_80), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_82), .B(n_118), .Y(n_516) );
INVx1_ASAP7_75t_L g807 ( .A(n_83), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_86), .B(n_134), .Y(n_133) );
AOI22xp33_ASAP7_75t_L g151 ( .A1(n_87), .A2(n_100), .B1(n_132), .B2(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_88), .B(n_187), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_91), .B(n_141), .Y(n_525) );
INVx1_ASAP7_75t_L g482 ( .A(n_92), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g848 ( .A(n_92), .B(n_849), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_93), .B(n_174), .Y(n_250) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_95), .A2(n_189), .B(n_212), .C(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g556 ( .A(n_96), .B(n_218), .Y(n_556) );
INVxp67_ASAP7_75t_SL g850 ( .A(n_97), .Y(n_850) );
NAND2xp33_ASAP7_75t_L g532 ( .A(n_98), .B(n_127), .Y(n_532) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_99), .Y(n_160) );
AO21x2_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_810), .B(n_820), .Y(n_102) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_805), .B1(n_806), .B2(n_809), .Y(n_103) );
INVxp33_ASAP7_75t_SL g809 ( .A(n_104), .Y(n_809) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_480), .B1(n_483), .B2(n_487), .Y(n_104) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_390), .Y(n_105) );
NAND4xp25_ASAP7_75t_L g106 ( .A(n_107), .B(n_295), .C(n_322), .D(n_358), .Y(n_106) );
AOI221x1_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_200), .B1(n_234), .B2(n_270), .C(n_274), .Y(n_107) );
NAND3xp33_ASAP7_75t_L g108 ( .A(n_109), .B(n_176), .C(n_198), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_143), .Y(n_111) );
INVx2_ASAP7_75t_L g235 ( .A(n_112), .Y(n_235) );
AND2x2_ASAP7_75t_L g408 ( .A(n_112), .B(n_352), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_112), .B(n_199), .Y(n_417) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g423 ( .A(n_113), .Y(n_423) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g268 ( .A(n_114), .Y(n_268) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OR2x2_ASAP7_75t_L g351 ( .A(n_115), .B(n_197), .Y(n_351) );
OAI21x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_140), .Y(n_115) );
OAI21xp5_ASAP7_75t_L g280 ( .A1(n_116), .A2(n_121), .B(n_140), .Y(n_280) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AO31x2_ASAP7_75t_L g537 ( .A1(n_117), .A2(n_538), .A3(n_542), .B(n_543), .Y(n_537) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g175 ( .A(n_118), .Y(n_175) );
INVx2_ASAP7_75t_L g195 ( .A(n_118), .Y(n_195) );
OAI21xp33_ASAP7_75t_L g522 ( .A1(n_118), .A2(n_216), .B(n_516), .Y(n_522) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_119), .Y(n_142) );
OAI21x1_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_130), .B(n_137), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_126), .B(n_128), .Y(n_122) );
INVx2_ASAP7_75t_SL g187 ( .A(n_124), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_124), .B(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_125), .Y(n_127) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_125), .Y(n_132) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_125), .Y(n_149) );
INVx1_ASAP7_75t_L g152 ( .A(n_125), .Y(n_152) );
INVx1_ASAP7_75t_L g162 ( .A(n_125), .Y(n_162) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_125), .Y(n_164) );
INVx1_ASAP7_75t_L g186 ( .A(n_125), .Y(n_186) );
INVx1_ASAP7_75t_L g212 ( .A(n_125), .Y(n_212) );
INVx3_ASAP7_75t_L g501 ( .A(n_125), .Y(n_501) );
INVx1_ASAP7_75t_L g515 ( .A(n_125), .Y(n_515) );
OAI22xp33_ASAP7_75t_L g552 ( .A1(n_127), .A2(n_152), .B1(n_553), .B2(n_554), .Y(n_552) );
INVx2_ASAP7_75t_L g563 ( .A(n_127), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g147 ( .A1(n_128), .A2(n_148), .B1(n_150), .B2(n_151), .Y(n_147) );
INVx6_ASAP7_75t_L g150 ( .A(n_128), .Y(n_150) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_128), .A2(n_165), .B1(n_222), .B2(n_223), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_128), .B(n_518), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_128), .A2(n_532), .B(n_533), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_L g575 ( .A1(n_128), .A2(n_512), .B(n_518), .C(n_522), .Y(n_575) );
BUFx8_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g135 ( .A(n_129), .Y(n_135) );
INVx2_ASAP7_75t_L g170 ( .A(n_129), .Y(n_170) );
INVx1_ASAP7_75t_L g189 ( .A(n_129), .Y(n_189) );
OAI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_133), .B(n_136), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g565 ( .A(n_132), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_132), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx4f_ASAP7_75t_L g165 ( .A(n_135), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_135), .B(n_589), .Y(n_588) );
AOI31xp67_ASAP7_75t_L g145 ( .A1(n_137), .A2(n_146), .A3(n_147), .B(n_153), .Y(n_145) );
OAI21x1_ASAP7_75t_L g158 ( .A1(n_137), .A2(n_159), .B(n_166), .Y(n_158) );
INVx1_ASAP7_75t_L g535 ( .A(n_137), .Y(n_535) );
AND2x2_ASAP7_75t_L g593 ( .A(n_137), .B(n_142), .Y(n_593) );
AO31x2_ASAP7_75t_L g632 ( .A1(n_137), .A2(n_146), .A3(n_633), .B(n_636), .Y(n_632) );
BUFx10_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g192 ( .A(n_138), .Y(n_192) );
INVx1_ASAP7_75t_L g216 ( .A(n_138), .Y(n_216) );
AO31x2_ASAP7_75t_L g226 ( .A1(n_138), .A2(n_183), .A3(n_227), .B(n_232), .Y(n_226) );
BUFx10_ASAP7_75t_L g542 ( .A(n_138), .Y(n_542) );
INVx2_ASAP7_75t_L g146 ( .A(n_141), .Y(n_146) );
NOR2x1_ASAP7_75t_L g534 ( .A(n_141), .B(n_535), .Y(n_534) );
INVx4_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_142), .B(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g157 ( .A(n_142), .Y(n_157) );
BUFx3_ASAP7_75t_L g183 ( .A(n_142), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_142), .B(n_233), .Y(n_232) );
INVx2_ASAP7_75t_SL g241 ( .A(n_142), .Y(n_241) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_143), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_143), .B(n_379), .Y(n_378) );
INVxp67_ASAP7_75t_L g421 ( .A(n_143), .Y(n_421) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_156), .Y(n_143) );
AND2x2_ASAP7_75t_L g199 ( .A(n_144), .B(n_182), .Y(n_199) );
INVx2_ASAP7_75t_L g277 ( .A(n_144), .Y(n_277) );
AND2x2_ASAP7_75t_L g342 ( .A(n_144), .B(n_280), .Y(n_342) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g197 ( .A(n_145), .Y(n_197) );
INVx3_ASAP7_75t_L g249 ( .A(n_149), .Y(n_249) );
INVxp67_ASAP7_75t_SL g519 ( .A(n_149), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g184 ( .A1(n_150), .A2(n_185), .B1(n_188), .B2(n_190), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g227 ( .A1(n_150), .A2(n_228), .B1(n_230), .B2(n_231), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_150), .A2(n_247), .B(n_248), .Y(n_246) );
OAI22x1_ASAP7_75t_L g538 ( .A1(n_150), .A2(n_539), .B1(n_540), .B2(n_541), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_150), .A2(n_541), .B1(n_562), .B2(n_564), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_150), .A2(n_231), .B1(n_634), .B2(n_635), .Y(n_633) );
INVx1_ASAP7_75t_L g171 ( .A(n_152), .Y(n_171) );
OAI22xp5_ASAP7_75t_L g207 ( .A1(n_152), .A2(n_164), .B1(n_208), .B2(n_209), .Y(n_207) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g269 ( .A(n_156), .Y(n_269) );
AND2x2_ASAP7_75t_L g279 ( .A(n_156), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g341 ( .A(n_156), .B(n_182), .Y(n_341) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_173), .Y(n_156) );
OA21x2_ASAP7_75t_L g179 ( .A1(n_157), .A2(n_158), .B(n_173), .Y(n_179) );
O2A1O1Ixp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_161), .B(n_163), .C(n_165), .Y(n_159) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_162), .B(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g229 ( .A(n_164), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_164), .B(n_497), .Y(n_496) );
OAI21xp5_ASAP7_75t_L g495 ( .A1(n_165), .A2(n_496), .B(n_498), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_169), .B1(n_171), .B2(n_172), .Y(n_166) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_168), .A2(n_528), .B(n_529), .C(n_530), .Y(n_527) );
INVx2_ASAP7_75t_SL g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
BUFx3_ASAP7_75t_L g215 ( .A(n_170), .Y(n_215) );
INVx2_ASAP7_75t_L g204 ( .A(n_174), .Y(n_204) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g306 ( .A(n_176), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_177), .B(n_180), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_178), .B(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_178), .B(n_321), .Y(n_320) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_178), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_178), .B(n_376), .Y(n_383) );
INVx2_ASAP7_75t_SL g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g352 ( .A(n_179), .B(n_327), .Y(n_352) );
OR2x2_ASAP7_75t_L g354 ( .A(n_179), .B(n_280), .Y(n_354) );
INVx1_ASAP7_75t_L g413 ( .A(n_179), .Y(n_413) );
BUFx2_ASAP7_75t_L g427 ( .A(n_179), .Y(n_427) );
OR2x2_ASAP7_75t_L g455 ( .A(n_179), .B(n_182), .Y(n_455) );
INVx1_ASAP7_75t_L g474 ( .A(n_180), .Y(n_474) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g321 ( .A(n_181), .Y(n_321) );
OR2x2_ASAP7_75t_L g334 ( .A(n_181), .B(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g353 ( .A(n_181), .B(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g181 ( .A(n_182), .B(n_196), .Y(n_181) );
INVx2_ASAP7_75t_L g273 ( .A(n_182), .Y(n_273) );
AND2x2_ASAP7_75t_L g289 ( .A(n_182), .B(n_196), .Y(n_289) );
INVx1_ASAP7_75t_L g327 ( .A(n_182), .Y(n_327) );
INVx1_ASAP7_75t_L g370 ( .A(n_182), .Y(n_370) );
AND2x2_ASAP7_75t_L g412 ( .A(n_182), .B(n_413), .Y(n_412) );
AO31x2_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .A3(n_191), .B(n_193), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_186), .B(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g520 ( .A(n_186), .Y(n_520) );
INVx1_ASAP7_75t_SL g188 ( .A(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g210 ( .A(n_189), .Y(n_210) );
INVx1_ASAP7_75t_L g541 ( .A(n_189), .Y(n_541) );
AO31x2_ASAP7_75t_L g560 ( .A1(n_191), .A2(n_493), .A3(n_561), .B(n_566), .Y(n_560) );
INVx2_ASAP7_75t_SL g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_SL g224 ( .A(n_192), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
INVx2_ASAP7_75t_L g218 ( .A(n_195), .Y(n_218) );
BUFx2_ASAP7_75t_L g493 ( .A(n_195), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_195), .B(n_544), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_195), .B(n_567), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_195), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g468 ( .A(n_198), .Y(n_468) );
AND2x4_ASAP7_75t_L g406 ( .A(n_199), .B(n_266), .Y(n_406) );
INVx2_ASAP7_75t_L g435 ( .A(n_199), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_199), .B(n_427), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_200), .B(n_425), .Y(n_424) );
AND2x4_ASAP7_75t_L g200 ( .A(n_201), .B(n_219), .Y(n_200) );
AND2x2_ASAP7_75t_L g346 ( .A(n_201), .B(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g367 ( .A(n_201), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
OR2x2_ASAP7_75t_L g238 ( .A(n_202), .B(n_239), .Y(n_238) );
OR2x2_ASAP7_75t_L g262 ( .A(n_202), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g293 ( .A(n_202), .Y(n_293) );
AND2x2_ASAP7_75t_L g333 ( .A(n_202), .B(n_225), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_202), .B(n_317), .Y(n_374) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g286 ( .A(n_203), .Y(n_286) );
AOI21x1_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_217), .Y(n_203) );
AO21x2_ASAP7_75t_L g546 ( .A1(n_204), .A2(n_547), .B(n_556), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_211), .B(n_216), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_207), .B(n_210), .Y(n_206) );
INVx2_ASAP7_75t_L g231 ( .A(n_215), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_216), .A2(n_495), .B(n_500), .Y(n_494) );
INVx3_ASAP7_75t_L g252 ( .A(n_219), .Y(n_252) );
AND2x2_ASAP7_75t_L g297 ( .A(n_219), .B(n_292), .Y(n_297) );
AND2x2_ASAP7_75t_L g452 ( .A(n_219), .B(n_256), .Y(n_452) );
AND2x4_ASAP7_75t_L g219 ( .A(n_220), .B(n_225), .Y(n_219) );
INVx1_ASAP7_75t_L g303 ( .A(n_220), .Y(n_303) );
AND2x2_ASAP7_75t_L g331 ( .A(n_220), .B(n_239), .Y(n_331) );
OAI21x1_ASAP7_75t_L g242 ( .A1(n_224), .A2(n_243), .B(n_246), .Y(n_242) );
AND2x4_ASAP7_75t_L g284 ( .A(n_225), .B(n_285), .Y(n_284) );
INVx3_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
OR2x2_ASAP7_75t_L g257 ( .A(n_226), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g294 ( .A(n_226), .B(n_258), .Y(n_294) );
AND2x2_ASAP7_75t_L g304 ( .A(n_226), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_226), .B(n_239), .Y(n_356) );
AND2x2_ASAP7_75t_L g362 ( .A(n_226), .B(n_286), .Y(n_362) );
AOI21x1_ASAP7_75t_L g243 ( .A1(n_231), .A2(n_244), .B(n_245), .Y(n_243) );
OAI21x1_ASAP7_75t_L g512 ( .A1(n_231), .A2(n_513), .B(n_516), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g590 ( .A1(n_231), .A2(n_591), .B(n_592), .Y(n_590) );
OAI21xp33_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B(n_253), .Y(n_234) );
OAI21xp33_ASAP7_75t_L g395 ( .A1(n_235), .A2(n_396), .B(n_400), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_235), .B(n_426), .Y(n_473) );
NAND2x1_ASAP7_75t_SL g236 ( .A(n_237), .B(n_251), .Y(n_236) );
INVx1_ASAP7_75t_L g479 ( .A(n_237), .Y(n_479) );
INVx3_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
BUFx2_ASAP7_75t_L g256 ( .A(n_239), .Y(n_256) );
INVx2_ASAP7_75t_L g261 ( .A(n_239), .Y(n_261) );
INVxp67_ASAP7_75t_L g282 ( .A(n_239), .Y(n_282) );
AND2x2_ASAP7_75t_L g302 ( .A(n_239), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g313 ( .A(n_239), .B(n_314), .Y(n_313) );
INVx3_ASAP7_75t_L g317 ( .A(n_239), .Y(n_317) );
INVx1_ASAP7_75t_L g335 ( .A(n_239), .Y(n_335) );
OR2x2_ASAP7_75t_L g368 ( .A(n_239), .B(n_303), .Y(n_368) );
INVx1_ASAP7_75t_L g439 ( .A(n_239), .Y(n_439) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
OAI21x1_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B(n_250), .Y(n_240) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
OAI21xp33_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_259), .B(n_264), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
OAI22xp33_ASAP7_75t_L g377 ( .A1(n_255), .A2(n_378), .B1(n_380), .B2(n_383), .Y(n_377) );
OR2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_256), .B(n_304), .Y(n_338) );
BUFx2_ASAP7_75t_L g397 ( .A(n_256), .Y(n_397) );
INVx2_ASAP7_75t_L g347 ( .A(n_257), .Y(n_347) );
OR2x2_ASAP7_75t_L g431 ( .A(n_257), .B(n_261), .Y(n_431) );
INVx1_ASAP7_75t_L g263 ( .A(n_258), .Y(n_263) );
INVx1_ASAP7_75t_L g312 ( .A(n_258), .Y(n_312) );
NOR2x1p5_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
INVxp67_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_261), .Y(n_382) );
OR2x2_ASAP7_75t_L g466 ( .A(n_261), .B(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g469 ( .A(n_261), .B(n_304), .Y(n_469) );
INVxp67_ASAP7_75t_SL g432 ( .A(n_262), .Y(n_432) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_266), .B(n_326), .Y(n_388) );
AND2x2_ASAP7_75t_L g478 ( .A(n_266), .B(n_276), .Y(n_478) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g387 ( .A(n_267), .B(n_276), .Y(n_387) );
NAND2x1p5_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
AND2x2_ASAP7_75t_L g344 ( .A(n_268), .B(n_277), .Y(n_344) );
AND2x2_ASAP7_75t_L g379 ( .A(n_268), .B(n_273), .Y(n_379) );
INVxp67_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g298 ( .A(n_271), .B(n_279), .Y(n_298) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g438 ( .A(n_273), .B(n_439), .Y(n_438) );
OAI22xp33_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_281), .B1(n_287), .B2(n_290), .Y(n_274) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_275), .A2(n_476), .B(n_477), .C(n_479), .Y(n_475) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g326 ( .A(n_277), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g394 ( .A(n_277), .Y(n_394) );
OR2x2_ASAP7_75t_L g441 ( .A(n_278), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AND2x2_ASAP7_75t_L g296 ( .A(n_282), .B(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g399 ( .A(n_285), .Y(n_399) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g305 ( .A(n_286), .Y(n_305) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_286), .Y(n_314) );
INVx1_ASAP7_75t_L g386 ( .A(n_286), .Y(n_386) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g442 ( .A(n_289), .Y(n_442) );
AND2x2_ASAP7_75t_L g464 ( .A(n_289), .B(n_427), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_290), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g316 ( .A(n_294), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g372 ( .A(n_294), .B(n_373), .Y(n_372) );
INVx2_ASAP7_75t_SL g467 ( .A(n_294), .Y(n_467) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_298), .B1(n_299), .B2(n_306), .C(n_307), .Y(n_295) );
INVxp67_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVx2_ASAP7_75t_L g389 ( .A(n_302), .Y(n_389) );
BUFx2_ASAP7_75t_L g409 ( .A(n_304), .Y(n_409) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_315), .B(n_318), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x4_ASAP7_75t_L g309 ( .A(n_310), .B(n_313), .Y(n_309) );
AND2x2_ASAP7_75t_L g451 ( .A(n_310), .B(n_373), .Y(n_451) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g357 ( .A(n_312), .Y(n_357) );
AND2x2_ASAP7_75t_L g447 ( .A(n_312), .B(n_317), .Y(n_447) );
INVx1_ASAP7_75t_L g330 ( .A(n_314), .Y(n_330) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AOI211xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_324), .B(n_336), .C(n_348), .Y(n_322) );
OAI22xp33_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_328), .B1(n_332), .B2(n_334), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
BUFx2_ASAP7_75t_L g364 ( .A(n_331), .Y(n_364) );
AND2x2_ASAP7_75t_L g457 ( .A(n_331), .B(n_399), .Y(n_457) );
OAI21xp33_ASAP7_75t_L g460 ( .A1(n_332), .A2(n_461), .B(n_463), .Y(n_460) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_339), .B1(n_343), .B2(n_345), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_339), .B(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVxp67_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x4_ASAP7_75t_L g411 ( .A(n_344), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x4_ASAP7_75t_L g398 ( .A(n_347), .B(n_399), .Y(n_398) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_347), .Y(n_414) );
AOI21xp33_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_353), .B(n_355), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
AND2x2_ASAP7_75t_L g425 ( .A(n_350), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g462 ( .A(n_350), .B(n_427), .Y(n_462) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g376 ( .A(n_351), .Y(n_376) );
OR2x2_ASAP7_75t_L g454 ( .A(n_351), .B(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g369 ( .A(n_354), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g401 ( .A(n_354), .Y(n_401) );
OR2x2_ASAP7_75t_L g434 ( .A(n_354), .B(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g405 ( .A(n_355), .Y(n_405) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
NOR3xp33_ASAP7_75t_L g358 ( .A(n_359), .B(n_377), .C(n_384), .Y(n_358) );
OAI322xp33_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_363), .A3(n_365), .B1(n_367), .B2(n_369), .C1(n_371), .C2(n_375), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
A2O1A1Ixp33_ASAP7_75t_L g436 ( .A1(n_361), .A2(n_401), .B(n_437), .C(n_440), .Y(n_436) );
BUFx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g381 ( .A(n_362), .B(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g418 ( .A(n_362), .Y(n_418) );
AND2x4_ASAP7_75t_L g446 ( .A(n_362), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AOI32xp33_ASAP7_75t_L g415 ( .A1(n_364), .A2(n_402), .A3(n_416), .B1(n_418), .B2(n_419), .Y(n_415) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g402 ( .A(n_368), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_370), .B(n_423), .Y(n_422) );
INVxp67_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
O2A1O1Ixp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_387), .B(n_388), .C(n_389), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_391), .B(n_448), .Y(n_390) );
AOI211xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_395), .B(n_403), .C(n_428), .Y(n_391) );
INVxp67_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
O2A1O1Ixp33_ASAP7_75t_SL g470 ( .A1(n_396), .A2(n_471), .B(n_472), .C(n_474), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
OAI31xp33_ASAP7_75t_L g450 ( .A1(n_398), .A2(n_451), .A3(n_452), .B(n_453), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
INVx2_ASAP7_75t_L g410 ( .A(n_402), .Y(n_410) );
NAND4xp25_ASAP7_75t_SL g403 ( .A(n_404), .B(n_407), .C(n_415), .D(n_424), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
AOI32xp33_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .A3(n_410), .B1(n_411), .B2(n_414), .Y(n_407) );
INVx1_ASAP7_75t_L g459 ( .A(n_411), .Y(n_459) );
INVx1_ASAP7_75t_L g471 ( .A(n_414), .Y(n_471) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NAND3xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_436), .C(n_443), .Y(n_428) );
OAI21xp5_ASAP7_75t_SL g429 ( .A1(n_430), .A2(n_432), .B(n_433), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx3_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_437), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_446), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
NOR4xp25_ASAP7_75t_L g448 ( .A(n_449), .B(n_460), .C(n_470), .D(n_475), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_456), .Y(n_449) );
OAI21xp33_ASAP7_75t_L g456 ( .A1(n_451), .A2(n_457), .B(n_458), .Y(n_456) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B1(n_468), .B2(n_469), .Y(n_463) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_467), .Y(n_476) );
INVxp67_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
BUFx8_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_481), .Y(n_486) );
AND2x2_ASAP7_75t_L g843 ( .A(n_481), .B(n_844), .Y(n_843) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx2_ASAP7_75t_L g829 ( .A(n_482), .Y(n_829) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx12f_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
XNOR2x1_ASAP7_75t_L g830 ( .A(n_487), .B(n_831), .Y(n_830) );
OR2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_705), .Y(n_487) );
NAND3xp33_ASAP7_75t_SL g488 ( .A(n_489), .B(n_608), .C(n_667), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_505), .B1(n_595), .B2(n_601), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OR2x2_ASAP7_75t_L g664 ( .A(n_491), .B(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_491), .B(n_582), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_491), .B(n_628), .Y(n_775) );
AND2x2_ASAP7_75t_L g781 ( .A(n_491), .B(n_607), .Y(n_781) );
INVxp67_ASAP7_75t_L g786 ( .A(n_491), .Y(n_786) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g599 ( .A(n_492), .Y(n_599) );
AOI21x1_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_494), .B(n_504), .Y(n_492) );
INVx4_ASAP7_75t_L g528 ( .A(n_501), .Y(n_528) );
OAI21xp5_ASAP7_75t_SL g505 ( .A1(n_506), .A2(n_557), .B(n_568), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_536), .Y(n_507) );
INVx1_ASAP7_75t_L g702 ( .A(n_508), .Y(n_702) );
AND2x2_ASAP7_75t_L g731 ( .A(n_508), .B(n_693), .Y(n_731) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_523), .Y(n_508) );
AND2x2_ASAP7_75t_L g625 ( .A(n_509), .B(n_546), .Y(n_625) );
INVx1_ASAP7_75t_L g680 ( .A(n_509), .Y(n_680) );
AND2x2_ASAP7_75t_L g730 ( .A(n_509), .B(n_545), .Y(n_730) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g605 ( .A(n_510), .B(n_545), .Y(n_605) );
AND2x4_ASAP7_75t_L g749 ( .A(n_510), .B(n_546), .Y(n_749) );
AOI21x1_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_517), .B(n_521), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_515), .B(n_550), .Y(n_549) );
OAI21xp33_ASAP7_75t_SL g585 ( .A1(n_520), .A2(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
BUFx2_ASAP7_75t_L g674 ( .A(n_523), .Y(n_674) );
AND2x2_ASAP7_75t_L g743 ( .A(n_523), .B(n_546), .Y(n_743) );
AND2x2_ASAP7_75t_L g750 ( .A(n_523), .B(n_576), .Y(n_750) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g572 ( .A(n_524), .Y(n_572) );
BUFx3_ASAP7_75t_L g607 ( .A(n_524), .Y(n_607) );
AND2x2_ASAP7_75t_L g618 ( .A(n_524), .B(n_604), .Y(n_618) );
AND2x2_ASAP7_75t_L g681 ( .A(n_524), .B(n_537), .Y(n_681) );
AND2x2_ASAP7_75t_L g686 ( .A(n_524), .B(n_546), .Y(n_686) );
NAND2x1p5_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
OAI21x1_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_531), .B(n_534), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_536), .B(n_692), .Y(n_794) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_545), .Y(n_536) );
INVx2_ASAP7_75t_L g576 ( .A(n_537), .Y(n_576) );
OR2x2_ASAP7_75t_L g579 ( .A(n_537), .B(n_546), .Y(n_579) );
INVx2_ASAP7_75t_L g604 ( .A(n_537), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_537), .B(n_574), .Y(n_620) );
AND2x2_ASAP7_75t_L g693 ( .A(n_537), .B(n_546), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_541), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g555 ( .A(n_542), .Y(n_555) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g621 ( .A(n_546), .Y(n_621) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_551), .B(n_555), .Y(n_547) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_558), .B(n_656), .Y(n_802) );
BUFx3_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g614 ( .A(n_559), .Y(n_614) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g594 ( .A(n_560), .Y(n_594) );
AND2x2_ASAP7_75t_L g600 ( .A(n_560), .B(n_582), .Y(n_600) );
INVx1_ASAP7_75t_L g648 ( .A(n_560), .Y(n_648) );
OR2x2_ASAP7_75t_L g653 ( .A(n_560), .B(n_632), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_560), .B(n_632), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_560), .B(n_631), .Y(n_734) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_560), .B(n_599), .Y(n_738) );
OAI21xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_577), .B(n_580), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
OR2x2_ASAP7_75t_L g578 ( .A(n_571), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g729 ( .A(n_571), .B(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_L g759 ( .A(n_571), .B(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_572), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g727 ( .A(n_572), .Y(n_727) );
OR2x2_ASAP7_75t_L g640 ( .A(n_573), .B(n_641), .Y(n_640) );
INVxp33_ASAP7_75t_L g758 ( .A(n_573), .Y(n_758) );
OR2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
INVx2_ASAP7_75t_L g662 ( .A(n_574), .Y(n_662) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g616 ( .A(n_576), .Y(n_616) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OAI221xp5_ASAP7_75t_SL g724 ( .A1(n_578), .A2(n_649), .B1(n_654), .B2(n_725), .C(n_728), .Y(n_724) );
OR2x2_ASAP7_75t_L g711 ( .A(n_579), .B(n_662), .Y(n_711) );
INVx2_ASAP7_75t_L g760 ( .A(n_579), .Y(n_760) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g660 ( .A(n_581), .Y(n_660) );
OR2x2_ASAP7_75t_L g663 ( .A(n_581), .B(n_664), .Y(n_663) );
INVxp67_ASAP7_75t_SL g704 ( .A(n_581), .Y(n_704) );
OR2x2_ASAP7_75t_L g717 ( .A(n_581), .B(n_718), .Y(n_717) );
OR2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_594), .Y(n_581) );
NAND2x1p5_ASAP7_75t_SL g613 ( .A(n_582), .B(n_598), .Y(n_613) );
INVx3_ASAP7_75t_L g628 ( .A(n_582), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_582), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g651 ( .A(n_582), .Y(n_651) );
AND2x2_ASAP7_75t_L g732 ( .A(n_582), .B(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g739 ( .A(n_582), .B(n_646), .Y(n_739) );
AND2x4_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
OAI21xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_590), .B(n_593), .Y(n_584) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_600), .Y(n_595) );
AND2x2_ASAP7_75t_L g791 ( .A(n_596), .B(n_650), .Y(n_791) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g695 ( .A(n_598), .B(n_665), .Y(n_695) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g630 ( .A(n_599), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g656 ( .A(n_599), .B(n_632), .Y(n_656) );
AND2x4_ASAP7_75t_L g753 ( .A(n_600), .B(n_723), .Y(n_753) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_606), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_605), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g672 ( .A(n_605), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_606), .B(n_693), .Y(n_777) );
AND2x2_ASAP7_75t_L g784 ( .A(n_606), .B(n_744), .Y(n_784) );
INVx3_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
BUFx2_ASAP7_75t_L g709 ( .A(n_607), .Y(n_709) );
AOI321xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_622), .A3(n_638), .B1(n_639), .B2(n_642), .C(n_657), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_610), .B(n_619), .Y(n_609) );
AOI21xp33_ASAP7_75t_SL g610 ( .A1(n_611), .A2(n_615), .B(n_617), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OAI21xp33_ASAP7_75t_L g622 ( .A1(n_612), .A2(n_623), .B(n_626), .Y(n_622) );
OR2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
OR2x2_ASAP7_75t_L g721 ( .A(n_613), .B(n_653), .Y(n_721) );
INVx1_ASAP7_75t_L g713 ( .A(n_614), .Y(n_713) );
INVx2_ASAP7_75t_L g698 ( .A(n_615), .Y(n_698) );
OAI32xp33_ASAP7_75t_L g801 ( .A1(n_615), .A2(n_763), .A3(n_774), .B1(n_802), .B2(n_803), .Y(n_801) );
INVx1_ASAP7_75t_L g716 ( .A(n_616), .Y(n_716) );
INVx1_ASAP7_75t_L g666 ( .A(n_617), .Y(n_666) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x4_ASAP7_75t_SL g754 ( .A(n_618), .B(n_661), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_619), .B(n_623), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_619), .A2(n_695), .B1(n_756), .B2(n_777), .Y(n_776) );
OR2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
INVx1_ASAP7_75t_L g744 ( .A(n_620), .Y(n_744) );
INVx1_ASAP7_75t_L g641 ( .A(n_621), .Y(n_641) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
BUFx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g726 ( .A(n_625), .Y(n_726) );
NAND4xp25_ASAP7_75t_L g642 ( .A(n_626), .B(n_643), .C(n_649), .D(n_654), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
INVxp67_ASAP7_75t_L g668 ( .A(n_627), .Y(n_668) );
AND2x2_ASAP7_75t_L g747 ( .A(n_627), .B(n_656), .Y(n_747) );
OR2x2_ASAP7_75t_L g756 ( .A(n_627), .B(n_630), .Y(n_756) );
AND2x2_ASAP7_75t_L g780 ( .A(n_627), .B(n_652), .Y(n_780) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g694 ( .A(n_628), .B(n_695), .Y(n_694) );
AND2x4_ASAP7_75t_L g701 ( .A(n_628), .B(n_648), .Y(n_701) );
INVx1_ASAP7_75t_L g765 ( .A(n_629), .Y(n_765) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g673 ( .A(n_630), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g723 ( .A(n_630), .Y(n_723) );
INVx1_ASAP7_75t_L g665 ( .A(n_631), .Y(n_665) );
INVx2_ASAP7_75t_SL g631 ( .A(n_632), .Y(n_631) );
BUFx2_ASAP7_75t_L g646 ( .A(n_632), .Y(n_646) );
INVx3_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
AND2x4_ASAP7_75t_L g659 ( .A(n_645), .B(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g700 ( .A(n_645), .Y(n_700) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_647), .Y(n_764) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AND2x4_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
AND2x2_ASAP7_75t_L g655 ( .A(n_651), .B(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx2_ASAP7_75t_L g741 ( .A(n_653), .Y(n_741) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g718 ( .A(n_656), .Y(n_718) );
AND2x2_ASAP7_75t_L g761 ( .A(n_656), .B(n_701), .Y(n_761) );
O2A1O1Ixp33_ASAP7_75t_SL g657 ( .A1(n_658), .A2(n_661), .B(n_663), .C(n_666), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g772 ( .A(n_661), .B(n_750), .Y(n_772) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g676 ( .A(n_664), .Y(n_676) );
AOI211xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B(n_682), .C(n_696), .Y(n_667) );
OAI21xp33_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_673), .B(n_675), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AOI21xp5_ASAP7_75t_L g778 ( .A1(n_671), .A2(n_779), .B(n_782), .Y(n_778) );
INVx3_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g692 ( .A(n_674), .Y(n_692) );
AND2x2_ASAP7_75t_L g752 ( .A(n_674), .B(n_749), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_679), .B(n_681), .Y(n_678) );
INVx1_ASAP7_75t_L g771 ( .A(n_679), .Y(n_771) );
AND2x2_ASAP7_75t_L g797 ( .A(n_679), .B(n_760), .Y(n_797) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g685 ( .A(n_680), .Y(n_685) );
INVx2_ASAP7_75t_L g736 ( .A(n_681), .Y(n_736) );
NAND2x1_ASAP7_75t_L g770 ( .A(n_681), .B(n_771), .Y(n_770) );
AOI33xp33_ASAP7_75t_L g788 ( .A1(n_681), .A2(n_701), .A3(n_739), .B1(n_749), .B2(n_781), .B3(n_863), .Y(n_788) );
OAI22xp33_ASAP7_75t_SL g682 ( .A1(n_683), .A2(n_687), .B1(n_690), .B2(n_694), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
AND2x2_ASAP7_75t_L g715 ( .A(n_686), .B(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_687), .B(n_774), .Y(n_773) );
OR2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
OR2x2_ASAP7_75t_L g800 ( .A(n_689), .B(n_734), .Y(n_800) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
OAI22xp33_ASAP7_75t_SL g696 ( .A1(n_697), .A2(n_699), .B1(n_702), .B2(n_703), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_700), .B(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_700), .B(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g722 ( .A(n_701), .B(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g787 ( .A(n_701), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_766), .Y(n_705) );
NOR4xp25_ASAP7_75t_L g706 ( .A(n_707), .B(n_724), .C(n_745), .D(n_762), .Y(n_706) );
OAI221xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_712), .B1(n_714), .B2(n_717), .C(n_719), .Y(n_707) );
O2A1O1Ixp33_ASAP7_75t_SL g762 ( .A1(n_708), .A2(n_763), .B(n_764), .C(n_765), .Y(n_762) );
NAND2x1_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g795 ( .A(n_711), .Y(n_795) );
INVx2_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
OAI21xp5_ASAP7_75t_L g719 ( .A1(n_715), .A2(n_720), .B(n_722), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
OR2x6_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
O2A1O1Ixp33_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_731), .B(n_732), .C(n_735), .Y(n_728) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OR2x2_ASAP7_75t_L g774 ( .A(n_734), .B(n_775), .Y(n_774) );
INVxp67_ASAP7_75t_SL g798 ( .A(n_734), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_737), .B1(n_740), .B2(n_742), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
OAI211xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_748), .B(n_751), .C(n_757), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
AOI221xp5_ASAP7_75t_L g796 ( .A1(n_749), .A2(n_797), .B1(n_798), .B2(n_799), .C(n_801), .Y(n_796) );
INVx3_ASAP7_75t_L g804 ( .A(n_749), .Y(n_804) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_753), .B1(n_754), .B2(n_755), .Y(n_751) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
OAI21xp33_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_759), .B(n_761), .Y(n_757) );
INVx1_ASAP7_75t_L g763 ( .A(n_760), .Y(n_763) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_789), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_768), .B(n_778), .Y(n_767) );
O2A1O1Ixp33_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_772), .B(n_773), .C(n_776), .Y(n_768) );
INVx2_ASAP7_75t_SL g769 ( .A(n_770), .Y(n_769) );
NOR3xp33_ASAP7_75t_L g792 ( .A(n_772), .B(n_793), .C(n_795), .Y(n_792) );
AND2x2_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
OAI21xp5_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_785), .B(n_788), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
OR2x2_ASAP7_75t_L g785 ( .A(n_786), .B(n_787), .Y(n_785) );
OAI21xp5_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_792), .B(n_796), .Y(n_789) );
INVx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx2_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx3_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx6_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
AND2x6_ASAP7_75t_SL g812 ( .A(n_813), .B(n_815), .Y(n_812) );
BUFx3_ASAP7_75t_L g821 ( .A(n_813), .Y(n_821) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
NOR2xp33_ASAP7_75t_L g841 ( .A(n_814), .B(n_842), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_816), .B(n_818), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
NOR2x1_ASAP7_75t_L g844 ( .A(n_817), .B(n_819), .Y(n_844) );
AND3x2_ASAP7_75t_L g826 ( .A(n_818), .B(n_827), .C(n_829), .Y(n_826) );
AND2x6_ASAP7_75t_SL g847 ( .A(n_818), .B(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
BUFx2_ASAP7_75t_L g855 ( .A(n_819), .Y(n_855) );
OAI21xp33_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_822), .B(n_837), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_823), .B(n_830), .Y(n_822) );
INVx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx3_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx4_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
NOR2x1p5_ASAP7_75t_L g856 ( .A(n_827), .B(n_857), .Y(n_856) );
HB1xp67_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g849 ( .A(n_828), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_829), .B(n_858), .Y(n_857) );
AOI22x1_ASAP7_75t_L g831 ( .A1(n_832), .A2(n_833), .B1(n_834), .B2(n_835), .Y(n_831) );
CKINVDCx5p33_ASAP7_75t_R g832 ( .A(n_833), .Y(n_832) );
CKINVDCx5p33_ASAP7_75t_R g835 ( .A(n_836), .Y(n_835) );
INVx3_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx6_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
BUFx10_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
NOR2xp33_ASAP7_75t_L g845 ( .A(n_846), .B(n_850), .Y(n_845) );
INVx3_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
BUFx6f_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx6_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx6_ASAP7_75t_L g861 ( .A(n_853), .Y(n_861) );
NAND2x2_ASAP7_75t_L g853 ( .A(n_854), .B(n_856), .Y(n_853) );
CKINVDCx5p33_ASAP7_75t_R g854 ( .A(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
endmodule