module fake_jpeg_5950_n_103 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_103);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_103;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_5),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

OR2x2_ASAP7_75t_SL g19 ( 
.A(n_8),
.B(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_26),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_0),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_13),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_30),
.A2(n_17),
.B1(n_21),
.B2(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_33),
.Y(n_34)
);

AND2x2_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_19),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_45),
.B(n_11),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_26),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_24),
.A2(n_17),
.B1(n_23),
.B2(n_12),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_28),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_30),
.A2(n_23),
.B1(n_12),
.B2(n_20),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_3),
.C(n_4),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_SL g45 ( 
.A(n_25),
.B(n_21),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_28),
.A2(n_15),
.B1(n_11),
.B2(n_13),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_32),
.B1(n_29),
.B2(n_31),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_47),
.A2(n_48),
.B(n_59),
.Y(n_69)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_51),
.Y(n_63)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_0),
.Y(n_53)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_54),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_1),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_56),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_33),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_57),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_35),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_33),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_58),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_66),
.A2(n_49),
.B1(n_56),
.B2(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_74),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_SL g75 ( 
.A1(n_72),
.A2(n_49),
.B(n_37),
.C(n_61),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_75),
.A2(n_78),
.B(n_79),
.Y(n_83)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_76),
.A2(n_77),
.B(n_80),
.Y(n_84)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_64),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_59),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g86 ( 
.A1(n_81),
.A2(n_45),
.B(n_72),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_65),
.C(n_59),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_39),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_86),
.B(n_81),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_62),
.Y(n_88)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_70),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_91),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_92),
.Y(n_93)
);

AOI322xp5_ASAP7_75t_SL g91 ( 
.A1(n_86),
.A2(n_75),
.A3(n_73),
.B1(n_70),
.B2(n_67),
.C1(n_60),
.C2(n_4),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_85),
.C(n_87),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_97),
.B(n_98),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_94),
.B(n_82),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_91),
.C(n_39),
.Y(n_98)
);

AOI21x1_ASAP7_75t_SL g100 ( 
.A1(n_98),
.A2(n_7),
.B(n_9),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_100),
.A2(n_10),
.B(n_99),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_74),
.C(n_58),
.Y(n_103)
);


endmodule