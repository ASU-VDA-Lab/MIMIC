module fake_jpeg_5584_n_63 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_63);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_63;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_38;
wire n_36;
wire n_62;
wire n_56;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_3),
.B(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_7),
.B(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_27),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_43),
.Y(n_50)
);

CKINVDCx12_ASAP7_75t_R g43 ( 
.A(n_39),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_45),
.B(n_1),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_46),
.A2(n_34),
.B1(n_4),
.B2(n_5),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_51),
.B(n_6),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_55),
.B1(n_52),
.B2(n_18),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_8),
.C(n_11),
.Y(n_54)
);

MAJx2_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_13),
.C(n_14),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_48),
.B(n_12),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_57),
.B(n_15),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_58),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_23),
.Y(n_60)
);

NAND3xp33_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_25),
.C(n_28),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_29),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_30),
.Y(n_63)
);


endmodule