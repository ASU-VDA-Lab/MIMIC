module fake_netlist_1_9915_n_643 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_643);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_643;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g74 ( .A(n_35), .Y(n_74) );
CKINVDCx5p33_ASAP7_75t_R g75 ( .A(n_37), .Y(n_75) );
INVx2_ASAP7_75t_L g76 ( .A(n_38), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_20), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_0), .Y(n_78) );
NOR2xp67_ASAP7_75t_L g79 ( .A(n_24), .B(n_5), .Y(n_79) );
INVx1_ASAP7_75t_SL g80 ( .A(n_45), .Y(n_80) );
INVxp67_ASAP7_75t_SL g81 ( .A(n_3), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_13), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_23), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_36), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_62), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_59), .Y(n_86) );
INVx2_ASAP7_75t_SL g87 ( .A(n_70), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_28), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_26), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_67), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_21), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_68), .Y(n_92) );
INVxp67_ASAP7_75t_L g93 ( .A(n_72), .Y(n_93) );
BUFx3_ASAP7_75t_L g94 ( .A(n_42), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_51), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_53), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_61), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_33), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_44), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_18), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_57), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_9), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_2), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_22), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_50), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_10), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_34), .Y(n_107) );
INVxp33_ASAP7_75t_L g108 ( .A(n_48), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_56), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_15), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_7), .Y(n_112) );
INVxp67_ASAP7_75t_L g113 ( .A(n_7), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_1), .Y(n_114) );
BUFx3_ASAP7_75t_L g115 ( .A(n_40), .Y(n_115) );
XOR2xp5_ASAP7_75t_L g116 ( .A(n_54), .B(n_66), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_60), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_1), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_74), .Y(n_119) );
OR2x2_ASAP7_75t_SL g120 ( .A(n_82), .B(n_0), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_118), .B(n_87), .Y(n_121) );
AND2x2_ASAP7_75t_L g122 ( .A(n_118), .B(n_3), .Y(n_122) );
AND2x2_ASAP7_75t_L g123 ( .A(n_108), .B(n_4), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_74), .Y(n_124) );
CKINVDCx16_ASAP7_75t_R g125 ( .A(n_116), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_94), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_94), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_102), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_77), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_77), .Y(n_130) );
BUFx2_ASAP7_75t_L g131 ( .A(n_102), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_83), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_76), .Y(n_133) );
NAND2xp33_ASAP7_75t_L g134 ( .A(n_75), .B(n_73), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_83), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_84), .Y(n_136) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_113), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_75), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_76), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_82), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_84), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_89), .Y(n_142) );
AOI22xp5_ASAP7_75t_SL g143 ( .A1(n_116), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_87), .B(n_6), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_78), .B(n_8), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_89), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_112), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_92), .B(n_8), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_90), .Y(n_149) );
OAI22xp5_ASAP7_75t_L g150 ( .A1(n_112), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_88), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g152 ( .A(n_88), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_114), .B(n_11), .Y(n_153) );
OR2x6_ASAP7_75t_L g154 ( .A(n_114), .B(n_12), .Y(n_154) );
BUFx8_ASAP7_75t_L g155 ( .A(n_90), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_91), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_91), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_96), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_121), .B(n_109), .Y(n_159) );
BUFx2_ASAP7_75t_L g160 ( .A(n_131), .Y(n_160) );
INVx4_ASAP7_75t_SL g161 ( .A(n_154), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_147), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_147), .Y(n_163) );
NAND3xp33_ASAP7_75t_L g164 ( .A(n_123), .B(n_103), .C(n_106), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_131), .B(n_97), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_147), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_126), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_126), .Y(n_168) );
BUFx10_ASAP7_75t_L g169 ( .A(n_138), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_119), .B(n_97), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_138), .B(n_151), .Y(n_171) );
INVx4_ASAP7_75t_L g172 ( .A(n_154), .Y(n_172) );
HB1xp67_ASAP7_75t_L g173 ( .A(n_128), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_122), .B(n_111), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_133), .Y(n_175) );
AO21x2_ASAP7_75t_L g176 ( .A1(n_145), .A2(n_96), .B(n_95), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_126), .Y(n_177) );
HB1xp67_ASAP7_75t_SL g178 ( .A(n_155), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_122), .B(n_117), .Y(n_179) );
INVxp67_ASAP7_75t_L g180 ( .A(n_128), .Y(n_180) );
INVx2_ASAP7_75t_SL g181 ( .A(n_123), .Y(n_181) );
INVx4_ASAP7_75t_L g182 ( .A(n_154), .Y(n_182) );
BUFx4f_ASAP7_75t_L g183 ( .A(n_154), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_126), .Y(n_184) );
OR2x6_ASAP7_75t_L g185 ( .A(n_150), .B(n_79), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_119), .B(n_117), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_124), .B(n_110), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_126), .Y(n_188) );
INVx4_ASAP7_75t_L g189 ( .A(n_127), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_127), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_127), .Y(n_191) );
BUFx10_ASAP7_75t_L g192 ( .A(n_151), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_152), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_137), .B(n_124), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_129), .B(n_110), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_129), .B(n_93), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_130), .B(n_99), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_133), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_130), .B(n_81), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_155), .A2(n_86), .B1(n_85), .B2(n_105), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_153), .Y(n_201) );
INVx2_ASAP7_75t_SL g202 ( .A(n_132), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_155), .B(n_107), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_132), .B(n_104), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_127), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_127), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_139), .Y(n_207) );
INVx3_ASAP7_75t_L g208 ( .A(n_139), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_146), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_135), .B(n_101), .Y(n_210) );
AO22x1_ASAP7_75t_L g211 ( .A1(n_153), .A2(n_100), .B1(n_98), .B2(n_115), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_146), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_162), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_170), .B(n_158), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_178), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_162), .Y(n_216) );
NOR2xp33_ASAP7_75t_R g217 ( .A(n_183), .B(n_125), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_181), .A2(n_144), .B1(n_148), .B2(n_158), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_186), .B(n_149), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_161), .B(n_183), .Y(n_220) );
NOR2x2_ASAP7_75t_L g221 ( .A(n_185), .B(n_183), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_181), .A2(n_142), .B1(n_135), .B2(n_149), .Y(n_222) );
INVx2_ASAP7_75t_SL g223 ( .A(n_161), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_199), .A2(n_142), .B1(n_141), .B2(n_136), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_162), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_201), .A2(n_136), .B(n_141), .C(n_157), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_187), .B(n_157), .Y(n_227) );
INVx3_ASAP7_75t_L g228 ( .A(n_172), .Y(n_228) );
NAND3xp33_ASAP7_75t_SL g229 ( .A(n_193), .B(n_80), .C(n_156), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_195), .B(n_156), .Y(n_230) );
INVx5_ASAP7_75t_L g231 ( .A(n_172), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_163), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_179), .B(n_140), .Y(n_233) );
BUFx2_ASAP7_75t_L g234 ( .A(n_160), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_193), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_179), .B(n_140), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_168), .Y(n_237) );
AOI22x1_ASAP7_75t_L g238 ( .A1(n_189), .A2(n_140), .B1(n_143), .B2(n_134), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_166), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_175), .Y(n_240) );
AND2x2_ASAP7_75t_L g241 ( .A(n_160), .B(n_115), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_159), .B(n_12), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_168), .Y(n_243) );
AOI22xp33_ASAP7_75t_SL g244 ( .A1(n_172), .A2(n_120), .B1(n_14), .B2(n_15), .Y(n_244) );
AO22x1_ASAP7_75t_L g245 ( .A1(n_182), .A2(n_120), .B1(n_14), .B2(n_13), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_175), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_159), .B(n_16), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_198), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_184), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_184), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_169), .Y(n_251) );
INVx3_ASAP7_75t_L g252 ( .A(n_182), .Y(n_252) );
NOR2xp67_ASAP7_75t_L g253 ( .A(n_182), .B(n_17), .Y(n_253) );
INVx3_ASAP7_75t_L g254 ( .A(n_208), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_198), .Y(n_255) );
AND2x4_ASAP7_75t_L g256 ( .A(n_161), .B(n_19), .Y(n_256) );
INVx1_ASAP7_75t_SL g257 ( .A(n_165), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_208), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_159), .B(n_25), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g260 ( .A1(n_194), .A2(n_27), .B1(n_29), .B2(n_30), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_188), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_161), .B(n_31), .Y(n_262) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_194), .Y(n_263) );
OAI22xp33_ASAP7_75t_L g264 ( .A1(n_185), .A2(n_32), .B1(n_39), .B2(n_41), .Y(n_264) );
INVx2_ASAP7_75t_SL g265 ( .A(n_199), .Y(n_265) );
INVx2_ASAP7_75t_SL g266 ( .A(n_169), .Y(n_266) );
BUFx3_ASAP7_75t_L g267 ( .A(n_199), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_202), .B(n_43), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_202), .B(n_46), .Y(n_269) );
INVx3_ASAP7_75t_L g270 ( .A(n_208), .Y(n_270) );
OR2x2_ASAP7_75t_L g271 ( .A(n_234), .B(n_173), .Y(n_271) );
NAND2x1_ASAP7_75t_L g272 ( .A(n_256), .B(n_212), .Y(n_272) );
AND2x4_ASAP7_75t_L g273 ( .A(n_266), .B(n_203), .Y(n_273) );
INVx1_ASAP7_75t_SL g274 ( .A(n_263), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_231), .B(n_192), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_214), .A2(n_176), .B(n_211), .Y(n_276) );
AOI21xp33_ASAP7_75t_L g277 ( .A1(n_247), .A2(n_176), .B(n_197), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_225), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_224), .B(n_257), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_225), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_265), .B(n_176), .Y(n_281) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_256), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_267), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_215), .Y(n_284) );
BUFx3_ASAP7_75t_L g285 ( .A(n_215), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_225), .Y(n_286) );
AND2x4_ASAP7_75t_L g287 ( .A(n_267), .B(n_265), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_219), .A2(n_211), .B(n_210), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g289 ( .A1(n_251), .A2(n_180), .B1(n_171), .B2(n_200), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_232), .Y(n_290) );
INVx2_ASAP7_75t_SL g291 ( .A(n_251), .Y(n_291) );
BUFx3_ASAP7_75t_L g292 ( .A(n_235), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_239), .Y(n_293) );
O2A1O1Ixp33_ASAP7_75t_L g294 ( .A1(n_226), .A2(n_204), .B(n_209), .C(n_212), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_254), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_235), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_227), .A2(n_196), .B(n_164), .Y(n_297) );
INVx5_ASAP7_75t_L g298 ( .A(n_256), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_222), .B(n_174), .Y(n_299) );
INVx4_ASAP7_75t_L g300 ( .A(n_231), .Y(n_300) );
AO32x2_ASAP7_75t_L g301 ( .A1(n_226), .A2(n_189), .A3(n_167), .B1(n_190), .B2(n_177), .Y(n_301) );
BUFx2_ASAP7_75t_L g302 ( .A(n_217), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_233), .Y(n_303) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_223), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_231), .B(n_192), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_230), .A2(n_174), .B(n_209), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_238), .A2(n_174), .B1(n_185), .B2(n_207), .Y(n_307) );
O2A1O1Ixp33_ASAP7_75t_L g308 ( .A1(n_236), .A2(n_185), .B(n_207), .C(n_205), .Y(n_308) );
INVxp67_ASAP7_75t_SL g309 ( .A(n_223), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_240), .B(n_192), .Y(n_310) );
BUFx12f_ASAP7_75t_L g311 ( .A(n_231), .Y(n_311) );
OAI22xp5_ASAP7_75t_SL g312 ( .A1(n_244), .A2(n_169), .B1(n_189), .B2(n_191), .Y(n_312) );
OR2x2_ASAP7_75t_L g313 ( .A(n_241), .B(n_205), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_259), .A2(n_206), .B(n_191), .Y(n_314) );
INVxp67_ASAP7_75t_SL g315 ( .A(n_228), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_290), .Y(n_316) );
AO21x2_ASAP7_75t_L g317 ( .A1(n_277), .A2(n_268), .B(n_262), .Y(n_317) );
INVx4_ASAP7_75t_L g318 ( .A(n_311), .Y(n_318) );
OAI21x1_ASAP7_75t_L g319 ( .A1(n_314), .A2(n_268), .B(n_262), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_277), .A2(n_220), .B(n_216), .Y(n_320) );
OA21x2_ASAP7_75t_L g321 ( .A1(n_314), .A2(n_269), .B(n_260), .Y(n_321) );
OAI21x1_ASAP7_75t_L g322 ( .A1(n_308), .A2(n_253), .B(n_220), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_299), .B(n_242), .Y(n_323) );
AOI22xp33_ASAP7_75t_SL g324 ( .A1(n_292), .A2(n_221), .B1(n_231), .B2(n_228), .Y(n_324) );
AND2x2_ASAP7_75t_SL g325 ( .A(n_282), .B(n_221), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_293), .Y(n_326) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_298), .A2(n_218), .B1(n_255), .B2(n_248), .Y(n_327) );
AO21x2_ASAP7_75t_L g328 ( .A1(n_276), .A2(n_264), .B(n_206), .Y(n_328) );
OAI21x1_ASAP7_75t_L g329 ( .A1(n_308), .A2(n_246), .B(n_261), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_303), .Y(n_330) );
AOI22xp33_ASAP7_75t_SL g331 ( .A1(n_302), .A2(n_228), .B1(n_252), .B2(n_245), .Y(n_331) );
OAI21x1_ASAP7_75t_L g332 ( .A1(n_272), .A2(n_261), .B(n_250), .Y(n_332) );
OAI21x1_ASAP7_75t_L g333 ( .A1(n_276), .A2(n_250), .B(n_249), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_279), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_281), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_299), .B(n_252), .Y(n_336) );
OR2x6_ASAP7_75t_L g337 ( .A(n_282), .B(n_252), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_274), .A2(n_279), .B1(n_271), .B2(n_287), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_296), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_287), .A2(n_229), .B1(n_254), .B2(n_270), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_310), .B(n_270), .Y(n_341) );
INVx5_ASAP7_75t_L g342 ( .A(n_300), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_298), .A2(n_270), .B1(n_254), .B2(n_258), .Y(n_343) );
AND2x4_ASAP7_75t_L g344 ( .A(n_273), .B(n_213), .Y(n_344) );
OAI21xp33_ASAP7_75t_L g345 ( .A1(n_331), .A2(n_307), .B(n_289), .Y(n_345) );
INVx3_ASAP7_75t_L g346 ( .A(n_342), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g347 ( .A1(n_330), .A2(n_338), .B1(n_316), .B2(n_326), .C(n_297), .Y(n_347) );
A2O1A1Ixp33_ASAP7_75t_L g348 ( .A1(n_335), .A2(n_288), .B(n_306), .C(n_297), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_330), .B(n_291), .Y(n_349) );
OA21x2_ASAP7_75t_L g350 ( .A1(n_329), .A2(n_281), .B(n_306), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_326), .Y(n_351) );
INVx4_ASAP7_75t_L g352 ( .A(n_318), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_335), .A2(n_298), .B1(n_282), .B2(n_310), .Y(n_353) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_325), .B(n_298), .Y(n_354) );
OAI222xp33_ASAP7_75t_L g355 ( .A1(n_324), .A2(n_288), .B1(n_300), .B2(n_275), .C1(n_305), .C2(n_294), .Y(n_355) );
OAI222xp33_ASAP7_75t_L g356 ( .A1(n_334), .A2(n_294), .B1(n_283), .B2(n_313), .C1(n_273), .C2(n_312), .Y(n_356) );
AOI22xp33_ASAP7_75t_SL g357 ( .A1(n_325), .A2(n_284), .B1(n_285), .B2(n_315), .Y(n_357) );
AOI21xp5_ASAP7_75t_L g358 ( .A1(n_320), .A2(n_286), .B(n_280), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_323), .B(n_295), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_344), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_344), .Y(n_361) );
OAI222xp33_ASAP7_75t_L g362 ( .A1(n_327), .A2(n_278), .B1(n_301), .B2(n_309), .C1(n_188), .C2(n_243), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_339), .A2(n_304), .B1(n_237), .B2(n_249), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_340), .A2(n_304), .B1(n_243), .B2(n_237), .C(n_190), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_339), .B(n_304), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g366 ( .A1(n_317), .A2(n_190), .B(n_177), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_344), .Y(n_367) );
AO21x2_ASAP7_75t_L g368 ( .A1(n_329), .A2(n_301), .B(n_190), .Y(n_368) );
AOI221xp5_ASAP7_75t_L g369 ( .A1(n_336), .A2(n_190), .B1(n_177), .B2(n_167), .C(n_301), .Y(n_369) );
AOI221xp5_ASAP7_75t_L g370 ( .A1(n_318), .A2(n_177), .B1(n_167), .B2(n_52), .C(n_55), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_347), .B(n_328), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_351), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_350), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_348), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_350), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_368), .Y(n_376) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_346), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_359), .B(n_342), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_360), .B(n_361), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_345), .A2(n_328), .B1(n_341), .B2(n_318), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_368), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_359), .B(n_342), .Y(n_382) );
BUFx2_ASAP7_75t_L g383 ( .A(n_346), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_367), .B(n_342), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_349), .B(n_328), .Y(n_385) );
INVxp67_ASAP7_75t_L g386 ( .A(n_365), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_357), .B(n_342), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_354), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_357), .B(n_333), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_353), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_358), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_363), .B(n_333), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_369), .B(n_332), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_366), .B(n_317), .Y(n_394) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_352), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_362), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_362), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_364), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_352), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_355), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_370), .A2(n_337), .B1(n_321), .B2(n_317), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_356), .B(n_322), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_355), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_385), .B(n_322), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_385), .B(n_337), .Y(n_405) );
BUFx3_ASAP7_75t_L g406 ( .A(n_383), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_372), .B(n_319), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_372), .B(n_319), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_373), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_374), .B(n_321), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_373), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_374), .B(n_321), .Y(n_412) );
BUFx2_ASAP7_75t_L g413 ( .A(n_375), .Y(n_413) );
BUFx2_ASAP7_75t_L g414 ( .A(n_375), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_376), .Y(n_415) );
AOI211x1_ASAP7_75t_SL g416 ( .A1(n_399), .A2(n_343), .B(n_356), .C(n_177), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_386), .B(n_337), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_383), .B(n_337), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_378), .Y(n_419) );
OAI221xp5_ASAP7_75t_L g420 ( .A1(n_380), .A2(n_167), .B1(n_332), .B2(n_58), .C(n_63), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_371), .A2(n_167), .B1(n_49), .B2(n_64), .C(n_65), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_389), .B(n_47), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_400), .B(n_69), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_389), .B(n_71), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_378), .Y(n_425) );
OAI31xp33_ASAP7_75t_L g426 ( .A1(n_395), .A2(n_382), .A3(n_387), .B(n_399), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_387), .B(n_392), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_376), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_381), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_382), .B(n_403), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_381), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_391), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_379), .B(n_384), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_400), .B(n_403), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_391), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_371), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_394), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_392), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_396), .B(n_397), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_396), .B(n_397), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_379), .B(n_393), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_393), .B(n_402), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_394), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_388), .B(n_384), .Y(n_444) );
INVx5_ASAP7_75t_SL g445 ( .A(n_377), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_402), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_377), .B(n_388), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_377), .Y(n_448) );
AND2x4_ASAP7_75t_L g449 ( .A(n_377), .B(n_390), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_377), .B(n_390), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_442), .B(n_398), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_428), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_433), .B(n_398), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_442), .B(n_401), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_441), .B(n_438), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_409), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_439), .B(n_440), .Y(n_457) );
AOI221xp5_ASAP7_75t_L g458 ( .A1(n_446), .A2(n_436), .B1(n_438), .B2(n_417), .C(n_444), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_435), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_413), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_435), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_428), .Y(n_462) );
INVx1_ASAP7_75t_SL g463 ( .A(n_413), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_432), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_406), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_441), .B(n_427), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_427), .B(n_407), .Y(n_467) );
NOR2x1_ASAP7_75t_L g468 ( .A(n_406), .B(n_418), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_428), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_432), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_432), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_431), .Y(n_472) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_449), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_431), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_419), .B(n_425), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_431), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_439), .B(n_440), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_427), .B(n_407), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_411), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_434), .B(n_430), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_427), .B(n_408), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_408), .B(n_430), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_446), .B(n_414), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_411), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_415), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_409), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_409), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_414), .B(n_450), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g489 ( .A1(n_423), .A2(n_434), .B(n_412), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_415), .Y(n_490) );
INVxp67_ASAP7_75t_L g491 ( .A(n_406), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_429), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_429), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_444), .B(n_405), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_450), .B(n_436), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_410), .B(n_412), .Y(n_496) );
INVx4_ASAP7_75t_L g497 ( .A(n_418), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_410), .B(n_443), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_405), .B(n_422), .Y(n_499) );
NOR2xp33_ASAP7_75t_SL g500 ( .A(n_426), .B(n_424), .Y(n_500) );
INVx3_ASAP7_75t_R g501 ( .A(n_449), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_426), .A2(n_424), .B1(n_422), .B2(n_421), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_437), .B(n_443), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_437), .B(n_443), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_437), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_482), .B(n_455), .Y(n_506) );
AND3x2_ASAP7_75t_L g507 ( .A(n_500), .B(n_447), .C(n_448), .Y(n_507) );
NAND2xp33_ASAP7_75t_L g508 ( .A(n_502), .B(n_448), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_459), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_505), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_451), .B(n_404), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_451), .B(n_404), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_505), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_455), .B(n_447), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_482), .B(n_478), .Y(n_515) );
INVxp67_ASAP7_75t_L g516 ( .A(n_465), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_480), .B(n_449), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_505), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_457), .B(n_449), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_459), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_457), .B(n_423), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_453), .B(n_420), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_467), .B(n_445), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_467), .B(n_445), .Y(n_524) );
NOR2xp67_ASAP7_75t_SL g525 ( .A(n_497), .B(n_445), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_461), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_454), .A2(n_416), .B1(n_445), .B2(n_500), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_477), .B(n_416), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_478), .B(n_445), .Y(n_529) );
AND2x4_ASAP7_75t_L g530 ( .A(n_495), .B(n_483), .Y(n_530) );
NAND2x1p5_ASAP7_75t_L g531 ( .A(n_468), .B(n_497), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_486), .Y(n_532) );
CKINVDCx16_ASAP7_75t_R g533 ( .A(n_475), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_494), .B(n_458), .Y(n_534) );
NOR2x1p5_ASAP7_75t_L g535 ( .A(n_497), .B(n_466), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_461), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_481), .B(n_466), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_496), .B(n_495), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_504), .B(n_496), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_498), .B(n_454), .Y(n_540) );
O2A1O1Ixp33_ASAP7_75t_L g541 ( .A1(n_491), .A2(n_489), .B(n_503), .C(n_460), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_498), .B(n_483), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_481), .B(n_488), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_488), .B(n_489), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_479), .Y(n_545) );
AND2x2_ASAP7_75t_SL g546 ( .A(n_497), .B(n_499), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_479), .B(n_484), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_468), .A2(n_463), .B1(n_460), .B2(n_484), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_485), .Y(n_549) );
INVxp67_ASAP7_75t_L g550 ( .A(n_463), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_485), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_492), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_504), .B(n_456), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_456), .B(n_490), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_539), .Y(n_555) );
INVxp67_ASAP7_75t_L g556 ( .A(n_528), .Y(n_556) );
AOI211xp5_ASAP7_75t_L g557 ( .A1(n_508), .A2(n_473), .B(n_493), .C(n_492), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_539), .Y(n_558) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_550), .Y(n_559) );
AOI21xp33_ASAP7_75t_SL g560 ( .A1(n_533), .A2(n_501), .B(n_493), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_514), .Y(n_561) );
OA21x2_ASAP7_75t_L g562 ( .A1(n_527), .A2(n_452), .B(n_476), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_547), .Y(n_563) );
OAI21xp5_ASAP7_75t_L g564 ( .A1(n_541), .A2(n_490), .B(n_464), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_546), .B(n_456), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_515), .B(n_473), .Y(n_566) );
INVx2_ASAP7_75t_SL g567 ( .A(n_535), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_546), .B(n_456), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_506), .B(n_464), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_548), .B(n_490), .Y(n_570) );
NAND2x1_ASAP7_75t_L g571 ( .A(n_525), .B(n_471), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_509), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_520), .Y(n_573) );
OAI21xp33_ASAP7_75t_L g574 ( .A1(n_544), .A2(n_471), .B(n_470), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_515), .B(n_473), .Y(n_575) );
OAI211xp5_ASAP7_75t_SL g576 ( .A1(n_508), .A2(n_470), .B(n_462), .C(n_469), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_532), .Y(n_577) );
OAI21xp5_ASAP7_75t_L g578 ( .A1(n_522), .A2(n_487), .B(n_486), .Y(n_578) );
NOR2xp33_ASAP7_75t_SL g579 ( .A(n_531), .B(n_487), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_506), .B(n_473), .Y(n_580) );
OAI22xp33_ASAP7_75t_L g581 ( .A1(n_531), .A2(n_473), .B1(n_487), .B2(n_486), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_534), .B(n_452), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_526), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_532), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_536), .Y(n_585) );
A2O1A1Ixp33_ASAP7_75t_L g586 ( .A1(n_522), .A2(n_501), .B(n_462), .C(n_469), .Y(n_586) );
INVx1_ASAP7_75t_SL g587 ( .A(n_523), .Y(n_587) );
OAI21xp33_ASAP7_75t_L g588 ( .A1(n_544), .A2(n_452), .B(n_462), .Y(n_588) );
XNOR2x1_ASAP7_75t_L g589 ( .A(n_587), .B(n_537), .Y(n_589) );
INVxp67_ASAP7_75t_L g590 ( .A(n_582), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_569), .Y(n_591) );
OAI21xp5_ASAP7_75t_L g592 ( .A1(n_556), .A2(n_516), .B(n_527), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_577), .Y(n_593) );
INVxp67_ASAP7_75t_SL g594 ( .A(n_570), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_555), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_558), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_561), .B(n_538), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_572), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_578), .B(n_540), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_574), .A2(n_521), .B1(n_512), .B2(n_511), .C(n_553), .Y(n_600) );
INVx3_ASAP7_75t_L g601 ( .A(n_571), .Y(n_601) );
AOI32xp33_ASAP7_75t_L g602 ( .A1(n_567), .A2(n_537), .A3(n_530), .B1(n_543), .B2(n_524), .Y(n_602) );
O2A1O1Ixp33_ASAP7_75t_L g603 ( .A1(n_565), .A2(n_552), .B(n_551), .C(n_549), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_580), .B(n_543), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_580), .B(n_530), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_563), .B(n_530), .Y(n_606) );
AOI221xp5_ASAP7_75t_L g607 ( .A1(n_588), .A2(n_553), .B1(n_542), .B2(n_545), .C(n_554), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_573), .Y(n_608) );
O2A1O1Ixp5_ASAP7_75t_SL g609 ( .A1(n_570), .A2(n_507), .B(n_519), .C(n_517), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_590), .B(n_559), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_589), .Y(n_611) );
AOI322xp5_ASAP7_75t_L g612 ( .A1(n_594), .A2(n_567), .A3(n_565), .B1(n_568), .B2(n_575), .C1(n_566), .C2(n_586), .Y(n_612) );
OAI211xp5_ASAP7_75t_L g613 ( .A1(n_592), .A2(n_560), .B(n_568), .C(n_586), .Y(n_613) );
OAI211xp5_ASAP7_75t_L g614 ( .A1(n_602), .A2(n_557), .B(n_564), .C(n_562), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_598), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_608), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_595), .Y(n_617) );
NOR2x1p5_ASAP7_75t_L g618 ( .A(n_601), .B(n_575), .Y(n_618) );
OAI21xp5_ASAP7_75t_L g619 ( .A1(n_609), .A2(n_576), .B(n_581), .Y(n_619) );
OAI21xp5_ASAP7_75t_L g620 ( .A1(n_603), .A2(n_579), .B(n_562), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_590), .A2(n_562), .B1(n_523), .B2(n_529), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_599), .A2(n_529), .B1(n_524), .B2(n_583), .Y(n_622) );
O2A1O1Ixp33_ASAP7_75t_L g623 ( .A1(n_611), .A2(n_601), .B(n_603), .C(n_596), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_613), .A2(n_600), .B1(n_607), .B2(n_591), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_618), .A2(n_607), .B1(n_600), .B2(n_606), .Y(n_625) );
O2A1O1Ixp33_ASAP7_75t_L g626 ( .A1(n_619), .A2(n_597), .B(n_593), .C(n_585), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_610), .A2(n_473), .B1(n_605), .B2(n_604), .Y(n_627) );
AOI211xp5_ASAP7_75t_L g628 ( .A1(n_614), .A2(n_554), .B(n_584), .C(n_577), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_622), .A2(n_584), .B1(n_510), .B2(n_513), .Y(n_629) );
XNOR2x1_ASAP7_75t_L g630 ( .A(n_624), .B(n_620), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_629), .Y(n_631) );
BUFx2_ASAP7_75t_L g632 ( .A(n_625), .Y(n_632) );
O2A1O1Ixp33_ASAP7_75t_L g633 ( .A1(n_623), .A2(n_621), .B(n_616), .C(n_615), .Y(n_633) );
AND2x4_ASAP7_75t_L g634 ( .A(n_632), .B(n_627), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_631), .Y(n_635) );
O2A1O1Ixp33_ASAP7_75t_L g636 ( .A1(n_633), .A2(n_626), .B(n_628), .C(n_630), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_634), .A2(n_621), .B1(n_617), .B2(n_612), .Y(n_637) );
A2O1A1Ixp33_ASAP7_75t_L g638 ( .A1(n_636), .A2(n_510), .B(n_513), .C(n_518), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_637), .A2(n_634), .B1(n_635), .B2(n_518), .Y(n_639) );
XNOR2x1_ASAP7_75t_L g640 ( .A(n_639), .B(n_638), .Y(n_640) );
AOI22xp33_ASAP7_75t_SL g641 ( .A1(n_640), .A2(n_469), .B1(n_472), .B2(n_474), .Y(n_641) );
AO221x2_ASAP7_75t_L g642 ( .A1(n_641), .A2(n_472), .B1(n_474), .B2(n_476), .C(n_635), .Y(n_642) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_642), .A2(n_476), .B(n_472), .Y(n_643) );
endmodule