module real_aes_8940_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_717;
wire n_359;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g455 ( .A1(n_0), .A2(n_155), .B(n_456), .C(n_459), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_1), .B(n_450), .Y(n_460) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_2), .B(n_89), .C(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g117 ( .A(n_2), .Y(n_117) );
INVx1_ASAP7_75t_L g153 ( .A(n_3), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_4), .B(n_156), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_5), .A2(n_445), .B(n_518), .Y(n_517) );
AO21x2_ASAP7_75t_L g525 ( .A1(n_6), .A2(n_178), .B(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_7), .A2(n_38), .B1(n_143), .B2(n_201), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_8), .A2(n_9), .B1(n_707), .B2(n_708), .Y(n_706) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_8), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_9), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_10), .B(n_178), .Y(n_186) );
AND2x6_ASAP7_75t_L g158 ( .A(n_11), .B(n_159), .Y(n_158) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_12), .A2(n_158), .B(n_436), .C(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_13), .B(n_106), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g118 ( .A(n_13), .B(n_39), .Y(n_118) );
INVx1_ASAP7_75t_L g137 ( .A(n_14), .Y(n_137) );
INVx1_ASAP7_75t_L g134 ( .A(n_15), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_16), .B(n_139), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_17), .B(n_156), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_18), .B(n_130), .Y(n_188) );
AO32x2_ASAP7_75t_L g239 ( .A1(n_19), .A2(n_129), .A3(n_172), .B1(n_178), .B2(n_240), .Y(n_239) );
OAI22xp5_ASAP7_75t_SL g727 ( .A1(n_20), .A2(n_30), .B1(n_120), .B2(n_728), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_20), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_21), .B(n_143), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_22), .B(n_130), .Y(n_160) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_23), .A2(n_56), .B1(n_143), .B2(n_201), .Y(n_242) );
AOI22xp33_ASAP7_75t_SL g203 ( .A1(n_24), .A2(n_81), .B1(n_139), .B2(n_143), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_25), .B(n_143), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g466 ( .A1(n_26), .A2(n_172), .B(n_436), .C(n_467), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_27), .A2(n_172), .B(n_436), .C(n_529), .Y(n_528) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_28), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_29), .B(n_174), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g119 ( .A1(n_30), .A2(n_120), .B1(n_121), .B2(n_122), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_30), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_31), .A2(n_445), .B(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_32), .B(n_174), .Y(n_216) );
INVx2_ASAP7_75t_L g141 ( .A(n_33), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_34), .A2(n_442), .B(n_485), .C(n_486), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_35), .B(n_143), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_36), .B(n_174), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_37), .B(n_223), .Y(n_530) );
INVx1_ASAP7_75t_L g106 ( .A(n_39), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_40), .B(n_465), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_41), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_42), .A2(n_103), .B1(n_111), .B2(n_736), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_43), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_44), .B(n_156), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_45), .B(n_445), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_46), .A2(n_442), .B(n_485), .C(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_47), .B(n_143), .Y(n_181) );
INVx1_ASAP7_75t_L g457 ( .A(n_48), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_49), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_50), .A2(n_90), .B1(n_201), .B2(n_202), .Y(n_200) );
INVx1_ASAP7_75t_L g510 ( .A(n_51), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_52), .B(n_143), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_53), .B(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_54), .B(n_445), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_55), .B(n_151), .Y(n_185) );
AOI22xp33_ASAP7_75t_SL g192 ( .A1(n_57), .A2(n_61), .B1(n_139), .B2(n_143), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_58), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_59), .B(n_143), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_60), .B(n_143), .Y(n_220) );
INVx1_ASAP7_75t_L g159 ( .A(n_62), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_63), .B(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_64), .B(n_450), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_65), .A2(n_145), .B(n_151), .C(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_66), .B(n_143), .Y(n_154) );
INVx1_ASAP7_75t_L g133 ( .A(n_67), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_68), .Y(n_720) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_69), .B(n_156), .Y(n_488) );
AO32x2_ASAP7_75t_L g198 ( .A1(n_70), .A2(n_172), .A3(n_178), .B1(n_199), .B2(n_204), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_71), .B(n_157), .Y(n_501) );
INVx1_ASAP7_75t_L g168 ( .A(n_72), .Y(n_168) );
INVx1_ASAP7_75t_L g211 ( .A(n_73), .Y(n_211) );
CKINVDCx16_ASAP7_75t_R g453 ( .A(n_74), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_75), .B(n_469), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g435 ( .A1(n_76), .A2(n_436), .B(n_438), .C(n_442), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_77), .B(n_139), .Y(n_212) );
CKINVDCx16_ASAP7_75t_R g519 ( .A(n_78), .Y(n_519) );
INVx1_ASAP7_75t_L g110 ( .A(n_79), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_80), .B(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_82), .B(n_201), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_83), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_84), .B(n_139), .Y(n_215) );
INVx2_ASAP7_75t_L g131 ( .A(n_85), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_86), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_87), .B(n_171), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_88), .B(n_139), .Y(n_182) );
OR2x2_ASAP7_75t_L g115 ( .A(n_89), .B(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g427 ( .A(n_89), .Y(n_427) );
OR2x2_ASAP7_75t_L g724 ( .A(n_89), .B(n_716), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_91), .A2(n_101), .B1(n_139), .B2(n_140), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_92), .B(n_445), .Y(n_483) );
INVx1_ASAP7_75t_L g487 ( .A(n_93), .Y(n_487) );
INVxp67_ASAP7_75t_L g522 ( .A(n_94), .Y(n_522) );
XNOR2xp5_ASAP7_75t_L g725 ( .A(n_95), .B(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_96), .B(n_139), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_97), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g439 ( .A(n_98), .Y(n_439) );
INVx1_ASAP7_75t_L g497 ( .A(n_99), .Y(n_497) );
AND2x2_ASAP7_75t_L g512 ( .A(n_100), .B(n_174), .Y(n_512) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
CKINVDCx6p67_ASAP7_75t_R g737 ( .A(n_104), .Y(n_737) );
OR2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_107), .Y(n_104) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
AO221x1_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_718), .B1(n_721), .B2(n_730), .C(n_732), .Y(n_111) );
OAI222xp33_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_706), .B1(n_709), .B2(n_713), .C1(n_714), .C2(n_717), .Y(n_112) );
AOI22xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_119), .B1(n_425), .B2(n_428), .Y(n_113) );
INVx2_ASAP7_75t_L g711 ( .A(n_114), .Y(n_711) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OR2x2_ASAP7_75t_L g426 ( .A(n_116), .B(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g716 ( .A(n_116), .Y(n_716) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
OAI22xp5_ASAP7_75t_SL g710 ( .A1(n_119), .A2(n_428), .B1(n_711), .B2(n_712), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_121), .A2(n_122), .B1(n_727), .B2(n_729), .Y(n_726) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OR5x1_ASAP7_75t_L g122 ( .A(n_123), .B(n_316), .C(n_374), .D(n_410), .E(n_417), .Y(n_122) );
NAND3xp33_ASAP7_75t_SL g123 ( .A(n_124), .B(n_262), .C(n_286), .Y(n_123) );
AOI221xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_194), .B1(n_228), .B2(n_233), .C(n_243), .Y(n_124) );
OAI21xp5_ASAP7_75t_SL g396 ( .A1(n_125), .A2(n_397), .B(n_399), .Y(n_396) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_175), .Y(n_125) );
NAND2x1p5_ASAP7_75t_L g386 ( .A(n_126), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_161), .Y(n_126) );
INVx2_ASAP7_75t_L g232 ( .A(n_127), .Y(n_232) );
AND2x2_ASAP7_75t_L g245 ( .A(n_127), .B(n_177), .Y(n_245) );
AND2x2_ASAP7_75t_L g299 ( .A(n_127), .B(n_176), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_127), .B(n_162), .Y(n_314) );
OA21x2_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_135), .B(n_160), .Y(n_127) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_128), .A2(n_163), .B(n_173), .Y(n_162) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_129), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_130), .Y(n_178) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
AND2x2_ASAP7_75t_SL g174 ( .A(n_131), .B(n_132), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
OAI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_149), .B(n_158), .Y(n_135) );
O2A1O1Ixp33_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_138), .B(n_142), .C(n_145), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_138), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_138), .A2(n_530), .B(n_531), .Y(n_529) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g144 ( .A(n_141), .Y(n_144) );
INVx1_ASAP7_75t_L g152 ( .A(n_141), .Y(n_152) );
INVx3_ASAP7_75t_L g210 ( .A(n_143), .Y(n_210) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_143), .Y(n_441) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g201 ( .A(n_144), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_144), .Y(n_202) );
AND2x6_ASAP7_75t_L g436 ( .A(n_144), .B(n_437), .Y(n_436) );
O2A1O1Ixp33_ASAP7_75t_L g438 ( .A1(n_145), .A2(n_439), .B(n_440), .C(n_441), .Y(n_438) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_146), .A2(n_214), .B(n_215), .Y(n_213) );
INVx4_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g469 ( .A(n_147), .Y(n_469) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx3_ASAP7_75t_L g157 ( .A(n_148), .Y(n_157) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_148), .Y(n_171) );
INVx1_ASAP7_75t_L g223 ( .A(n_148), .Y(n_223) );
INVx1_ASAP7_75t_L g437 ( .A(n_148), .Y(n_437) );
AND2x2_ASAP7_75t_L g446 ( .A(n_148), .B(n_152), .Y(n_446) );
O2A1O1Ixp33_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_153), .B(n_154), .C(n_155), .Y(n_149) );
O2A1O1Ixp5_ASAP7_75t_L g167 ( .A1(n_150), .A2(n_168), .B(n_169), .C(n_170), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_150), .A2(n_468), .B(n_470), .Y(n_467) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_155), .A2(n_184), .B(n_185), .Y(n_183) );
OAI22xp5_ASAP7_75t_L g190 ( .A1(n_155), .A2(n_171), .B1(n_191), .B2(n_192), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_155), .A2(n_171), .B1(n_241), .B2(n_242), .Y(n_240) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_156), .A2(n_165), .B(n_166), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_156), .A2(n_181), .B(n_182), .Y(n_180) );
O2A1O1Ixp5_ASAP7_75t_SL g209 ( .A1(n_156), .A2(n_210), .B(n_211), .C(n_212), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_156), .B(n_522), .Y(n_521) );
INVx5_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
OAI22xp5_ASAP7_75t_SL g199 ( .A1(n_157), .A2(n_171), .B1(n_200), .B2(n_203), .Y(n_199) );
BUFx3_ASAP7_75t_L g172 ( .A(n_158), .Y(n_172) );
OAI21xp5_ASAP7_75t_L g179 ( .A1(n_158), .A2(n_180), .B(n_183), .Y(n_179) );
OAI21xp5_ASAP7_75t_L g208 ( .A1(n_158), .A2(n_209), .B(n_213), .Y(n_208) );
OAI21xp5_ASAP7_75t_L g218 ( .A1(n_158), .A2(n_219), .B(n_224), .Y(n_218) );
INVx4_ASAP7_75t_SL g443 ( .A(n_158), .Y(n_443) );
AND2x4_ASAP7_75t_L g445 ( .A(n_158), .B(n_446), .Y(n_445) );
NAND2x1p5_ASAP7_75t_L g498 ( .A(n_158), .B(n_446), .Y(n_498) );
AND2x2_ASAP7_75t_L g332 ( .A(n_161), .B(n_273), .Y(n_332) );
AND2x2_ASAP7_75t_L g365 ( .A(n_161), .B(n_177), .Y(n_365) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
OR2x2_ASAP7_75t_L g272 ( .A(n_162), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g285 ( .A(n_162), .B(n_177), .Y(n_285) );
AND2x2_ASAP7_75t_L g292 ( .A(n_162), .B(n_273), .Y(n_292) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_162), .Y(n_301) );
AND2x2_ASAP7_75t_L g308 ( .A(n_162), .B(n_176), .Y(n_308) );
INVx1_ASAP7_75t_L g339 ( .A(n_162), .Y(n_339) );
OAI21xp5_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_167), .B(n_172), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_170), .A2(n_225), .B(n_226), .Y(n_224) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx4_ASAP7_75t_L g458 ( .A(n_171), .Y(n_458) );
NAND3xp33_ASAP7_75t_L g189 ( .A(n_172), .B(n_190), .C(n_193), .Y(n_189) );
INVx2_ASAP7_75t_L g204 ( .A(n_174), .Y(n_204) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_174), .A2(n_208), .B(n_216), .Y(n_207) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_174), .A2(n_218), .B(n_227), .Y(n_217) );
INVx1_ASAP7_75t_L g475 ( .A(n_174), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_174), .A2(n_483), .B(n_484), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_174), .A2(n_507), .B(n_508), .Y(n_506) );
INVx1_ASAP7_75t_L g315 ( .A(n_175), .Y(n_315) );
AND2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_187), .Y(n_175) );
INVx2_ASAP7_75t_L g271 ( .A(n_176), .Y(n_271) );
AND2x2_ASAP7_75t_L g293 ( .A(n_176), .B(n_232), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_176), .B(n_339), .Y(n_344) );
INVx3_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_177), .B(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g416 ( .A(n_177), .B(n_380), .Y(n_416) );
OA21x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_186), .Y(n_177) );
INVx4_ASAP7_75t_L g193 ( .A(n_178), .Y(n_193) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_178), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_178), .A2(n_527), .B(n_528), .Y(n_526) );
INVx2_ASAP7_75t_L g230 ( .A(n_187), .Y(n_230) );
INVx3_ASAP7_75t_L g331 ( .A(n_187), .Y(n_331) );
OR2x2_ASAP7_75t_L g361 ( .A(n_187), .B(n_362), .Y(n_361) );
NOR2x1_ASAP7_75t_L g387 ( .A(n_187), .B(n_271), .Y(n_387) );
AND2x4_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
INVx1_ASAP7_75t_L g274 ( .A(n_188), .Y(n_274) );
AO21x1_ASAP7_75t_L g273 ( .A1(n_190), .A2(n_193), .B(n_274), .Y(n_273) );
AO21x2_ASAP7_75t_L g433 ( .A1(n_193), .A2(n_434), .B(n_447), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_193), .B(n_448), .Y(n_447) );
INVx3_ASAP7_75t_L g450 ( .A(n_193), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_193), .B(n_491), .Y(n_490) );
AO21x2_ASAP7_75t_L g495 ( .A1(n_193), .A2(n_496), .B(n_503), .Y(n_495) );
AOI33xp33_ASAP7_75t_L g407 ( .A1(n_194), .A2(n_245), .A3(n_259), .B1(n_331), .B2(n_408), .B3(n_409), .Y(n_407) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
OR2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_205), .Y(n_195) );
OR2x2_ASAP7_75t_L g260 ( .A(n_196), .B(n_261), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_196), .B(n_257), .Y(n_319) );
OR2x2_ASAP7_75t_L g372 ( .A(n_196), .B(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g298 ( .A(n_197), .B(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g323 ( .A(n_197), .B(n_205), .Y(n_323) );
AND2x2_ASAP7_75t_L g390 ( .A(n_197), .B(n_235), .Y(n_390) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_197), .A2(n_290), .B(n_416), .Y(n_415) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g237 ( .A(n_198), .Y(n_237) );
INVx1_ASAP7_75t_L g250 ( .A(n_198), .Y(n_250) );
AND2x2_ASAP7_75t_L g269 ( .A(n_198), .B(n_239), .Y(n_269) );
AND2x2_ASAP7_75t_L g318 ( .A(n_198), .B(n_238), .Y(n_318) );
INVx2_ASAP7_75t_L g459 ( .A(n_202), .Y(n_459) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_202), .Y(n_489) );
INVx1_ASAP7_75t_L g472 ( .A(n_204), .Y(n_472) );
INVx2_ASAP7_75t_SL g360 ( .A(n_205), .Y(n_360) );
OR2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_217), .Y(n_205) );
INVx2_ASAP7_75t_L g280 ( .A(n_206), .Y(n_280) );
INVx1_ASAP7_75t_L g411 ( .A(n_206), .Y(n_411) );
AND2x2_ASAP7_75t_L g424 ( .A(n_206), .B(n_305), .Y(n_424) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g251 ( .A(n_207), .Y(n_251) );
OR2x2_ASAP7_75t_L g257 ( .A(n_207), .B(n_258), .Y(n_257) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_207), .Y(n_268) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_217), .Y(n_235) );
AND2x2_ASAP7_75t_L g252 ( .A(n_217), .B(n_238), .Y(n_252) );
INVx1_ASAP7_75t_L g258 ( .A(n_217), .Y(n_258) );
INVx1_ASAP7_75t_L g265 ( .A(n_217), .Y(n_265) );
AND2x2_ASAP7_75t_L g290 ( .A(n_217), .B(n_239), .Y(n_290) );
INVx2_ASAP7_75t_L g306 ( .A(n_217), .Y(n_306) );
AND2x2_ASAP7_75t_L g399 ( .A(n_217), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_217), .B(n_280), .Y(n_420) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_222), .Y(n_219) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_SL g228 ( .A(n_229), .Y(n_228) );
OR2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
INVx2_ASAP7_75t_L g254 ( .A(n_230), .Y(n_254) );
INVx1_ASAP7_75t_L g283 ( .A(n_230), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_230), .B(n_314), .Y(n_380) );
INVx1_ASAP7_75t_SL g340 ( .A(n_231), .Y(n_340) );
INVx2_ASAP7_75t_L g261 ( .A(n_232), .Y(n_261) );
AND2x2_ASAP7_75t_L g330 ( .A(n_232), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g346 ( .A(n_232), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_236), .Y(n_233) );
INVx1_ASAP7_75t_L g408 ( .A(n_234), .Y(n_408) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g263 ( .A(n_236), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g366 ( .A(n_236), .B(n_356), .Y(n_366) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_236), .A2(n_377), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
AND2x2_ASAP7_75t_L g279 ( .A(n_237), .B(n_280), .Y(n_279) );
BUFx2_ASAP7_75t_L g304 ( .A(n_237), .Y(n_304) );
INVx1_ASAP7_75t_L g328 ( .A(n_237), .Y(n_328) );
OR2x2_ASAP7_75t_L g392 ( .A(n_238), .B(n_251), .Y(n_392) );
NOR2xp67_ASAP7_75t_L g400 ( .A(n_238), .B(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g305 ( .A(n_239), .B(n_306), .Y(n_305) );
BUFx2_ASAP7_75t_L g312 ( .A(n_239), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_246), .B1(n_253), .B2(n_255), .Y(n_243) );
OR2x2_ASAP7_75t_L g322 ( .A(n_244), .B(n_272), .Y(n_322) );
INVx1_ASAP7_75t_SL g244 ( .A(n_245), .Y(n_244) );
AOI222xp33_ASAP7_75t_L g363 ( .A1(n_245), .A2(n_364), .B1(n_366), .B2(n_367), .C1(n_368), .C2(n_371), .Y(n_363) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_252), .Y(n_247) );
INVx1_ASAP7_75t_SL g248 ( .A(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g310 ( .A(n_249), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
AND2x2_ASAP7_75t_SL g264 ( .A(n_251), .B(n_265), .Y(n_264) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_251), .Y(n_335) );
AND2x2_ASAP7_75t_L g383 ( .A(n_251), .B(n_252), .Y(n_383) );
INVx1_ASAP7_75t_L g401 ( .A(n_251), .Y(n_401) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g367 ( .A(n_254), .B(n_293), .Y(n_367) );
AND2x2_ASAP7_75t_L g409 ( .A(n_254), .B(n_285), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_259), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_256), .B(n_304), .Y(n_391) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_257), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g284 ( .A(n_261), .B(n_285), .Y(n_284) );
INVx3_ASAP7_75t_L g352 ( .A(n_261), .Y(n_352) );
O2A1O1Ixp33_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_266), .B(n_270), .C(n_275), .Y(n_262) );
INVxp67_ASAP7_75t_L g276 ( .A(n_263), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_264), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_264), .B(n_311), .Y(n_406) );
BUFx3_ASAP7_75t_L g370 ( .A(n_265), .Y(n_370) );
INVx1_ASAP7_75t_L g277 ( .A(n_266), .Y(n_277) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_269), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g296 ( .A(n_268), .B(n_290), .Y(n_296) );
INVx1_ASAP7_75t_SL g336 ( .A(n_269), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
INVx1_ASAP7_75t_L g326 ( .A(n_271), .Y(n_326) );
AND2x2_ASAP7_75t_L g349 ( .A(n_271), .B(n_332), .Y(n_349) );
INVx1_ASAP7_75t_SL g320 ( .A(n_272), .Y(n_320) );
INVx1_ASAP7_75t_L g347 ( .A(n_273), .Y(n_347) );
AOI31xp33_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_277), .A3(n_278), .B(n_281), .Y(n_275) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g368 ( .A(n_279), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g342 ( .A(n_280), .Y(n_342) );
BUFx2_ASAP7_75t_L g356 ( .A(n_280), .Y(n_356) );
AND2x2_ASAP7_75t_L g384 ( .A(n_280), .B(n_305), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_SL g357 ( .A(n_284), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_285), .B(n_352), .Y(n_398) );
AND2x2_ASAP7_75t_L g405 ( .A(n_285), .B(n_331), .Y(n_405) );
AOI211xp5_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_291), .B(n_294), .C(n_309), .Y(n_286) );
INVxp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AOI221xp5_ASAP7_75t_L g317 ( .A1(n_291), .A2(n_318), .B1(n_319), .B2(n_320), .C(n_321), .Y(n_317) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
AND2x2_ASAP7_75t_L g325 ( .A(n_292), .B(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g362 ( .A(n_293), .Y(n_362) );
OAI32xp33_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_297), .A3(n_300), .B1(n_302), .B2(n_307), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
O2A1O1Ixp33_ASAP7_75t_L g348 ( .A1(n_296), .A2(n_349), .B(n_350), .C(n_353), .Y(n_348) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
OAI21xp5_ASAP7_75t_SL g412 ( .A1(n_304), .A2(n_413), .B(n_414), .Y(n_412) );
INVx1_ASAP7_75t_L g373 ( .A(n_305), .Y(n_373) );
INVxp67_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_310), .B(n_313), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_311), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g359 ( .A(n_311), .B(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g376 ( .A(n_313), .Y(n_376) );
OR2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
NAND4xp25_ASAP7_75t_SL g316 ( .A(n_317), .B(n_329), .C(n_348), .D(n_363), .Y(n_316) );
AND2x2_ASAP7_75t_L g355 ( .A(n_318), .B(n_356), .Y(n_355) );
AND2x4_ASAP7_75t_L g377 ( .A(n_318), .B(n_370), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_320), .B(n_352), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_323), .B1(n_324), .B2(n_327), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_322), .A2(n_373), .B1(n_404), .B2(n_406), .Y(n_403) );
O2A1O1Ixp33_ASAP7_75t_L g410 ( .A1(n_322), .A2(n_411), .B(n_412), .C(n_415), .Y(n_410) );
INVx2_ASAP7_75t_L g381 ( .A(n_323), .Y(n_381) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AOI222xp33_ASAP7_75t_L g375 ( .A1(n_325), .A2(n_359), .B1(n_376), .B2(n_377), .C1(n_378), .C2(n_381), .Y(n_375) );
O2A1O1Ixp33_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_332), .B(n_333), .C(n_337), .Y(n_329) );
INVx1_ASAP7_75t_L g395 ( .A(n_330), .Y(n_395) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OAI22xp33_ASAP7_75t_L g337 ( .A1(n_334), .A2(n_338), .B1(n_341), .B2(n_343), .Y(n_337) );
OR2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g364 ( .A(n_346), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g422 ( .A(n_349), .Y(n_422) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OAI22xp33_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_357), .B1(n_358), .B2(n_361), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_356), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g413 ( .A(n_361), .Y(n_413) );
INVx1_ASAP7_75t_L g394 ( .A(n_365), .Y(n_394) );
CKINVDCx16_ASAP7_75t_R g421 ( .A(n_367), .Y(n_421) );
INVxp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND5xp2_ASAP7_75t_L g374 ( .A(n_375), .B(n_382), .C(n_396), .D(n_402), .E(n_407), .Y(n_374) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
O2A1O1Ixp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_384), .B(n_385), .C(n_388), .Y(n_382) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AOI31xp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_391), .A3(n_392), .B(n_393), .Y(n_388) );
INVx1_ASAP7_75t_L g414 ( .A(n_390), .Y(n_414) );
OR2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OAI222xp33_ASAP7_75t_L g417 ( .A1(n_404), .A2(n_406), .B1(n_418), .B2(n_421), .C1(n_422), .C2(n_423), .Y(n_417) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g712 ( .A(n_425), .Y(n_712) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NOR2x2_ASAP7_75t_L g715 ( .A(n_427), .B(n_716), .Y(n_715) );
OR3x1_ASAP7_75t_L g428 ( .A(n_429), .B(n_614), .C(n_663), .Y(n_428) );
NAND5xp2_ASAP7_75t_L g429 ( .A(n_430), .B(n_548), .C(n_577), .D(n_585), .E(n_600), .Y(n_429) );
O2A1O1Ixp33_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_476), .B(n_492), .C(n_532), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_432), .B(n_461), .Y(n_431) );
AND2x2_ASAP7_75t_L g543 ( .A(n_432), .B(n_540), .Y(n_543) );
AND2x2_ASAP7_75t_L g576 ( .A(n_432), .B(n_462), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_432), .B(n_480), .Y(n_669) );
AND2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_449), .Y(n_432) );
INVx2_ASAP7_75t_L g479 ( .A(n_433), .Y(n_479) );
BUFx2_ASAP7_75t_L g643 ( .A(n_433), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_444), .Y(n_434) );
INVx5_ASAP7_75t_L g454 ( .A(n_436), .Y(n_454) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
O2A1O1Ixp33_ASAP7_75t_SL g452 ( .A1(n_443), .A2(n_453), .B(n_454), .C(n_455), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_L g518 ( .A1(n_443), .A2(n_454), .B(n_519), .C(n_520), .Y(n_518) );
BUFx2_ASAP7_75t_L g465 ( .A(n_445), .Y(n_465) );
AND2x2_ASAP7_75t_L g461 ( .A(n_449), .B(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g541 ( .A(n_449), .Y(n_541) );
AND2x2_ASAP7_75t_L g627 ( .A(n_449), .B(n_540), .Y(n_627) );
AND2x2_ASAP7_75t_L g682 ( .A(n_449), .B(n_479), .Y(n_682) );
OA21x2_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_451), .B(n_460), .Y(n_449) );
INVx2_ASAP7_75t_L g485 ( .A(n_454), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
INVx1_ASAP7_75t_L g599 ( .A(n_461), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_461), .B(n_480), .Y(n_646) );
INVx5_ASAP7_75t_L g540 ( .A(n_462), .Y(n_540) );
AND2x4_ASAP7_75t_L g561 ( .A(n_462), .B(n_541), .Y(n_561) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_462), .Y(n_583) );
AND2x2_ASAP7_75t_L g658 ( .A(n_462), .B(n_643), .Y(n_658) );
AND2x2_ASAP7_75t_L g661 ( .A(n_462), .B(n_481), .Y(n_661) );
OR2x6_ASAP7_75t_L g462 ( .A(n_463), .B(n_473), .Y(n_462) );
AOI21xp5_ASAP7_75t_SL g463 ( .A1(n_464), .A2(n_466), .B(n_472), .Y(n_463) );
INVx2_ASAP7_75t_L g471 ( .A(n_469), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g486 ( .A1(n_471), .A2(n_487), .B(n_488), .C(n_489), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_L g509 ( .A1(n_471), .A2(n_489), .B(n_510), .C(n_511), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_476), .B(n_541), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_476), .B(n_672), .Y(n_671) );
INVx2_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_480), .Y(n_477) );
AND2x2_ASAP7_75t_L g566 ( .A(n_478), .B(n_541), .Y(n_566) );
AND2x2_ASAP7_75t_L g584 ( .A(n_478), .B(n_481), .Y(n_584) );
INVx1_ASAP7_75t_L g604 ( .A(n_478), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_478), .B(n_540), .Y(n_649) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_478), .Y(n_691) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_479), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_480), .B(n_539), .Y(n_538) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_480), .Y(n_593) );
O2A1O1Ixp33_ASAP7_75t_L g596 ( .A1(n_480), .A2(n_536), .B(n_597), .C(n_599), .Y(n_596) );
AND2x2_ASAP7_75t_L g603 ( .A(n_480), .B(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g612 ( .A(n_480), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g616 ( .A(n_480), .B(n_540), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_480), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g631 ( .A(n_480), .B(n_541), .Y(n_631) );
AND2x2_ASAP7_75t_L g681 ( .A(n_480), .B(n_682), .Y(n_681) );
INVx5_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
BUFx2_ASAP7_75t_L g545 ( .A(n_481), .Y(n_545) );
AND2x2_ASAP7_75t_L g586 ( .A(n_481), .B(n_539), .Y(n_586) );
AND2x2_ASAP7_75t_L g598 ( .A(n_481), .B(n_573), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_481), .B(n_627), .Y(n_645) );
OR2x6_ASAP7_75t_L g481 ( .A(n_482), .B(n_490), .Y(n_481) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_513), .Y(n_492) );
INVx1_ASAP7_75t_L g534 ( .A(n_493), .Y(n_534) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_505), .Y(n_493) );
OR2x2_ASAP7_75t_L g536 ( .A(n_494), .B(n_505), .Y(n_536) );
NAND3xp33_ASAP7_75t_L g542 ( .A(n_494), .B(n_543), .C(n_544), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_494), .B(n_515), .Y(n_553) );
OR2x2_ASAP7_75t_L g568 ( .A(n_494), .B(n_556), .Y(n_568) );
AND2x2_ASAP7_75t_L g574 ( .A(n_494), .B(n_524), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_494), .B(n_705), .Y(n_704) );
INVx5_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_495), .B(n_515), .Y(n_571) );
AND2x2_ASAP7_75t_L g610 ( .A(n_495), .B(n_525), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_495), .B(n_524), .Y(n_638) );
OR2x2_ASAP7_75t_L g641 ( .A(n_495), .B(n_524), .Y(n_641) );
OAI21xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B(n_499), .Y(n_496) );
INVx5_ASAP7_75t_SL g556 ( .A(n_505), .Y(n_556) );
OR2x2_ASAP7_75t_L g562 ( .A(n_505), .B(n_514), .Y(n_562) );
AND2x2_ASAP7_75t_L g578 ( .A(n_505), .B(n_579), .Y(n_578) );
AOI321xp33_ASAP7_75t_L g585 ( .A1(n_505), .A2(n_586), .A3(n_587), .B1(n_588), .B2(n_594), .C(n_596), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_505), .B(n_513), .Y(n_595) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_505), .Y(n_608) );
OR2x2_ASAP7_75t_L g655 ( .A(n_505), .B(n_553), .Y(n_655) );
AND2x2_ASAP7_75t_L g677 ( .A(n_505), .B(n_574), .Y(n_677) );
AND2x2_ASAP7_75t_L g696 ( .A(n_505), .B(n_515), .Y(n_696) );
OR2x6_ASAP7_75t_L g505 ( .A(n_506), .B(n_512), .Y(n_505) );
INVx1_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_524), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_515), .B(n_524), .Y(n_537) );
AND2x2_ASAP7_75t_L g546 ( .A(n_515), .B(n_547), .Y(n_546) );
INVx3_ASAP7_75t_L g573 ( .A(n_515), .Y(n_573) );
AND2x2_ASAP7_75t_L g579 ( .A(n_515), .B(n_574), .Y(n_579) );
INVxp67_ASAP7_75t_L g609 ( .A(n_515), .Y(n_609) );
OR2x2_ASAP7_75t_L g651 ( .A(n_515), .B(n_556), .Y(n_651) );
OA21x2_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_517), .B(n_523), .Y(n_515) );
OR2x2_ASAP7_75t_L g533 ( .A(n_524), .B(n_534), .Y(n_533) );
INVx1_ASAP7_75t_SL g547 ( .A(n_524), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_524), .B(n_536), .Y(n_580) );
AND2x2_ASAP7_75t_L g629 ( .A(n_524), .B(n_573), .Y(n_629) );
AND2x2_ASAP7_75t_L g667 ( .A(n_524), .B(n_556), .Y(n_667) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_525), .B(n_556), .Y(n_555) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_535), .B(n_538), .C(n_542), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_533), .A2(n_535), .B1(n_660), .B2(n_662), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_535), .A2(n_558), .B1(n_613), .B2(n_699), .Y(n_698) );
OR2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
INVx1_ASAP7_75t_SL g687 ( .A(n_536), .Y(n_687) );
INVx1_ASAP7_75t_SL g587 ( .A(n_537), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_539), .B(n_559), .Y(n_589) );
AOI222xp33_ASAP7_75t_L g600 ( .A1(n_539), .A2(n_580), .B1(n_587), .B2(n_601), .C1(n_605), .C2(n_611), .Y(n_600) );
AND2x2_ASAP7_75t_L g690 ( .A(n_539), .B(n_691), .Y(n_690) );
AND2x4_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
INVx2_ASAP7_75t_L g565 ( .A(n_540), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_540), .B(n_560), .Y(n_635) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_540), .Y(n_672) );
AND2x2_ASAP7_75t_L g675 ( .A(n_540), .B(n_584), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_540), .B(n_691), .Y(n_701) );
INVx1_ASAP7_75t_L g592 ( .A(n_541), .Y(n_592) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_541), .Y(n_620) );
O2A1O1Ixp33_ASAP7_75t_L g683 ( .A1(n_543), .A2(n_684), .B(n_685), .C(n_688), .Y(n_683) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
NAND3xp33_ASAP7_75t_L g606 ( .A(n_545), .B(n_607), .C(n_610), .Y(n_606) );
OR2x2_ASAP7_75t_L g634 ( .A(n_545), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_545), .B(n_561), .Y(n_662) );
OR2x2_ASAP7_75t_L g567 ( .A(n_547), .B(n_568), .Y(n_567) );
AOI211xp5_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_551), .B(n_557), .C(n_569), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_550), .B(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g656 ( .A(n_551), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_554), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_552), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g570 ( .A(n_555), .B(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_556), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g624 ( .A(n_556), .B(n_574), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_556), .B(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_556), .B(n_573), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_562), .B1(n_563), .B2(n_567), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_559), .B(n_631), .Y(n_630) );
BUFx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_561), .B(n_603), .Y(n_602) );
OAI221xp5_ASAP7_75t_SL g625 ( .A1(n_562), .A2(n_626), .B1(n_628), .B2(n_630), .C(n_632), .Y(n_625) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
AND2x2_ASAP7_75t_L g680 ( .A(n_565), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g693 ( .A(n_565), .B(n_682), .Y(n_693) );
INVx1_ASAP7_75t_L g613 ( .A(n_566), .Y(n_613) );
INVx1_ASAP7_75t_L g684 ( .A(n_567), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_568), .A2(n_651), .B(n_674), .Y(n_673) );
AOI21xp33_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_572), .B(n_575), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OAI21xp5_ASAP7_75t_SL g577 ( .A1(n_578), .A2(n_580), .B(n_581), .Y(n_577) );
INVx1_ASAP7_75t_L g617 ( .A(n_578), .Y(n_617) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_579), .A2(n_665), .B1(n_668), .B2(n_670), .C(n_673), .Y(n_664) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_587), .A2(n_677), .B1(n_678), .B2(n_680), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx1_ASAP7_75t_L g653 ( .A(n_589), .Y(n_653) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NOR2xp67_ASAP7_75t_SL g591 ( .A(n_592), .B(n_593), .Y(n_591) );
AND2x2_ASAP7_75t_L g657 ( .A(n_593), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g622 ( .A(n_598), .Y(n_622) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_603), .B(n_627), .Y(n_679) );
INVxp67_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_609), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g695 ( .A(n_610), .B(n_696), .Y(n_695) );
AND2x4_ASAP7_75t_L g702 ( .A(n_610), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OAI211xp5_ASAP7_75t_SL g614 ( .A1(n_615), .A2(n_617), .B(n_618), .C(n_652), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AOI211xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_621), .B(n_625), .C(n_644), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_SL g705 ( .A(n_629), .Y(n_705) );
AND2x2_ASAP7_75t_L g642 ( .A(n_631), .B(n_643), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_636), .B1(n_640), .B2(n_642), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OR2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
OR2x2_ASAP7_75t_L g650 ( .A(n_638), .B(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g703 ( .A(n_639), .Y(n_703) );
INVxp67_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AOI31xp33_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_646), .A3(n_647), .B(n_650), .Y(n_644) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AOI211xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_654), .B(n_656), .C(n_659), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
CKINVDCx16_ASAP7_75t_R g660 ( .A(n_661), .Y(n_660) );
NAND5xp2_ASAP7_75t_L g663 ( .A(n_664), .B(n_676), .C(n_683), .D(n_697), .E(n_700), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_675), .A2(n_701), .B1(n_702), .B2(n_704), .Y(n_700) );
INVx1_ASAP7_75t_SL g699 ( .A(n_677), .Y(n_699) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AOI21xp33_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_692), .B(n_694), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVxp67_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g713 ( .A(n_706), .Y(n_713) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
BUFx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_SL g731 ( .A(n_719), .Y(n_731) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVxp67_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_725), .Y(n_722) );
BUFx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g735 ( .A(n_724), .Y(n_735) );
INVx1_ASAP7_75t_L g729 ( .A(n_727), .Y(n_729) );
BUFx3_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
INVx1_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_737), .Y(n_736) );
endmodule