module fake_jpeg_29889_n_408 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_408);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_408;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_SL g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_47),
.Y(n_129)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_51),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_17),
.B(n_14),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_52),
.B(n_73),
.Y(n_112)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_54),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_55),
.Y(n_126)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_57),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_58),
.Y(n_147)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_60),
.Y(n_132)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_61),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_62),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_17),
.B(n_13),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_63),
.B(n_74),
.Y(n_138)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx11_ASAP7_75t_L g152 ( 
.A(n_65),
.Y(n_152)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_66),
.Y(n_153)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_20),
.B(n_13),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_68),
.B(n_71),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_20),
.B(n_11),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_SL g140 ( 
.A(n_72),
.B(n_75),
.Y(n_140)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_24),
.B(n_12),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_31),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_80),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_78),
.B(n_79),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_24),
.B(n_9),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_87),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_40),
.B(n_0),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_82),
.B(n_83),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_40),
.B(n_44),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_89),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_37),
.B(n_0),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_91),
.B(n_95),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

BUFx10_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_96),
.B(n_97),
.Y(n_130)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

AND2x4_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_26),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_103),
.B(n_37),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_68),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_105),
.B(n_117),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_71),
.B(n_44),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_108),
.B(n_149),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_79),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_82),
.A2(n_64),
.B1(n_92),
.B2(n_86),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_118),
.A2(n_120),
.B1(n_122),
.B2(n_124),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_50),
.A2(n_66),
.B1(n_67),
.B2(n_26),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_46),
.A2(n_33),
.B1(n_41),
.B2(n_15),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_70),
.A2(n_33),
.B1(n_15),
.B2(n_38),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_70),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_131),
.B(n_143),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_49),
.A2(n_33),
.B1(n_85),
.B2(n_84),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_135),
.A2(n_18),
.B1(n_45),
.B2(n_4),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_93),
.A2(n_33),
.B1(n_42),
.B2(n_32),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_136),
.A2(n_35),
.B1(n_34),
.B2(n_29),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_51),
.A2(n_27),
.B1(n_42),
.B2(n_32),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_139),
.A2(n_15),
.B1(n_23),
.B2(n_38),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_77),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_55),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_62),
.B(n_27),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_150),
.B(n_5),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_99),
.Y(n_154)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

INVx3_ASAP7_75t_SL g155 ( 
.A(n_107),
.Y(n_155)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_155),
.Y(n_211)
);

AND2x2_ASAP7_75t_SL g156 ( 
.A(n_103),
.B(n_69),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_156),
.B(n_133),
.C(n_101),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_146),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_157),
.B(n_178),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_158),
.A2(n_163),
.B1(n_174),
.B2(n_188),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_159),
.B(n_168),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_35),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_160),
.B(n_164),
.Y(n_209)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_162),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_34),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_L g165 ( 
.A1(n_152),
.A2(n_65),
.B1(n_45),
.B2(n_29),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_165),
.A2(n_133),
.B1(n_125),
.B2(n_101),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_121),
.B(n_23),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_166),
.B(n_167),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_103),
.B(n_1),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_110),
.Y(n_168)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_169),
.Y(n_217)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_170),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_130),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_171),
.B(n_176),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_115),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_172),
.Y(n_218)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_109),
.Y(n_173)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_173),
.Y(n_220)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_175),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_127),
.B(n_2),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_2),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_177),
.B(n_8),
.Y(n_229)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_128),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_137),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_179),
.B(n_181),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_140),
.A2(n_18),
.B1(n_3),
.B2(n_4),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_180),
.A2(n_184),
.B1(n_189),
.B2(n_190),
.Y(n_227)
);

O2A1O1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_124),
.A2(n_2),
.B(n_5),
.C(n_7),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_111),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_182),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_151),
.B(n_112),
.Y(n_183)
);

AOI21xp33_ASAP7_75t_L g224 ( 
.A1(n_183),
.A2(n_191),
.B(n_104),
.Y(n_224)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_99),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_111),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_185),
.Y(n_216)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_132),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_187),
.Y(n_225)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_122),
.A2(n_2),
.B1(n_5),
.B2(n_7),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_132),
.Y(n_189)
);

INVx4_ASAP7_75t_SL g190 ( 
.A(n_104),
.Y(n_190)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_98),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_142),
.Y(n_228)
);

INVx4_ASAP7_75t_SL g193 ( 
.A(n_104),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_142),
.A2(n_8),
.B1(n_123),
.B2(n_145),
.Y(n_194)
);

OA22x2_ASAP7_75t_L g239 ( 
.A1(n_199),
.A2(n_184),
.B1(n_189),
.B2(n_186),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_195),
.A2(n_163),
.B1(n_152),
.B2(n_165),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_200),
.A2(n_219),
.B1(n_223),
.B2(n_193),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_202),
.B(n_206),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_160),
.A2(n_135),
.B1(n_120),
.B2(n_126),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_204),
.A2(n_187),
.B1(n_155),
.B2(n_168),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_156),
.B(n_98),
.C(n_126),
.Y(n_206)
);

AOI211xp5_ASAP7_75t_L g207 ( 
.A1(n_196),
.A2(n_156),
.B(n_159),
.C(n_167),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_207),
.A2(n_190),
.B(n_116),
.C(n_123),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_159),
.A2(n_125),
.B1(n_106),
.B2(n_144),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_164),
.B(n_119),
.C(n_142),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_229),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_172),
.A2(n_106),
.B1(n_102),
.B2(n_144),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_224),
.B(n_192),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_177),
.B(n_102),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_233),
.Y(n_246)
);

NOR2x1_ASAP7_75t_SL g231 ( 
.A(n_166),
.B(n_119),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_231),
.A2(n_169),
.B(n_185),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_119),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_197),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_234),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_232),
.A2(n_181),
.B(n_175),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_235),
.A2(n_250),
.B(n_252),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_236),
.B(n_241),
.Y(n_273)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_237),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_238),
.A2(n_258),
.B1(n_259),
.B2(n_227),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_239),
.B(n_223),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_173),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_209),
.B(n_161),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_243),
.B(n_257),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_244),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_247),
.A2(n_248),
.B1(n_254),
.B2(n_255),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_232),
.A2(n_102),
.B1(n_114),
.B2(n_116),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_249),
.B(n_253),
.Y(n_275)
);

AO21x2_ASAP7_75t_L g250 ( 
.A1(n_231),
.A2(n_154),
.B(n_116),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_205),
.Y(n_251)
);

INVx11_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_214),
.A2(n_114),
.B(n_123),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_209),
.B(n_114),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_204),
.A2(n_134),
.B1(n_144),
.B2(n_145),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_206),
.A2(n_134),
.B1(n_145),
.B2(n_199),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_226),
.Y(n_256)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_256),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_134),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_201),
.A2(n_207),
.B1(n_214),
.B2(n_233),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_201),
.A2(n_202),
.B1(n_221),
.B2(n_219),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_212),
.B(n_203),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_211),
.Y(n_285)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_256),
.Y(n_262)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_262),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_214),
.C(n_210),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_264),
.C(n_267),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_210),
.C(n_222),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_229),
.C(n_216),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_215),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_268),
.B(n_248),
.Y(n_307)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_237),
.Y(n_269)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_269),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_226),
.C(n_220),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_270),
.B(n_263),
.Y(n_308)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_241),
.Y(n_271)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_271),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_259),
.Y(n_287)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_239),
.Y(n_278)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_278),
.Y(n_306)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_279),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_260),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_282),
.Y(n_290)
);

INVx8_ASAP7_75t_L g282 ( 
.A(n_251),
.Y(n_282)
);

NOR3xp33_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_212),
.C(n_211),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_285),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_283),
.A2(n_249),
.B(n_245),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_286),
.B(n_292),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_287),
.A2(n_265),
.B1(n_270),
.B2(n_267),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_266),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_291),
.B(n_293),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_283),
.A2(n_236),
.B(n_250),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_261),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_243),
.Y(n_295)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_295),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_277),
.A2(n_250),
.B(n_244),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_299),
.Y(n_313)
);

XNOR2x2_ASAP7_75t_L g297 ( 
.A(n_268),
.B(n_250),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_297),
.B(n_275),
.Y(n_310)
);

O2A1O1Ixp33_ASAP7_75t_L g298 ( 
.A1(n_277),
.A2(n_250),
.B(n_239),
.C(n_247),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_298),
.B(n_307),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_268),
.A2(n_250),
.B(n_258),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_266),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_266),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_234),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g318 ( 
.A(n_302),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_278),
.A2(n_238),
.B1(n_253),
.B2(n_242),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_304),
.A2(n_276),
.B1(n_255),
.B2(n_254),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_242),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_310),
.B(n_299),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_311),
.B(n_314),
.Y(n_337)
);

OAI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_305),
.A2(n_274),
.B1(n_279),
.B2(n_273),
.Y(n_312)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_312),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_289),
.A2(n_265),
.B1(n_274),
.B2(n_279),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_305),
.Y(n_315)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_315),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_302),
.B(n_281),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_316),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_317),
.B(n_327),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_319),
.A2(n_324),
.B1(n_307),
.B2(n_297),
.Y(n_343)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_290),
.Y(n_320)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_320),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_295),
.B(n_290),
.Y(n_323)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_323),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_304),
.A2(n_275),
.B1(n_257),
.B2(n_239),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_328),
.C(n_288),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_294),
.B(n_264),
.Y(n_326)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_326),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_306),
.B(n_262),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_308),
.B(n_252),
.C(n_261),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_294),
.B(n_217),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_329),
.B(n_301),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_332),
.B(n_333),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_316),
.B(n_293),
.Y(n_334)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_334),
.Y(n_350)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_335),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_325),
.B(n_288),
.C(n_287),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_338),
.B(n_345),
.C(n_347),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_318),
.B(n_301),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_339),
.B(n_323),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_343),
.A2(n_298),
.B1(n_330),
.B2(n_327),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_328),
.B(n_292),
.C(n_286),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_314),
.A2(n_297),
.B1(n_289),
.B2(n_306),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_346),
.B(n_322),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_311),
.B(n_296),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_310),
.B(n_303),
.C(n_269),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_348),
.B(n_324),
.C(n_309),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_341),
.A2(n_320),
.B1(n_309),
.B2(n_315),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_352),
.A2(n_336),
.B1(n_337),
.B2(n_348),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_346),
.A2(n_313),
.B(n_321),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_353),
.A2(n_356),
.B(n_343),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_355),
.A2(n_344),
.B1(n_298),
.B2(n_332),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_347),
.A2(n_321),
.B(n_322),
.Y(n_356)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_357),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_359),
.B(n_360),
.C(n_354),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_338),
.B(n_319),
.C(n_330),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_340),
.Y(n_361)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_361),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_340),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_362),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_363),
.A2(n_331),
.B1(n_337),
.B2(n_342),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_364),
.B(n_366),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_365),
.B(n_369),
.Y(n_381)
);

INVxp33_ASAP7_75t_L g368 ( 
.A(n_353),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_368),
.B(n_370),
.Y(n_377)
);

FAx1_ASAP7_75t_SL g369 ( 
.A(n_355),
.B(n_333),
.CI(n_345),
.CON(n_369),
.SN(n_369)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_350),
.Y(n_371)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_371),
.Y(n_378)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_363),
.B(n_349),
.Y(n_372)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_372),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_375),
.B(n_359),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_379),
.B(n_377),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_373),
.A2(n_358),
.B1(n_360),
.B2(n_354),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_382),
.B(n_383),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_374),
.B(n_356),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_367),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_384),
.B(n_385),
.Y(n_390)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_372),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_381),
.A2(n_365),
.B(n_375),
.Y(n_386)
);

OAI21x1_ASAP7_75t_L g394 ( 
.A1(n_386),
.A2(n_393),
.B(n_379),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_387),
.B(n_389),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_376),
.Y(n_389)
);

AOI322xp5_ASAP7_75t_L g391 ( 
.A1(n_380),
.A2(n_368),
.A3(n_366),
.B1(n_291),
.B2(n_300),
.C1(n_303),
.C2(n_369),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_391),
.A2(n_282),
.B1(n_272),
.B2(n_251),
.Y(n_396)
);

CKINVDCx14_ASAP7_75t_R g392 ( 
.A(n_376),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_392),
.A2(n_351),
.B1(n_378),
.B2(n_282),
.Y(n_395)
);

OAI21x1_ASAP7_75t_L g393 ( 
.A1(n_384),
.A2(n_369),
.B(n_351),
.Y(n_393)
);

A2O1A1Ixp33_ASAP7_75t_L g403 ( 
.A1(n_394),
.A2(n_239),
.B(n_225),
.C(n_208),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_395),
.B(n_396),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_387),
.B(n_388),
.C(n_390),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_398),
.B(n_399),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_387),
.B(n_205),
.C(n_272),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_397),
.A2(n_225),
.B(n_220),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_402),
.B(n_398),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_403),
.B(n_399),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_404),
.B(n_405),
.Y(n_406)
);

NAND3xp33_ASAP7_75t_SL g407 ( 
.A(n_406),
.B(n_401),
.C(n_400),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_407),
.B(n_225),
.Y(n_408)
);


endmodule