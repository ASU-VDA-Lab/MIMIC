module fake_jpeg_22455_n_257 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_33),
.Y(n_54)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_25),
.B(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_39),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_41),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_28),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_41),
.A2(n_17),
.B1(n_27),
.B2(n_28),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_43),
.B1(n_45),
.B2(n_59),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_39),
.A2(n_17),
.B1(n_27),
.B2(n_28),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_17),
.B1(n_19),
.B2(n_21),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_40),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_46),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_28),
.C(n_23),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_38),
.Y(n_62)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_26),
.Y(n_52)
);

OA22x2_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_28),
.B1(n_23),
.B2(n_22),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_43),
.B(n_42),
.C(n_23),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_26),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_52),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_19),
.B1(n_21),
.B2(n_26),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_60),
.B(n_16),
.Y(n_110)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_35),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_64),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_38),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_65),
.B(n_73),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_22),
.B1(n_44),
.B2(n_32),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_21),
.B1(n_19),
.B2(n_18),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_70),
.A2(n_55),
.B(n_53),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_71),
.A2(n_81),
.B(n_45),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_30),
.Y(n_72)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_38),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_22),
.B1(n_31),
.B2(n_32),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_32),
.B1(n_31),
.B2(n_30),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_31),
.B1(n_29),
.B2(n_24),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_47),
.A2(n_36),
.B1(n_34),
.B2(n_29),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_85),
.B1(n_16),
.B2(n_33),
.Y(n_103)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_79),
.Y(n_88)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_59),
.A2(n_18),
.B(n_38),
.C(n_35),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_35),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_82),
.B(n_56),
.Y(n_90)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_55),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_24),
.Y(n_84)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_43),
.A2(n_36),
.B1(n_34),
.B2(n_20),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_87),
.A2(n_95),
.B(n_100),
.Y(n_130)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_108),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_99),
.C(n_105),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_62),
.A2(n_50),
.B1(n_54),
.B2(n_53),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_92),
.A2(n_102),
.B1(n_103),
.B2(n_109),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_0),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_108),
.Y(n_133)
);

NAND2x1_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_35),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_55),
.Y(n_98)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_65),
.B(n_33),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_67),
.A2(n_54),
.B1(n_53),
.B2(n_33),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_16),
.B(n_1),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_66),
.B(n_16),
.Y(n_107)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_0),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_71),
.A2(n_16),
.B1(n_1),
.B2(n_0),
.Y(n_109)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_97),
.B(n_72),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_112),
.B(n_124),
.Y(n_156)
);

NAND2x1p5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_81),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_113),
.A2(n_105),
.B(n_99),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_115),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_79),
.C(n_67),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_128),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_95),
.B(n_64),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_120),
.C(n_122),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_95),
.A2(n_71),
.B1(n_81),
.B2(n_63),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_63),
.Y(n_120)
);

MAJx2_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_84),
.C(n_83),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_97),
.B(n_60),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_68),
.C(n_80),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_99),
.C(n_105),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_68),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_127),
.Y(n_146)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_132),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_88),
.B(n_68),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_94),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_86),
.A2(n_80),
.B1(n_61),
.B2(n_1),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_135),
.A2(n_102),
.B1(n_93),
.B2(n_87),
.Y(n_142)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_106),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_141),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_115),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_140),
.Y(n_179)
);

OAI32xp33_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_109),
.A3(n_91),
.B1(n_92),
.B2(n_94),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_142),
.A2(n_143),
.B1(n_148),
.B2(n_151),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_113),
.A2(n_86),
.B1(n_103),
.B2(n_93),
.Y(n_143)
);

OAI221xp5_ASAP7_75t_L g177 ( 
.A1(n_147),
.A2(n_15),
.B1(n_3),
.B2(n_5),
.C(n_7),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_116),
.A2(n_119),
.B1(n_125),
.B2(n_130),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_163),
.C(n_131),
.Y(n_173)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_152),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_130),
.A2(n_91),
.B1(n_94),
.B2(n_99),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_107),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_154),
.Y(n_170)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_134),
.B(n_108),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_157),
.Y(n_183)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_108),
.Y(n_158)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_106),
.Y(n_160)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_116),
.A2(n_110),
.B(n_101),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g169 ( 
.A1(n_161),
.A2(n_114),
.B(n_123),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_101),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_162),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_61),
.C(n_1),
.Y(n_163)
);

OAI22x1_ASAP7_75t_SL g165 ( 
.A1(n_147),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_165),
.A2(n_172),
.B1(n_163),
.B2(n_138),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_173),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_150),
.A2(n_123),
.B1(n_121),
.B2(n_4),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_15),
.C(n_3),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_176),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_137),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_175),
.B(n_180),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_157),
.C(n_161),
.Y(n_176)
);

XNOR2x1_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_2),
.Y(n_203)
);

INVxp33_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_185),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_137),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_154),
.Y(n_182)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_156),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_184),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_2),
.C(n_7),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_170),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_186),
.B(n_187),
.Y(n_218)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_165),
.A2(n_139),
.B(n_162),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_189),
.A2(n_190),
.B(n_199),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_168),
.A2(n_159),
.B(n_145),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_164),
.A2(n_159),
.B1(n_143),
.B2(n_160),
.Y(n_191)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_155),
.Y(n_194)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_142),
.B1(n_151),
.B2(n_149),
.Y(n_195)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_146),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_198),
.B(n_171),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_179),
.B(n_156),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_178),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_201),
.A2(n_202),
.B(n_203),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_164),
.A2(n_141),
.B1(n_158),
.B2(n_140),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_181),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_205),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_176),
.C(n_173),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_207),
.C(n_211),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_166),
.C(n_181),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_208),
.B(n_213),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_214),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_166),
.C(n_171),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_183),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_211),
.B(n_198),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_219),
.B(n_223),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_209),
.A2(n_188),
.B1(n_194),
.B2(n_190),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_222),
.A2(n_228),
.B1(n_212),
.B2(n_174),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_207),
.B(n_189),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_191),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_224),
.B(n_226),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_196),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_9),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_214),
.B(n_197),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_217),
.A2(n_203),
.B1(n_200),
.B2(n_185),
.Y(n_228)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_230),
.Y(n_244)
);

OAI221xp5_ASAP7_75t_L g231 ( 
.A1(n_220),
.A2(n_183),
.B1(n_218),
.B2(n_215),
.C(n_216),
.Y(n_231)
);

NOR2xp67_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_221),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_227),
.A2(n_196),
.B1(n_7),
.B2(n_8),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_224),
.A2(n_2),
.B1(n_8),
.B2(n_9),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_233),
.B(n_227),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_8),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_237),
.C(n_238),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_9),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_225),
.C(n_221),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_235),
.C(n_236),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_242),
.A2(n_12),
.B(n_13),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_245),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_11),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_246),
.A2(n_247),
.B(n_250),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_238),
.C(n_13),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_12),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_14),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_248),
.A2(n_241),
.B1(n_239),
.B2(n_14),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_251),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_252),
.A2(n_14),
.B(n_253),
.Y(n_254)
);

BUFx24_ASAP7_75t_SL g256 ( 
.A(n_254),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_255),
.Y(n_257)
);


endmodule