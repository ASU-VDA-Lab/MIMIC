module real_jpeg_4252_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_400;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_0),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_0),
.B(n_182),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_0),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_0),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_0),
.B(n_287),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_0),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_0),
.B(n_376),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_0),
.B(n_105),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_1),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_1),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_1),
.Y(n_261)
);

INVx8_ASAP7_75t_L g312 ( 
.A(n_1),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_1),
.Y(n_332)
);

BUFx5_ASAP7_75t_L g349 ( 
.A(n_1),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_2),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_2),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_2),
.B(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_2),
.B(n_152),
.Y(n_151)
);

AND2x2_ASAP7_75t_SL g177 ( 
.A(n_2),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_2),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_2),
.B(n_215),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_3),
.Y(n_162)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_3),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_3),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_4),
.B(n_35),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_4),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_4),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_4),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_4),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_4),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_4),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_4),
.B(n_260),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_5),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_6),
.B(n_66),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_6),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_6),
.B(n_142),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_6),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_6),
.B(n_220),
.Y(n_219)
);

AND2x2_ASAP7_75t_SL g284 ( 
.A(n_6),
.B(n_200),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_6),
.B(n_373),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_6),
.B(n_193),
.Y(n_413)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_7),
.Y(n_86)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_7),
.Y(n_140)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_7),
.Y(n_232)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_8),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_9),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_9),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_9),
.B(n_307),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_9),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_9),
.B(n_353),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_9),
.B(n_96),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_9),
.B(n_292),
.Y(n_398)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_10),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_10),
.Y(n_180)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_10),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_10),
.Y(n_316)
);

BUFx5_ASAP7_75t_L g370 ( 
.A(n_10),
.Y(n_370)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_12),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_12),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_12),
.Y(n_272)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_14),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_14),
.B(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_14),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_14),
.B(n_292),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_14),
.B(n_332),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_14),
.B(n_347),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_14),
.B(n_409),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_15),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_15),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_15),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_15),
.B(n_310),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_15),
.B(n_329),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_15),
.B(n_180),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_15),
.B(n_385),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_15),
.B(n_356),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_16),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_16),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_16),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_16),
.B(n_340),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_16),
.B(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_16),
.B(n_388),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_16),
.B(n_400),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_17),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_17),
.B(n_59),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_17),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_17),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_17),
.B(n_96),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_17),
.B(n_270),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_17),
.B(n_289),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_17),
.B(n_310),
.Y(n_414)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_19),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_19),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_19),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_19),
.B(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_19),
.B(n_193),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_526),
.B(n_529),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_40),
.B(n_75),
.C(n_525),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_48),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_24),
.B(n_48),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_38),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.C(n_34),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_26),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_26),
.A2(n_30),
.B1(n_39),
.B2(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_28),
.Y(n_221)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_28),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_30),
.A2(n_52),
.B1(n_56),
.B2(n_57),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_30),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_30),
.B(n_52),
.C(n_58),
.Y(n_72)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_32),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_33),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_34),
.B(n_74),
.Y(n_73)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_37),
.Y(n_149)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_71),
.C(n_73),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_49),
.B(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_60),
.C(n_61),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_50),
.B(n_115),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_58),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_52),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_52),
.A2(n_57),
.B1(n_67),
.B2(n_108),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_54),
.Y(n_145)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_54),
.Y(n_275)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_55),
.Y(n_132)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_55),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_62),
.C(n_67),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_60),
.B(n_61),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_62),
.A2(n_63),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_65),
.Y(n_283)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_67),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_67),
.A2(n_103),
.B1(n_104),
.B2(n_108),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_69),
.Y(n_205)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_69),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_69),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_69),
.Y(n_409)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_71),
.A2(n_72),
.B1(n_73),
.B2(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

AO21x1_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_119),
.B(n_524),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_116),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_77),
.B(n_116),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_113),
.C(n_114),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_78),
.A2(n_79),
.B1(n_520),
.B2(n_521),
.Y(n_519)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_101),
.C(n_109),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_80),
.A2(n_81),
.B1(n_501),
.B2(n_503),
.Y(n_500)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_90),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_87),
.C(n_90),
.Y(n_113)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_89),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_89),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_89),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_89),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.C(n_97),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_91),
.B(n_491),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_92),
.A2(n_93),
.B1(n_97),
.B2(n_98),
.Y(n_491)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx6_ASAP7_75t_SL g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_101),
.A2(n_109),
.B1(n_110),
.B2(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_101),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.C(n_108),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g496 ( 
.A(n_102),
.B(n_497),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_103),
.A2(n_104),
.B1(n_192),
.B2(n_195),
.Y(n_191)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_104),
.B(n_188),
.C(n_192),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_107),
.Y(n_290)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_113),
.B(n_114),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_518),
.B(n_523),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_484),
.B(n_515),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_295),
.B(n_483),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_245),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_123),
.B(n_245),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_185),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_124),
.B(n_186),
.C(n_222),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_159),
.C(n_168),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_125),
.B(n_248),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_136),
.C(n_146),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_126),
.B(n_468),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_130),
.C(n_133),
.Y(n_167)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_128),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_136),
.A2(n_137),
.B1(n_146),
.B2(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.C(n_144),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_138),
.B(n_144),
.Y(n_458)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_141),
.B(n_458),
.Y(n_457)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_146),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_147),
.B(n_151),
.C(n_156),
.Y(n_242)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_155),
.B1(n_156),
.B2(n_158),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_151),
.Y(n_158)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_154),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_154),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_155),
.B(n_192),
.C(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_155),
.A2(n_156),
.B1(n_192),
.B2(n_195),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_159),
.B(n_168),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_167),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_163),
.B1(n_165),
.B2(n_166),
.Y(n_160)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_161),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_163),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_163),
.B(n_165),
.C(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_163),
.A2(n_166),
.B1(n_234),
.B2(n_238),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_166),
.B(n_227),
.C(n_238),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_167),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_179),
.C(n_181),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_169),
.B(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.C(n_177),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_170),
.B(n_257),
.Y(n_256)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_174),
.B(n_177),
.Y(n_257)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_179),
.B(n_181),
.Y(n_278)
);

INVx4_ASAP7_75t_SL g182 ( 
.A(n_183),
.Y(n_182)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_222),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_196),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_187),
.B(n_197),
.C(n_206),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_192),
.Y(n_195)
);

BUFx8_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_206),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.C(n_203),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_198),
.B(n_203),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_199),
.B(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_201),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx8_ASAP7_75t_L g353 ( 
.A(n_205),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_219),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_214),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_208),
.B(n_214),
.C(n_219),
.Y(n_499)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_213),
.Y(n_357)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_218),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_239),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_224),
.B(n_226),
.C(n_239),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_233),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_228),
.B(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx6_ASAP7_75t_L g267 ( 
.A(n_232),
.Y(n_267)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_234),
.Y(n_238)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx8_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.C(n_243),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_243),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_249),
.C(n_252),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_247),
.B(n_250),
.Y(n_478)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_252),
.B(n_478),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_276),
.C(n_279),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_254),
.B(n_471),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.C(n_264),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_255),
.A2(n_256),
.B1(n_449),
.B2(n_450),
.Y(n_448)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_258),
.A2(n_259),
.B(n_262),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_258),
.B(n_264),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

MAJx2_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_268),
.C(n_273),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_265),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_426)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_272),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_272),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_273),
.B(n_426),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_274),
.B(n_369),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_276),
.A2(n_277),
.B1(n_279),
.B2(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_279),
.Y(n_472)
);

MAJx2_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_288),
.C(n_291),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_281),
.B(n_460),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.C(n_285),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_282),
.B(n_438),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g439 ( 
.A(n_284),
.Y(n_439)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_288),
.B(n_291),
.Y(n_460)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx6_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

AOI21x1_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_476),
.B(n_482),
.Y(n_295)
);

OAI21x1_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_463),
.B(n_475),
.Y(n_296)
);

AOI21x1_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_445),
.B(n_462),
.Y(n_297)
);

OAI21x1_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_419),
.B(n_444),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_300),
.A2(n_393),
.B(n_418),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_361),
.B(n_392),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_342),
.B(n_360),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_323),
.B(n_341),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_317),
.B(n_322),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_313),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_313),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_309),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_318),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_309),
.Y(n_324)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx8_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_312),
.Y(n_321)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_312),
.Y(n_373)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_324),
.B(n_325),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_326),
.A2(n_327),
.B1(n_333),
.B2(n_334),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_326),
.B(n_336),
.C(n_338),
.Y(n_359)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_331),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_328),
.B(n_331),
.Y(n_350)
);

INVx8_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_335),
.A2(n_336),
.B1(n_338),
.B2(n_339),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_343),
.B(n_359),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_343),
.B(n_359),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_351),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_350),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_345),
.B(n_350),
.C(n_363),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_348),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_346),
.B(n_348),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_351),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_354),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_352),
.B(n_381),
.C(n_382),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_358),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_355),
.Y(n_381)
);

INVx6_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_358),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_364),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_362),
.B(n_364),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_379),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_365),
.B(n_380),
.C(n_383),
.Y(n_417)
);

XOR2x2_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_366),
.B(n_368),
.C(n_371),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_371),
.Y(n_367)
);

INVx4_ASAP7_75t_SL g369 ( 
.A(n_370),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_372),
.A2(n_374),
.B1(n_375),
.B2(n_378),
.Y(n_371)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_372),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_374),
.B(n_378),
.Y(n_402)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_383),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_386),
.Y(n_383)
);

MAJx2_ASAP7_75t_L g416 ( 
.A(n_384),
.B(n_389),
.C(n_390),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_387),
.A2(n_389),
.B1(n_390),
.B2(n_391),
.Y(n_386)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_387),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_389),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_394),
.B(n_417),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_394),
.B(n_417),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_395),
.B(n_404),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_403),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_396),
.B(n_403),
.C(n_443),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_402),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_399),
.Y(n_397)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_398),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_399),
.Y(n_434)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_402),
.B(n_433),
.C(n_434),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_404),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_410),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_405),
.B(n_412),
.C(n_415),
.Y(n_422)
);

BUFx24_ASAP7_75t_SL g532 ( 
.A(n_405),
.Y(n_532)
);

FAx1_ASAP7_75t_SL g405 ( 
.A(n_406),
.B(n_407),
.CI(n_408),
.CON(n_405),
.SN(n_405)
);

MAJx2_ASAP7_75t_L g430 ( 
.A(n_406),
.B(n_407),
.C(n_408),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_411),
.A2(n_412),
.B1(n_415),
.B2(n_416),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_414),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_413),
.B(n_414),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_416),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_420),
.B(n_442),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_420),
.B(n_442),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_431),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_422),
.B(n_423),
.C(n_431),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_424),
.A2(n_425),
.B1(n_427),
.B2(n_428),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_424),
.B(n_454),
.C(n_455),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.Y(n_428)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_429),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_430),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g431 ( 
.A(n_432),
.B(n_435),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_432),
.B(n_436),
.C(n_441),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_436),
.A2(n_437),
.B1(n_440),
.B2(n_441),
.Y(n_435)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_436),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_437),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_446),
.B(n_461),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_446),
.B(n_461),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_447),
.B(n_452),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_451),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_448),
.B(n_451),
.C(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_449),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_452),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_453),
.B(n_456),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_453),
.B(n_457),
.C(n_459),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_459),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_464),
.B(n_473),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_473),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_466),
.Y(n_464)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_465),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_470),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_467),
.B(n_480),
.C(n_481),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_470),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_477),
.B(n_479),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_477),
.B(n_479),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_512),
.Y(n_484)
);

OAI21xp33_ASAP7_75t_L g515 ( 
.A1(n_485),
.A2(n_516),
.B(n_517),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_486),
.B(n_505),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_486),
.B(n_505),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_487),
.A2(n_488),
.B1(n_494),
.B2(n_504),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_487),
.B(n_495),
.C(n_500),
.Y(n_522)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_490),
.C(n_492),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_489),
.B(n_507),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_490),
.A2(n_492),
.B1(n_493),
.B2(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_490),
.Y(n_508)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_494),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_500),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_498),
.C(n_499),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_496),
.B(n_510),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_498),
.B(n_499),
.Y(n_510)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_501),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_509),
.C(n_511),
.Y(n_505)
);

FAx1_ASAP7_75t_SL g513 ( 
.A(n_506),
.B(n_509),
.CI(n_511),
.CON(n_513),
.SN(n_513)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_513),
.B(n_514),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_513),
.B(n_514),
.Y(n_516)
);

BUFx24_ASAP7_75t_SL g533 ( 
.A(n_513),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_522),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_519),
.B(n_522),
.Y(n_523)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_520),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx5_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx6_ASAP7_75t_L g530 ( 
.A(n_528),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_530),
.B(n_531),
.Y(n_529)
);


endmodule