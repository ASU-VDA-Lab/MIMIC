module fake_aes_12341_n_686 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_93, n_51, n_39, n_686);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_93;
input n_51;
input n_39;
output n_686;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_482;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx6f_ASAP7_75t_L g95 ( .A(n_86), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_28), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_44), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_42), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_38), .Y(n_99) );
OR2x2_ASAP7_75t_L g100 ( .A(n_3), .B(n_50), .Y(n_100) );
BUFx3_ASAP7_75t_L g101 ( .A(n_79), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_85), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_11), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_83), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_23), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_14), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_72), .Y(n_107) );
BUFx3_ASAP7_75t_L g108 ( .A(n_67), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_62), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_61), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_31), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_24), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_6), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_55), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_88), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_89), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_93), .Y(n_117) );
BUFx3_ASAP7_75t_L g118 ( .A(n_43), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_69), .Y(n_119) );
INVxp33_ASAP7_75t_L g120 ( .A(n_40), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_18), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_91), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_22), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_7), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_35), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_21), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_77), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_46), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_15), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_57), .Y(n_130) );
CKINVDCx14_ASAP7_75t_R g131 ( .A(n_56), .Y(n_131) );
NOR2xp67_ASAP7_75t_L g132 ( .A(n_15), .B(n_59), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_73), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_68), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_25), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_2), .Y(n_136) );
BUFx2_ASAP7_75t_L g137 ( .A(n_36), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_0), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_117), .B(n_0), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_117), .B(n_1), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_137), .B(n_1), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_105), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_137), .B(n_2), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_95), .Y(n_144) );
BUFx8_ASAP7_75t_L g145 ( .A(n_95), .Y(n_145) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_113), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_104), .B(n_3), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_125), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_125), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_120), .B(n_4), .Y(n_150) );
CKINVDCx11_ASAP7_75t_R g151 ( .A(n_124), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_131), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_105), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_106), .B(n_4), .Y(n_154) );
AND2x4_ASAP7_75t_L g155 ( .A(n_106), .B(n_5), .Y(n_155) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_107), .A2(n_45), .B(n_92), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_107), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_144), .Y(n_158) );
NAND2xp33_ASAP7_75t_R g159 ( .A(n_152), .B(n_113), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_155), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_146), .B(n_96), .Y(n_161) );
AO22x2_ASAP7_75t_L g162 ( .A1(n_155), .A2(n_100), .B1(n_130), .B2(n_109), .Y(n_162) );
OR2x6_ASAP7_75t_L g163 ( .A(n_139), .B(n_100), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_144), .Y(n_164) );
OAI22xp33_ASAP7_75t_L g165 ( .A1(n_141), .A2(n_138), .B1(n_103), .B2(n_129), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_156), .Y(n_166) );
AOI22xp5_ASAP7_75t_L g167 ( .A1(n_139), .A2(n_138), .B1(n_136), .B2(n_103), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_155), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_155), .Y(n_169) );
OR2x2_ASAP7_75t_L g170 ( .A(n_143), .B(n_129), .Y(n_170) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_150), .A2(n_126), .B1(n_121), .B2(n_102), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_144), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_154), .Y(n_173) );
INVx2_ASAP7_75t_SL g174 ( .A(n_145), .Y(n_174) );
INVx3_ASAP7_75t_L g175 ( .A(n_148), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_148), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_150), .B(n_121), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_149), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_152), .B(n_98), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_142), .B(n_98), .Y(n_180) );
INVx2_ASAP7_75t_SL g181 ( .A(n_145), .Y(n_181) );
INVx3_ASAP7_75t_L g182 ( .A(n_149), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_163), .B(n_173), .Y(n_183) );
AND2x6_ASAP7_75t_SL g184 ( .A(n_163), .B(n_151), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_158), .Y(n_185) );
BUFx12f_ASAP7_75t_L g186 ( .A(n_163), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_177), .B(n_142), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_159), .Y(n_188) );
INVxp67_ASAP7_75t_L g189 ( .A(n_163), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_174), .B(n_147), .Y(n_190) );
OR2x2_ASAP7_75t_L g191 ( .A(n_171), .B(n_140), .Y(n_191) );
AND2x4_ASAP7_75t_L g192 ( .A(n_177), .B(n_170), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_160), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_158), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_170), .B(n_154), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_174), .B(n_99), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_160), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_180), .B(n_153), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_162), .A2(n_157), .B1(n_153), .B2(n_145), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_162), .B(n_157), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_179), .B(n_99), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_181), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_161), .B(n_102), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_168), .B(n_145), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_164), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_176), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_169), .B(n_109), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_181), .B(n_97), .Y(n_208) );
AOI21x1_ASAP7_75t_L g209 ( .A1(n_164), .A2(n_156), .B(n_110), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_162), .B(n_110), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_172), .Y(n_211) );
INVx5_ASAP7_75t_L g212 ( .A(n_175), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_176), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_178), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_178), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_185), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_192), .B(n_162), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_192), .B(n_167), .Y(n_218) );
BUFx3_ASAP7_75t_L g219 ( .A(n_202), .Y(n_219) );
CKINVDCx10_ASAP7_75t_R g220 ( .A(n_184), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_204), .A2(n_166), .B(n_156), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g222 ( .A1(n_195), .A2(n_165), .B1(n_175), .B2(n_182), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_192), .B(n_182), .Y(n_223) );
OAI22x1_ASAP7_75t_L g224 ( .A1(n_183), .A2(n_156), .B1(n_128), .B2(n_130), .Y(n_224) );
OA22x2_ASAP7_75t_L g225 ( .A1(n_183), .A2(n_182), .B1(n_175), .B2(n_128), .Y(n_225) );
CKINVDCx14_ASAP7_75t_R g226 ( .A(n_186), .Y(n_226) );
INVx3_ASAP7_75t_L g227 ( .A(n_212), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_202), .B(n_166), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_192), .B(n_166), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_L g230 ( .A1(n_210), .A2(n_116), .B(n_135), .C(n_134), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g231 ( .A1(n_186), .A2(n_166), .B1(n_123), .B2(n_115), .Y(n_231) );
INVx1_ASAP7_75t_SL g232 ( .A(n_186), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_187), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_190), .A2(n_193), .B(n_197), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_183), .B(n_166), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_184), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_193), .A2(n_172), .B(n_111), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_189), .B(n_112), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_197), .A2(n_127), .B(n_118), .Y(n_239) );
NAND3xp33_ASAP7_75t_L g240 ( .A(n_199), .B(n_132), .C(n_118), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_202), .B(n_95), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_183), .B(n_101), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_206), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_185), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_200), .B(n_101), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g246 ( .A1(n_222), .A2(n_191), .B(n_203), .C(n_207), .Y(n_246) );
BUFx4f_ASAP7_75t_SL g247 ( .A(n_232), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_228), .A2(n_208), .B(n_196), .Y(n_248) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_226), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_233), .B(n_191), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_243), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_218), .B(n_200), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_217), .A2(n_215), .B1(n_214), .B2(n_213), .Y(n_253) );
OAI21xp5_ASAP7_75t_L g254 ( .A1(n_234), .A2(n_215), .B(n_214), .Y(n_254) );
AO31x2_ASAP7_75t_L g255 ( .A1(n_224), .A2(n_213), .A3(n_206), .B(n_194), .Y(n_255) );
AO21x2_ASAP7_75t_L g256 ( .A1(n_221), .A2(n_209), .B(n_198), .Y(n_256) );
BUFx2_ASAP7_75t_L g257 ( .A(n_226), .Y(n_257) );
INVx1_ASAP7_75t_SL g258 ( .A(n_216), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_SL g259 ( .A1(n_241), .A2(n_211), .B(n_205), .C(n_185), .Y(n_259) );
AO31x2_ASAP7_75t_L g260 ( .A1(n_229), .A2(n_211), .A3(n_205), .B(n_194), .Y(n_260) );
BUFx10_ASAP7_75t_L g261 ( .A(n_245), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_228), .A2(n_211), .B(n_205), .Y(n_262) );
BUFx3_ASAP7_75t_L g263 ( .A(n_216), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_223), .B(n_201), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_238), .B(n_188), .Y(n_265) );
BUFx4f_ASAP7_75t_SL g266 ( .A(n_220), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_244), .B(n_212), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_244), .Y(n_268) );
OAI21x1_ASAP7_75t_L g269 ( .A1(n_241), .A2(n_209), .B(n_194), .Y(n_269) );
OA21x2_ASAP7_75t_L g270 ( .A1(n_269), .A2(n_240), .B(n_239), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_268), .Y(n_271) );
INVx3_ASAP7_75t_L g272 ( .A(n_263), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_263), .Y(n_273) );
INVx2_ASAP7_75t_SL g274 ( .A(n_261), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_268), .Y(n_275) );
AND2x4_ASAP7_75t_L g276 ( .A(n_251), .B(n_227), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_251), .Y(n_277) );
AO21x2_ASAP7_75t_L g278 ( .A1(n_254), .A2(n_235), .B(n_242), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_258), .Y(n_279) );
INVxp67_ASAP7_75t_L g280 ( .A(n_267), .Y(n_280) );
OAI21x1_ASAP7_75t_L g281 ( .A1(n_269), .A2(n_225), .B(n_237), .Y(n_281) );
A2O1A1Ixp33_ASAP7_75t_L g282 ( .A1(n_246), .A2(n_230), .B(n_245), .C(n_219), .Y(n_282) );
AND2x4_ASAP7_75t_L g283 ( .A(n_258), .B(n_267), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_260), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_250), .A2(n_225), .B1(n_245), .B2(n_236), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_256), .Y(n_286) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_260), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_260), .Y(n_288) );
AO31x2_ASAP7_75t_L g289 ( .A1(n_252), .A2(n_231), .A3(n_119), .B(n_122), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_260), .Y(n_290) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_287), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_277), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_271), .B(n_253), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_271), .B(n_253), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_277), .B(n_260), .Y(n_295) );
AND3x1_ASAP7_75t_L g296 ( .A(n_285), .B(n_266), .C(n_236), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_286), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_275), .Y(n_298) );
BUFx3_ASAP7_75t_L g299 ( .A(n_273), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_275), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_284), .Y(n_301) );
AO21x1_ASAP7_75t_SL g302 ( .A1(n_288), .A2(n_261), .B(n_259), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_284), .B(n_255), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_284), .B(n_261), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_284), .Y(n_305) );
AO21x2_ASAP7_75t_L g306 ( .A1(n_286), .A2(n_256), .B(n_262), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_286), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_288), .Y(n_308) );
BUFx2_ASAP7_75t_L g309 ( .A(n_273), .Y(n_309) );
AO31x2_ASAP7_75t_L g310 ( .A1(n_290), .A2(n_264), .A3(n_248), .B(n_255), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_290), .B(n_257), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_285), .A2(n_265), .B1(n_257), .B2(n_261), .Y(n_312) );
INVx2_ASAP7_75t_SL g313 ( .A(n_273), .Y(n_313) );
AO21x1_ASAP7_75t_SL g314 ( .A1(n_287), .A2(n_273), .B(n_272), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_279), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_280), .B(n_255), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_297), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_301), .B(n_283), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_297), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_301), .B(n_283), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_293), .B(n_276), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_308), .Y(n_322) );
BUFx3_ASAP7_75t_L g323 ( .A(n_309), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_305), .B(n_283), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_308), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_305), .B(n_283), .Y(n_326) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_311), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_304), .B(n_283), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_295), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_291), .B(n_279), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_304), .B(n_279), .Y(n_331) );
AND2x4_ASAP7_75t_SL g332 ( .A(n_313), .B(n_272), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_297), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_299), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_291), .B(n_289), .Y(n_335) );
INVx2_ASAP7_75t_SL g336 ( .A(n_299), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_295), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_292), .B(n_272), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_307), .Y(n_339) );
INVx5_ASAP7_75t_SL g340 ( .A(n_314), .Y(n_340) );
OR2x6_ASAP7_75t_L g341 ( .A(n_309), .B(n_272), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_311), .B(n_289), .Y(n_342) );
BUFx2_ASAP7_75t_L g343 ( .A(n_299), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_292), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_293), .B(n_276), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_316), .B(n_289), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_298), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_298), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_303), .B(n_272), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_294), .B(n_276), .Y(n_350) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_313), .Y(n_351) );
NAND2x1p5_ASAP7_75t_SL g352 ( .A(n_313), .B(n_274), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_300), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_307), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_307), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_316), .B(n_289), .Y(n_356) );
BUFx2_ASAP7_75t_L g357 ( .A(n_315), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_315), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_300), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_322), .Y(n_360) );
OAI21xp5_ASAP7_75t_SL g361 ( .A1(n_340), .A2(n_312), .B(n_294), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_349), .B(n_303), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_342), .B(n_303), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_322), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_325), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_317), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_325), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_349), .B(n_314), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_344), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_318), .B(n_315), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_344), .Y(n_371) );
NOR2xp67_ASAP7_75t_L g372 ( .A(n_335), .B(n_274), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_347), .Y(n_373) );
INVx3_ASAP7_75t_L g374 ( .A(n_340), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_318), .B(n_310), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_317), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_347), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_320), .B(n_324), .Y(n_378) );
BUFx2_ASAP7_75t_L g379 ( .A(n_352), .Y(n_379) );
INVx1_ASAP7_75t_SL g380 ( .A(n_334), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_320), .B(n_310), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_317), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_351), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_319), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_324), .B(n_310), .Y(n_385) );
NOR2xp67_ASAP7_75t_SL g386 ( .A(n_340), .B(n_274), .Y(n_386) );
INVxp67_ASAP7_75t_SL g387 ( .A(n_357), .Y(n_387) );
NAND2x1_ASAP7_75t_SL g388 ( .A(n_340), .B(n_270), .Y(n_388) );
OR2x2_ASAP7_75t_L g389 ( .A(n_342), .B(n_310), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_326), .B(n_310), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_327), .B(n_310), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_335), .B(n_310), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_326), .B(n_306), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_321), .B(n_247), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_348), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_329), .B(n_306), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_348), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_329), .B(n_306), .Y(n_398) );
INVx3_ASAP7_75t_L g399 ( .A(n_340), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_337), .B(n_306), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_337), .B(n_302), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_331), .B(n_302), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_331), .B(n_289), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_319), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_339), .B(n_289), .Y(n_405) );
NOR2x1_ASAP7_75t_L g406 ( .A(n_341), .B(n_282), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_353), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_353), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_359), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_359), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_339), .B(n_289), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_330), .Y(n_412) );
INVx3_ASAP7_75t_L g413 ( .A(n_339), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_333), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_339), .B(n_289), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_328), .B(n_278), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_328), .B(n_278), .Y(n_417) );
AND2x4_ASAP7_75t_L g418 ( .A(n_338), .B(n_323), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_330), .Y(n_419) );
AND2x4_ASAP7_75t_L g420 ( .A(n_338), .B(n_278), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_333), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_354), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_346), .B(n_278), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_346), .B(n_278), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_368), .B(n_343), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_396), .B(n_356), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_363), .B(n_356), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_360), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_366), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_368), .B(n_343), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_372), .B(n_323), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_378), .B(n_323), .Y(n_432) );
INVxp67_ASAP7_75t_L g433 ( .A(n_379), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_360), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_364), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_364), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_378), .B(n_336), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_366), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_365), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_383), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_366), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_363), .B(n_345), .Y(n_442) );
NAND2x1_ASAP7_75t_L g443 ( .A(n_374), .B(n_341), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_365), .Y(n_444) );
NAND2x1p5_ASAP7_75t_L g445 ( .A(n_386), .B(n_374), .Y(n_445) );
AND2x4_ASAP7_75t_L g446 ( .A(n_372), .B(n_336), .Y(n_446) );
INVx1_ASAP7_75t_SL g447 ( .A(n_379), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_362), .B(n_341), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_362), .B(n_341), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_396), .B(n_400), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_376), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_412), .B(n_350), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_367), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_400), .B(n_354), .Y(n_454) );
NOR2x1p5_ASAP7_75t_SL g455 ( .A(n_398), .B(n_355), .Y(n_455) );
INVxp33_ASAP7_75t_L g456 ( .A(n_386), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_376), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_419), .B(n_357), .Y(n_458) );
NAND2x1_ASAP7_75t_SL g459 ( .A(n_374), .B(n_355), .Y(n_459) );
NAND2xp33_ASAP7_75t_R g460 ( .A(n_374), .B(n_341), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_402), .B(n_418), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_402), .B(n_332), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_367), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_369), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_376), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_369), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_371), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_418), .B(n_332), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_418), .B(n_332), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_389), .B(n_352), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_423), .B(n_358), .Y(n_471) );
NOR2x1_ASAP7_75t_L g472 ( .A(n_399), .B(n_358), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_399), .B(n_296), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_371), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_423), .B(n_352), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_382), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_389), .B(n_5), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_418), .B(n_296), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_375), .B(n_95), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_373), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_392), .B(n_6), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_375), .B(n_381), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_373), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_377), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_392), .B(n_7), .Y(n_485) );
INVxp67_ASAP7_75t_L g486 ( .A(n_387), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_381), .B(n_95), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_385), .B(n_8), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_424), .B(n_282), .Y(n_489) );
INVx2_ASAP7_75t_SL g490 ( .A(n_380), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_377), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_385), .B(n_119), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_390), .B(n_119), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_382), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_424), .B(n_270), .Y(n_495) );
OR2x6_ASAP7_75t_L g496 ( .A(n_399), .B(n_276), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_361), .B(n_8), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_395), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_394), .A2(n_276), .B1(n_280), .B2(n_270), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_391), .B(n_270), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_395), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_401), .B(n_119), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_390), .B(n_270), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_382), .Y(n_504) );
INVx4_ASAP7_75t_L g505 ( .A(n_399), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_384), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_497), .A2(n_401), .B1(n_393), .B2(n_420), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_450), .B(n_427), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_504), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_479), .B(n_393), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_440), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_461), .B(n_416), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_486), .Y(n_513) );
INVx2_ASAP7_75t_SL g514 ( .A(n_490), .Y(n_514) );
NAND2xp33_ASAP7_75t_L g515 ( .A(n_456), .B(n_406), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_482), .B(n_416), .Y(n_516) );
AND2x4_ASAP7_75t_L g517 ( .A(n_455), .B(n_405), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_428), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_497), .B(n_397), .Y(n_519) );
NAND3xp33_ASAP7_75t_L g520 ( .A(n_487), .B(n_406), .C(n_119), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_504), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_450), .B(n_403), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_492), .B(n_493), .Y(n_523) );
OAI211xp5_ASAP7_75t_SL g524 ( .A1(n_473), .A2(n_249), .B(n_398), .C(n_397), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_488), .B(n_407), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_434), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_426), .B(n_417), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_458), .Y(n_528) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_502), .Y(n_529) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_473), .A2(n_388), .B(n_403), .C(n_405), .Y(n_530) );
BUFx3_ASAP7_75t_L g531 ( .A(n_437), .Y(n_531) );
OAI22xp33_ASAP7_75t_SL g532 ( .A1(n_477), .A2(n_409), .B1(n_407), .B2(n_408), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_481), .A2(n_411), .B1(n_415), .B2(n_417), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_432), .B(n_370), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_478), .B(n_408), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_435), .Y(n_536) );
INVx1_ASAP7_75t_SL g537 ( .A(n_447), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_476), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_426), .B(n_370), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_471), .B(n_442), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_436), .Y(n_541) );
AOI221xp5_ASAP7_75t_SL g542 ( .A1(n_433), .A2(n_410), .B1(n_409), .B2(n_415), .C(n_411), .Y(n_542) );
INVx1_ASAP7_75t_SL g543 ( .A(n_447), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_471), .B(n_410), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_425), .B(n_420), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_439), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_452), .B(n_420), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_476), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_444), .Y(n_549) );
INVx2_ASAP7_75t_SL g550 ( .A(n_430), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_489), .A2(n_420), .B1(n_413), .B2(n_133), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_453), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_463), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_475), .B(n_414), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_464), .Y(n_555) );
AND2x2_ASAP7_75t_SL g556 ( .A(n_505), .B(n_413), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_466), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_502), .B(n_414), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_467), .B(n_422), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_474), .B(n_422), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_485), .B(n_384), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_480), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_448), .B(n_413), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_449), .B(n_413), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_483), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_484), .B(n_384), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_491), .B(n_404), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_498), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_468), .B(n_421), .Y(n_569) );
INVxp67_ASAP7_75t_SL g570 ( .A(n_486), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_501), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_469), .B(n_421), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_454), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_462), .B(n_421), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_454), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_475), .B(n_404), .Y(n_576) );
INVx2_ASAP7_75t_SL g577 ( .A(n_446), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_470), .B(n_404), .Y(n_578) );
CKINVDCx20_ASAP7_75t_R g579 ( .A(n_505), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_506), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_579), .A2(n_456), .B1(n_445), .B2(n_443), .Y(n_581) );
OA22x2_ASAP7_75t_L g582 ( .A1(n_507), .A2(n_433), .B1(n_496), .B2(n_431), .Y(n_582) );
AOI32xp33_ASAP7_75t_L g583 ( .A1(n_524), .A2(n_446), .A3(n_431), .B1(n_472), .B2(n_499), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_509), .Y(n_584) );
OAI31xp33_ASAP7_75t_SL g585 ( .A1(n_570), .A2(n_460), .A3(n_445), .B(n_459), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_519), .A2(n_460), .B1(n_496), .B2(n_489), .Y(n_586) );
OAI31xp33_ASAP7_75t_L g587 ( .A1(n_532), .A2(n_503), .A3(n_499), .B(n_495), .Y(n_587) );
NOR4xp25_ASAP7_75t_SL g588 ( .A(n_511), .B(n_496), .C(n_388), .D(n_500), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_530), .A2(n_495), .B1(n_500), .B2(n_494), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_513), .Y(n_590) );
NAND2xp33_ASAP7_75t_SL g591 ( .A(n_577), .B(n_429), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_544), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_573), .B(n_465), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_544), .Y(n_594) );
AOI221xp5_ASAP7_75t_L g595 ( .A1(n_532), .A2(n_133), .B1(n_122), .B2(n_441), .C(n_438), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_554), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_575), .B(n_451), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_512), .B(n_457), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_518), .Y(n_599) );
AOI222xp33_ASAP7_75t_L g600 ( .A1(n_533), .A2(n_133), .B1(n_122), .B2(n_114), .C1(n_108), .C2(n_281), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_533), .A2(n_270), .B1(n_122), .B2(n_133), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_531), .A2(n_122), .B1(n_133), .B2(n_108), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_542), .B(n_255), .Y(n_603) );
AND2x4_ASAP7_75t_L g604 ( .A(n_517), .B(n_281), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_514), .B(n_9), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_516), .B(n_281), .Y(n_606) );
AOI32xp33_ASAP7_75t_L g607 ( .A1(n_515), .A2(n_114), .A3(n_227), .B1(n_11), .B2(n_12), .Y(n_607) );
AOI322xp5_ASAP7_75t_L g608 ( .A1(n_542), .A2(n_527), .A3(n_525), .B1(n_535), .B2(n_550), .C1(n_534), .C2(n_545), .Y(n_608) );
AO22x1_ASAP7_75t_L g609 ( .A1(n_517), .A2(n_9), .B1(n_10), .B2(n_12), .Y(n_609) );
AO22x1_ASAP7_75t_L g610 ( .A1(n_529), .A2(n_10), .B1(n_13), .B2(n_14), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_563), .B(n_255), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_564), .B(n_256), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_526), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_536), .Y(n_614) );
INVxp67_ASAP7_75t_L g615 ( .A(n_537), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_569), .B(n_16), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g617 ( .A1(n_520), .A2(n_16), .B(n_17), .Y(n_617) );
AOI32xp33_ASAP7_75t_L g618 ( .A1(n_537), .A2(n_17), .A3(n_18), .B1(n_219), .B2(n_20), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_572), .B(n_19), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_576), .B(n_26), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_541), .Y(n_621) );
INVx1_ASAP7_75t_SL g622 ( .A(n_543), .Y(n_622) );
AOI22x1_ASAP7_75t_L g623 ( .A1(n_543), .A2(n_27), .B1(n_29), .B2(n_30), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_523), .A2(n_556), .B1(n_529), .B2(n_510), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_546), .Y(n_625) );
OAI221xp5_ASAP7_75t_SL g626 ( .A1(n_608), .A2(n_551), .B1(n_508), .B2(n_547), .C(n_540), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_590), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_596), .Y(n_628) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_587), .A2(n_528), .B1(n_552), .B2(n_553), .C(n_571), .Y(n_629) );
AO21x1_ASAP7_75t_L g630 ( .A1(n_591), .A2(n_558), .B(n_549), .Y(n_630) );
OAI221xp5_ASAP7_75t_L g631 ( .A1(n_583), .A2(n_561), .B1(n_555), .B2(n_562), .C(n_568), .Y(n_631) );
O2A1O1Ixp5_ASAP7_75t_SL g632 ( .A1(n_602), .A2(n_557), .B(n_565), .C(n_580), .Y(n_632) );
OAI22xp33_ASAP7_75t_SL g633 ( .A1(n_589), .A2(n_522), .B1(n_539), .B2(n_559), .Y(n_633) );
O2A1O1Ixp33_ASAP7_75t_L g634 ( .A1(n_617), .A2(n_521), .B(n_560), .C(n_559), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_592), .B(n_578), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_594), .Y(n_636) );
AO21x1_ASAP7_75t_L g637 ( .A1(n_581), .A2(n_560), .B(n_567), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_582), .A2(n_574), .B1(n_567), .B2(n_566), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_585), .A2(n_566), .B(n_548), .Y(n_639) );
OAI21xp33_ASAP7_75t_SL g640 ( .A1(n_624), .A2(n_538), .B(n_33), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_599), .Y(n_641) );
OAI221xp5_ASAP7_75t_SL g642 ( .A1(n_586), .A2(n_32), .B1(n_34), .B2(n_37), .C(n_39), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_624), .B(n_41), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_613), .Y(n_644) );
AOI21xp33_ASAP7_75t_SL g645 ( .A1(n_609), .A2(n_47), .B(n_48), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_584), .Y(n_646) );
AOI222xp33_ASAP7_75t_L g647 ( .A1(n_605), .A2(n_49), .B1(n_51), .B2(n_52), .C1(n_53), .C2(n_54), .Y(n_647) );
NAND2x1_ASAP7_75t_L g648 ( .A(n_586), .B(n_94), .Y(n_648) );
AOI211xp5_ASAP7_75t_L g649 ( .A1(n_610), .A2(n_58), .B(n_60), .C(n_63), .Y(n_649) );
NOR3xp33_ASAP7_75t_L g650 ( .A(n_595), .B(n_64), .C(n_65), .Y(n_650) );
NOR4xp25_ASAP7_75t_L g651 ( .A(n_622), .B(n_66), .C(n_70), .D(n_71), .Y(n_651) );
O2A1O1Ixp5_ASAP7_75t_L g652 ( .A1(n_603), .A2(n_74), .B(n_75), .C(n_76), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_606), .B(n_78), .Y(n_653) );
AOI211xp5_ASAP7_75t_L g654 ( .A1(n_616), .A2(n_80), .B(n_81), .C(n_82), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_598), .Y(n_655) );
A2O1A1Ixp33_ASAP7_75t_L g656 ( .A1(n_618), .A2(n_84), .B(n_87), .C(n_90), .Y(n_656) );
NAND2xp5_ASAP7_75t_SL g657 ( .A(n_615), .B(n_601), .Y(n_657) );
O2A1O1Ixp33_ASAP7_75t_L g658 ( .A1(n_600), .A2(n_625), .B(n_614), .C(n_621), .Y(n_658) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_607), .A2(n_593), .B1(n_597), .B2(n_611), .C(n_612), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_604), .A2(n_619), .B1(n_620), .B2(n_601), .Y(n_660) );
OAI21xp33_ASAP7_75t_L g661 ( .A1(n_604), .A2(n_623), .B(n_588), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_582), .A2(n_579), .B1(n_624), .B2(n_586), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_644), .Y(n_663) );
AOI21xp33_ASAP7_75t_L g664 ( .A1(n_662), .A2(n_661), .B(n_634), .Y(n_664) );
OR2x2_ASAP7_75t_L g665 ( .A(n_628), .B(n_657), .Y(n_665) );
OAI211xp5_ASAP7_75t_SL g666 ( .A1(n_631), .A2(n_659), .B(n_629), .C(n_647), .Y(n_666) );
NAND4xp25_ASAP7_75t_L g667 ( .A(n_626), .B(n_647), .C(n_649), .D(n_656), .Y(n_667) );
NOR4xp25_ASAP7_75t_L g668 ( .A(n_638), .B(n_658), .C(n_642), .D(n_627), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_641), .Y(n_669) );
NOR3xp33_ASAP7_75t_L g670 ( .A(n_664), .B(n_640), .C(n_645), .Y(n_670) );
NAND4xp25_ASAP7_75t_L g671 ( .A(n_667), .B(n_649), .C(n_654), .D(n_652), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_665), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_663), .Y(n_673) );
AND4x1_ASAP7_75t_L g674 ( .A(n_670), .B(n_668), .C(n_651), .D(n_643), .Y(n_674) );
NOR2x1_ASAP7_75t_L g675 ( .A(n_671), .B(n_666), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_672), .A2(n_637), .B1(n_630), .B2(n_669), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_675), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_674), .B(n_673), .Y(n_678) );
INVxp67_ASAP7_75t_L g679 ( .A(n_678), .Y(n_679) );
XNOR2x1_ASAP7_75t_L g680 ( .A(n_677), .B(n_676), .Y(n_680) );
OAI22x1_ASAP7_75t_L g681 ( .A1(n_679), .A2(n_636), .B1(n_660), .B2(n_655), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_680), .B(n_633), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_682), .A2(n_648), .B(n_639), .Y(n_683) );
NAND3xp33_ASAP7_75t_L g684 ( .A(n_683), .B(n_681), .C(n_632), .Y(n_684) );
OR2x6_ASAP7_75t_L g685 ( .A(n_684), .B(n_646), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_685), .A2(n_653), .B1(n_635), .B2(n_650), .Y(n_686) );
endmodule