module fake_netlist_6_3610_n_1792 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1792);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1792;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_116),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_120),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_146),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_50),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_124),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_107),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_46),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_80),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_37),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_48),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_134),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_132),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_139),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_141),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_5),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_158),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_133),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_92),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_67),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_108),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_150),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_98),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_90),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_38),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_95),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_60),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_96),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_29),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_82),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_109),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_48),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_76),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_129),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_138),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_15),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_156),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_30),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_88),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

BUFx8_ASAP7_75t_SL g202 ( 
.A(n_101),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_24),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_32),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_12),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_144),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_13),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_36),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_41),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_145),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_71),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_19),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_74),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_93),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_152),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_52),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_121),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_52),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_44),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_7),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_56),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_3),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_16),
.Y(n_223)
);

BUFx10_ASAP7_75t_L g224 ( 
.A(n_22),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_24),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_62),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_73),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_135),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_32),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_28),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_64),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_126),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_75),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_29),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_97),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_143),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_102),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_11),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_15),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_6),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_81),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_50),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_119),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_45),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_103),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_127),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_70),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_128),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_37),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_151),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_30),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_38),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_58),
.Y(n_253)
);

INVxp33_ASAP7_75t_L g254 ( 
.A(n_35),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_6),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_100),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_79),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_12),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_112),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_148),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_41),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_94),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_83),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_89),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_7),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_155),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_57),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_131),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_42),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_0),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_13),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_31),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_21),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_9),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_0),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_14),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_3),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_61),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_99),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_57),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_58),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_142),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_154),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_105),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_17),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_160),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_19),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_56),
.Y(n_288)
);

INVxp67_ASAP7_75t_SL g289 ( 
.A(n_72),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_118),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_136),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_106),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_86),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_125),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_23),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_113),
.Y(n_296)
);

BUFx5_ASAP7_75t_L g297 ( 
.A(n_2),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_4),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_65),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_4),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_115),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_43),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_23),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_137),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_51),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_9),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_63),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_25),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_54),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_53),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_54),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_104),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_10),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_77),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_111),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_1),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_45),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_1),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_36),
.Y(n_319)
);

NOR2xp67_ASAP7_75t_L g320 ( 
.A(n_225),
.B(n_2),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_178),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_202),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_245),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_161),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_163),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_182),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_183),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_297),
.B(n_5),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_297),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_297),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_195),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_297),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_165),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_245),
.B(n_8),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_244),
.B(n_8),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_297),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_276),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_276),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_297),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_297),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_233),
.B(n_10),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_168),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_260),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_211),
.Y(n_344)
);

NOR2xp67_ASAP7_75t_L g345 ( 
.A(n_225),
.B(n_11),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_260),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_291),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_313),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_171),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_297),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_297),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_267),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_172),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_267),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_267),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_267),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_317),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_267),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_271),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_271),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_173),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_174),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_176),
.Y(n_363)
);

INVxp33_ASAP7_75t_SL g364 ( 
.A(n_170),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_180),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_271),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_184),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_271),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_271),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_167),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_240),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_232),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_189),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_192),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_240),
.Y(n_375)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_162),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_167),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_194),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_196),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_206),
.Y(n_380)
);

INVxp67_ASAP7_75t_SL g381 ( 
.A(n_162),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_232),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_210),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_212),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_232),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_213),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_166),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_212),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_232),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_214),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_215),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_234),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_313),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_175),
.Y(n_394)
);

NOR2xp67_ASAP7_75t_L g395 ( 
.A(n_234),
.B(n_14),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_329),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_357),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_352),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_352),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_347),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_354),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_385),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_320),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_354),
.Y(n_404)
);

BUFx8_ASAP7_75t_L g405 ( 
.A(n_394),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_385),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_355),
.Y(n_407)
);

INVx4_ASAP7_75t_L g408 ( 
.A(n_385),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_366),
.B(n_233),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_355),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_329),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_329),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_356),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_368),
.B(n_226),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_385),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_356),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_376),
.B(n_227),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_385),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_358),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_385),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_330),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_358),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_359),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_359),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_360),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_381),
.B(n_166),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_360),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_387),
.B(n_231),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_369),
.B(n_181),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_330),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_369),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_372),
.Y(n_432)
);

OR2x6_ASAP7_75t_L g433 ( 
.A(n_328),
.B(n_181),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_372),
.Y(n_434)
);

AND2x6_ASAP7_75t_L g435 ( 
.A(n_332),
.B(n_198),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_371),
.B(n_177),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_394),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_341),
.B(n_254),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_332),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_336),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_372),
.Y(n_441)
);

OA21x2_ASAP7_75t_L g442 ( 
.A1(n_328),
.A2(n_255),
.B(n_169),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_382),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_382),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_382),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_336),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_389),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_375),
.B(n_177),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_334),
.B(n_268),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_348),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_343),
.B(n_237),
.Y(n_451)
);

NAND3xp33_ASAP7_75t_L g452 ( 
.A(n_335),
.B(n_169),
.C(n_164),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_339),
.B(n_198),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_389),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_389),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_339),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_346),
.B(n_241),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_340),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_340),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_350),
.B(n_200),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_350),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_351),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_351),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_323),
.B(n_179),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_370),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_337),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_370),
.B(n_246),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_449),
.B(n_324),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_458),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_403),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_396),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_402),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_414),
.B(n_325),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_458),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_458),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_462),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_396),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_450),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_402),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g480 ( 
.A(n_403),
.Y(n_480)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_442),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_396),
.Y(n_482)
);

AND2x6_ASAP7_75t_L g483 ( 
.A(n_426),
.B(n_200),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_396),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_436),
.B(n_377),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_462),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_449),
.B(n_364),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_402),
.Y(n_488)
);

NAND2xp33_ASAP7_75t_L g489 ( 
.A(n_451),
.B(n_333),
.Y(n_489)
);

BUFx10_ASAP7_75t_L g490 ( 
.A(n_438),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_402),
.Y(n_491)
);

BUFx6f_ASAP7_75t_SL g492 ( 
.A(n_433),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_442),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_411),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_433),
.B(n_179),
.Y(n_495)
);

INVxp33_ASAP7_75t_L g496 ( 
.A(n_397),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_436),
.B(n_377),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_411),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_462),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_456),
.Y(n_500)
);

AO22x2_ASAP7_75t_L g501 ( 
.A1(n_452),
.A2(n_338),
.B1(n_252),
.B2(n_220),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_411),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_442),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_438),
.B(n_342),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_411),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_412),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_412),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_436),
.B(n_384),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_412),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_456),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_437),
.B(n_353),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_412),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_L g513 ( 
.A1(n_433),
.A2(n_338),
.B1(n_345),
.B2(n_320),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_433),
.A2(n_345),
.B1(n_395),
.B2(n_255),
.Y(n_514)
);

AND3x1_ASAP7_75t_L g515 ( 
.A(n_464),
.B(n_203),
.C(n_164),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_451),
.B(n_362),
.Y(n_516)
);

BUFx10_ASAP7_75t_L g517 ( 
.A(n_464),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_456),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_421),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_414),
.B(n_365),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_421),
.Y(n_521)
);

INVx4_ASAP7_75t_L g522 ( 
.A(n_442),
.Y(n_522)
);

OR2x6_ASAP7_75t_L g523 ( 
.A(n_433),
.B(n_185),
.Y(n_523)
);

NOR2x1p5_ASAP7_75t_L g524 ( 
.A(n_452),
.B(n_322),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_405),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_421),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_437),
.B(n_367),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_450),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_421),
.Y(n_529)
);

INVxp33_ASAP7_75t_SL g530 ( 
.A(n_400),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_402),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_457),
.B(n_373),
.Y(n_532)
);

OR2x6_ASAP7_75t_L g533 ( 
.A(n_433),
.B(n_185),
.Y(n_533)
);

OAI22xp33_ASAP7_75t_L g534 ( 
.A1(n_433),
.A2(n_300),
.B1(n_308),
.B2(n_253),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_456),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_457),
.B(n_374),
.Y(n_536)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_442),
.Y(n_537)
);

BUFx4f_ASAP7_75t_L g538 ( 
.A(n_442),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_448),
.B(n_384),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_453),
.Y(n_540)
);

BUFx4f_ASAP7_75t_L g541 ( 
.A(n_435),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_430),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_426),
.A2(n_448),
.B1(n_460),
.B2(n_453),
.Y(n_543)
);

BUFx10_ASAP7_75t_L g544 ( 
.A(n_397),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_430),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_426),
.A2(n_395),
.B1(n_269),
.B2(n_258),
.Y(n_546)
);

NAND2xp33_ASAP7_75t_L g547 ( 
.A(n_417),
.B(n_380),
.Y(n_547)
);

NOR3xp33_ASAP7_75t_L g548 ( 
.A(n_466),
.B(n_393),
.C(n_348),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_402),
.Y(n_549)
);

AND2x6_ASAP7_75t_L g550 ( 
.A(n_448),
.B(n_232),
.Y(n_550)
);

INVx4_ASAP7_75t_L g551 ( 
.A(n_453),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_461),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_430),
.Y(n_553)
);

INVx8_ASAP7_75t_L g554 ( 
.A(n_435),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_450),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_417),
.B(n_248),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_430),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_453),
.A2(n_272),
.B1(n_319),
.B2(n_318),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_466),
.A2(n_251),
.B1(n_270),
.B2(n_273),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_402),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_461),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_467),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_428),
.B(n_349),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_402),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_439),
.Y(n_565)
);

NAND2xp33_ASAP7_75t_L g566 ( 
.A(n_428),
.B(n_243),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_461),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_461),
.Y(n_568)
);

OR2x6_ASAP7_75t_L g569 ( 
.A(n_467),
.B(n_187),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_461),
.Y(n_570)
);

OR2x6_ASAP7_75t_L g571 ( 
.A(n_409),
.B(n_187),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_405),
.B(n_361),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_408),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_409),
.B(n_363),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_439),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_463),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_439),
.Y(n_577)
);

AND2x6_ASAP7_75t_L g578 ( 
.A(n_453),
.B(n_243),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_439),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_408),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_440),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_440),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_440),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g584 ( 
.A(n_400),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_440),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_446),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_405),
.B(n_378),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_405),
.B(n_379),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_453),
.B(n_188),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_463),
.Y(n_590)
);

BUFx4f_ASAP7_75t_L g591 ( 
.A(n_435),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_463),
.B(n_383),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_463),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_463),
.Y(n_594)
);

NAND3xp33_ASAP7_75t_L g595 ( 
.A(n_460),
.B(n_191),
.C(n_188),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_446),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_460),
.A2(n_203),
.B1(n_220),
.B2(n_252),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_460),
.A2(n_258),
.B1(n_269),
.B2(n_272),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_465),
.B(n_386),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_446),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_465),
.B(n_390),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_446),
.Y(n_602)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_460),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_459),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_459),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_460),
.A2(n_280),
.B1(n_190),
.B2(n_287),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_432),
.Y(n_607)
);

INVx4_ASAP7_75t_L g608 ( 
.A(n_432),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_459),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_459),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_404),
.Y(n_611)
);

AND3x2_ASAP7_75t_L g612 ( 
.A(n_429),
.B(n_393),
.C(n_201),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_405),
.Y(n_613)
);

AND3x2_ASAP7_75t_L g614 ( 
.A(n_429),
.B(n_201),
.C(n_191),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_404),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_404),
.Y(n_616)
);

AND3x2_ASAP7_75t_L g617 ( 
.A(n_429),
.B(n_235),
.C(n_217),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_398),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_487),
.B(n_391),
.Y(n_619)
);

OAI22xp33_ASAP7_75t_L g620 ( 
.A1(n_571),
.A2(n_319),
.B1(n_318),
.B2(n_309),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_526),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_541),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_544),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_555),
.B(n_321),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_538),
.B(n_405),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_516),
.B(n_562),
.Y(n_626)
);

NAND2xp33_ASAP7_75t_L g627 ( 
.A(n_483),
.B(n_250),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_526),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_618),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_618),
.Y(n_630)
);

INVxp67_ASAP7_75t_L g631 ( 
.A(n_478),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_470),
.B(n_186),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_470),
.B(n_193),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_493),
.A2(n_309),
.B1(n_288),
.B2(n_290),
.Y(n_634)
);

NAND2xp33_ASAP7_75t_L g635 ( 
.A(n_483),
.B(n_256),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_530),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_603),
.B(n_429),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_603),
.B(n_429),
.Y(n_638)
);

INVx4_ASAP7_75t_L g639 ( 
.A(n_540),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_555),
.B(n_326),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_478),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_543),
.A2(n_344),
.B1(n_331),
.B2(n_327),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_528),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_584),
.Y(n_644)
);

A2O1A1Ixp33_ASAP7_75t_L g645 ( 
.A1(n_538),
.A2(n_429),
.B(n_294),
.C(n_307),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_500),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_480),
.B(n_197),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_500),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_538),
.B(n_243),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_541),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_528),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_473),
.B(n_398),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_584),
.Y(n_653)
);

INVx8_ASAP7_75t_L g654 ( 
.A(n_483),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_520),
.B(n_399),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_490),
.B(n_257),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_526),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_510),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_540),
.Y(n_659)
);

INVxp67_ASAP7_75t_L g660 ( 
.A(n_599),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_471),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_541),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_471),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_532),
.B(n_536),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_556),
.B(n_510),
.Y(n_665)
);

OAI22x1_ASAP7_75t_SL g666 ( 
.A1(n_559),
.A2(n_204),
.B1(n_205),
.B2(n_199),
.Y(n_666)
);

OR2x2_ASAP7_75t_L g667 ( 
.A(n_480),
.B(n_207),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_490),
.B(n_208),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_540),
.B(n_243),
.Y(n_669)
);

OR2x6_ASAP7_75t_L g670 ( 
.A(n_572),
.B(n_587),
.Y(n_670)
);

NAND2xp33_ASAP7_75t_L g671 ( 
.A(n_483),
.B(n_259),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_540),
.B(n_243),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_518),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_551),
.B(n_262),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_551),
.B(n_263),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_490),
.B(n_209),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_485),
.B(n_217),
.Y(n_677)
);

INVxp33_ASAP7_75t_L g678 ( 
.A(n_496),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_518),
.B(n_399),
.Y(n_679)
);

INVx5_ASAP7_75t_L g680 ( 
.A(n_578),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_535),
.B(n_401),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_469),
.B(n_474),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_469),
.B(n_401),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g684 ( 
.A(n_601),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_493),
.A2(n_288),
.B1(n_286),
.B2(n_279),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_474),
.B(n_407),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_475),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_490),
.B(n_216),
.Y(n_688)
);

INVx4_ASAP7_75t_L g689 ( 
.A(n_551),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_476),
.B(n_486),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_544),
.Y(n_691)
);

NAND2x1_ASAP7_75t_L g692 ( 
.A(n_551),
.B(n_408),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_476),
.B(n_407),
.Y(n_693)
);

NAND3xp33_ASAP7_75t_L g694 ( 
.A(n_513),
.B(n_265),
.C(n_281),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_486),
.B(n_435),
.Y(n_695)
);

NAND2x1p5_ASAP7_75t_L g696 ( 
.A(n_613),
.B(n_228),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_504),
.B(n_218),
.Y(n_697)
);

NAND2xp33_ASAP7_75t_SL g698 ( 
.A(n_524),
.B(n_219),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_499),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_499),
.B(n_435),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_574),
.B(n_264),
.Y(n_701)
);

A2O1A1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_493),
.A2(n_495),
.B(n_514),
.C(n_589),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_477),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_485),
.B(n_435),
.Y(n_704)
);

INVx4_ASAP7_75t_L g705 ( 
.A(n_554),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_497),
.B(n_435),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_495),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_592),
.A2(n_289),
.B1(n_284),
.B2(n_283),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_497),
.B(n_224),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_517),
.B(n_221),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_495),
.B(n_266),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_495),
.B(n_278),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_508),
.B(n_435),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_477),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_611),
.Y(n_715)
);

NAND2xp33_ASAP7_75t_L g716 ( 
.A(n_483),
.B(n_282),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_611),
.Y(n_717)
);

A2O1A1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_589),
.A2(n_539),
.B(n_508),
.C(n_552),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_539),
.B(n_435),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_589),
.B(n_228),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_483),
.A2(n_293),
.B1(n_312),
.B2(n_301),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_483),
.B(n_435),
.Y(n_722)
);

NOR2xp67_ASAP7_75t_SL g723 ( 
.A(n_613),
.B(n_235),
.Y(n_723)
);

NAND2xp33_ASAP7_75t_L g724 ( 
.A(n_550),
.B(n_296),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_615),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_511),
.Y(n_726)
);

O2A1O1Ixp33_ASAP7_75t_L g727 ( 
.A1(n_571),
.A2(n_247),
.B(n_279),
.C(n_286),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_481),
.A2(n_307),
.B1(n_236),
.B2(n_290),
.Y(n_728)
);

BUFx6f_ASAP7_75t_SL g729 ( 
.A(n_544),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_569),
.B(n_435),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_482),
.Y(n_731)
);

AND2x4_ASAP7_75t_SL g732 ( 
.A(n_544),
.B(n_224),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_569),
.B(n_410),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_569),
.B(n_552),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_481),
.B(n_315),
.Y(n_735)
);

INVxp67_ASAP7_75t_SL g736 ( 
.A(n_573),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_517),
.B(n_548),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_468),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_481),
.B(n_236),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_517),
.B(n_222),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_591),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_559),
.B(n_606),
.Y(n_742)
);

INVxp67_ASAP7_75t_L g743 ( 
.A(n_527),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_482),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_569),
.B(n_410),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_481),
.B(n_247),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_591),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_484),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_615),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_503),
.B(n_292),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_569),
.B(n_561),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_561),
.B(n_410),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_567),
.B(n_413),
.Y(n_753)
);

NAND2x1p5_ASAP7_75t_L g754 ( 
.A(n_591),
.B(n_292),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_616),
.Y(n_755)
);

NOR2xp67_ASAP7_75t_L g756 ( 
.A(n_525),
.B(n_413),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_503),
.B(n_294),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_503),
.A2(n_299),
.B1(n_304),
.B2(n_314),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_517),
.B(n_299),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_484),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_534),
.B(n_563),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_503),
.B(n_223),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_606),
.B(n_304),
.Y(n_763)
);

NOR2xp67_ASAP7_75t_L g764 ( 
.A(n_525),
.B(n_595),
.Y(n_764)
);

INVxp67_ASAP7_75t_L g765 ( 
.A(n_515),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_515),
.B(n_314),
.Y(n_766)
);

AND2x2_ASAP7_75t_SL g767 ( 
.A(n_522),
.B(n_408),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_501),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_547),
.A2(n_413),
.B1(n_416),
.B2(n_419),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_616),
.Y(n_770)
);

INVx1_ASAP7_75t_SL g771 ( 
.A(n_612),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_571),
.B(n_224),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_494),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_494),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_522),
.B(n_408),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_522),
.B(n_229),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_522),
.B(n_432),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_568),
.B(n_416),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_537),
.B(n_230),
.Y(n_779)
);

AO22x2_ASAP7_75t_L g780 ( 
.A1(n_588),
.A2(n_388),
.B1(n_392),
.B2(n_416),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_498),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_568),
.B(n_419),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_571),
.B(n_261),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_537),
.B(n_238),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_589),
.B(n_524),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_554),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_660),
.B(n_537),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_707),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_749),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_664),
.B(n_537),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_626),
.B(n_546),
.Y(n_791)
);

INVx4_ASAP7_75t_L g792 ( 
.A(n_786),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_652),
.B(n_571),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_659),
.A2(n_580),
.B(n_573),
.Y(n_794)
);

AO21x1_ASAP7_75t_L g795 ( 
.A1(n_649),
.A2(n_566),
.B(n_489),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_707),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_659),
.A2(n_580),
.B(n_573),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_637),
.A2(n_580),
.B(n_573),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_644),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_655),
.B(n_570),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_684),
.B(n_576),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_638),
.A2(n_580),
.B(n_554),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_736),
.B(n_576),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_705),
.A2(n_775),
.B(n_777),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_705),
.A2(n_554),
.B(n_491),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_775),
.A2(n_554),
.B(n_491),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_777),
.A2(n_491),
.B(n_488),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_622),
.B(n_590),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_702),
.A2(n_492),
.B1(n_523),
.B2(n_533),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_728),
.A2(n_492),
.B1(n_523),
.B2(n_533),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_786),
.A2(n_491),
.B(n_488),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_786),
.A2(n_491),
.B(n_488),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_653),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_749),
.Y(n_814)
);

OR2x2_ASAP7_75t_L g815 ( 
.A(n_631),
.B(n_523),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_786),
.A2(n_649),
.B(n_622),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_622),
.B(n_590),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_687),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_622),
.A2(n_531),
.B(n_488),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_699),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_629),
.B(n_630),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_646),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_665),
.B(n_728),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_650),
.B(n_662),
.Y(n_824)
);

AOI21x1_ASAP7_75t_L g825 ( 
.A1(n_739),
.A2(n_594),
.B(n_593),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_758),
.B(n_593),
.Y(n_826)
);

O2A1O1Ixp33_ASAP7_75t_SL g827 ( 
.A1(n_718),
.A2(n_594),
.B(n_595),
.C(n_596),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_650),
.A2(n_531),
.B(n_488),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_758),
.B(n_550),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_685),
.B(n_550),
.Y(n_830)
);

CKINVDCx10_ASAP7_75t_R g831 ( 
.A(n_729),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_650),
.A2(n_741),
.B(n_662),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_648),
.Y(n_833)
);

OR2x2_ASAP7_75t_L g834 ( 
.A(n_643),
.B(n_523),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_L g835 ( 
.A1(n_739),
.A2(n_602),
.B(n_596),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_650),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_662),
.A2(n_549),
.B(n_531),
.Y(n_837)
);

O2A1O1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_768),
.A2(n_523),
.B(n_533),
.C(n_605),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_662),
.A2(n_549),
.B(n_531),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_685),
.B(n_550),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_762),
.A2(n_492),
.B1(n_533),
.B2(n_550),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_658),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_741),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_741),
.A2(n_549),
.B(n_531),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_639),
.Y(n_845)
);

O2A1O1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_763),
.A2(n_533),
.B(n_605),
.C(n_602),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_762),
.B(n_550),
.Y(n_847)
);

CKINVDCx20_ASAP7_75t_R g848 ( 
.A(n_636),
.Y(n_848)
);

BUFx2_ASAP7_75t_L g849 ( 
.A(n_641),
.Y(n_849)
);

O2A1O1Ixp33_ASAP7_75t_L g850 ( 
.A1(n_766),
.A2(n_558),
.B(n_597),
.C(n_598),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_738),
.B(n_549),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_R g852 ( 
.A(n_698),
.B(n_550),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_673),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_776),
.B(n_501),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_634),
.A2(n_501),
.B1(n_560),
.B2(n_564),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_741),
.A2(n_549),
.B(n_608),
.Y(n_856)
);

INVxp67_ASAP7_75t_L g857 ( 
.A(n_709),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_776),
.B(n_501),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_710),
.B(n_472),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_747),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_779),
.B(n_519),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_747),
.A2(n_608),
.B(n_607),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_747),
.A2(n_608),
.B(n_607),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_710),
.B(n_472),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_747),
.A2(n_608),
.B(n_607),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_779),
.B(n_519),
.Y(n_866)
);

BUFx8_ASAP7_75t_L g867 ( 
.A(n_729),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_651),
.Y(n_868)
);

O2A1O1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_765),
.A2(n_542),
.B(n_521),
.C(n_610),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_692),
.A2(n_607),
.B(n_560),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_784),
.B(n_521),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_639),
.A2(n_607),
.B(n_560),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_654),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_689),
.A2(n_479),
.B(n_560),
.Y(n_874)
);

NOR2x1_ASAP7_75t_L g875 ( 
.A(n_656),
.B(n_472),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_624),
.B(n_261),
.Y(n_876)
);

AO21x1_ASAP7_75t_L g877 ( 
.A1(n_735),
.A2(n_545),
.B(n_529),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_784),
.B(n_634),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_689),
.A2(n_479),
.B(n_564),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_654),
.A2(n_479),
.B(n_564),
.Y(n_880)
);

BUFx4f_ASAP7_75t_L g881 ( 
.A(n_670),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_654),
.A2(n_479),
.B(n_564),
.Y(n_882)
);

OAI321xp33_ASAP7_75t_L g883 ( 
.A1(n_761),
.A2(n_392),
.A3(n_388),
.B1(n_261),
.B2(n_431),
.C(n_419),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_632),
.B(n_529),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_746),
.A2(n_472),
.B(n_610),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_715),
.Y(n_886)
);

CKINVDCx20_ASAP7_75t_R g887 ( 
.A(n_642),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_632),
.B(n_542),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_746),
.A2(n_575),
.B(n_609),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_750),
.A2(n_757),
.B(n_706),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_750),
.A2(n_575),
.B(n_609),
.Y(n_891)
);

OAI21xp5_ASAP7_75t_L g892 ( 
.A1(n_757),
.A2(n_577),
.B(n_604),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_697),
.A2(n_578),
.B1(n_545),
.B2(n_604),
.Y(n_893)
);

OAI21xp5_ASAP7_75t_L g894 ( 
.A1(n_704),
.A2(n_577),
.B(n_600),
.Y(n_894)
);

INVx1_ASAP7_75t_SL g895 ( 
.A(n_640),
.Y(n_895)
);

O2A1O1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_759),
.A2(n_553),
.B(n_557),
.C(n_600),
.Y(n_896)
);

NOR2x1_ASAP7_75t_L g897 ( 
.A(n_737),
.B(n_553),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_767),
.B(n_557),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_633),
.B(n_565),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_667),
.Y(n_900)
);

AOI21x1_ASAP7_75t_L g901 ( 
.A1(n_669),
.A2(n_565),
.B(n_579),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_713),
.A2(n_579),
.B(n_586),
.Y(n_902)
);

OAI21xp5_ASAP7_75t_L g903 ( 
.A1(n_719),
.A2(n_581),
.B(n_586),
.Y(n_903)
);

O2A1O1Ixp33_ASAP7_75t_SL g904 ( 
.A1(n_645),
.A2(n_581),
.B(n_582),
.C(n_585),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_767),
.B(n_734),
.Y(n_905)
);

NAND3x1_ASAP7_75t_L g906 ( 
.A(n_619),
.B(n_249),
.C(n_316),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_785),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_717),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_751),
.B(n_582),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_725),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_633),
.B(n_583),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_647),
.B(n_239),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_680),
.B(n_583),
.Y(n_913)
);

INVxp67_ASAP7_75t_L g914 ( 
.A(n_647),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_627),
.A2(n_585),
.B(n_505),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_755),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_635),
.A2(n_506),
.B(n_502),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_740),
.B(n_498),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_671),
.A2(n_506),
.B(n_505),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_716),
.A2(n_735),
.B(n_690),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_682),
.A2(n_507),
.B(n_512),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_785),
.B(n_614),
.Y(n_922)
);

BUFx3_ASAP7_75t_L g923 ( 
.A(n_732),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_619),
.B(n_242),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_726),
.B(n_274),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_770),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_683),
.Y(n_927)
);

O2A1O1Ixp5_ASAP7_75t_L g928 ( 
.A1(n_669),
.A2(n_502),
.B(n_507),
.C(n_512),
.Y(n_928)
);

INVxp67_ASAP7_75t_L g929 ( 
.A(n_772),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_743),
.B(n_275),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_677),
.B(n_509),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_742),
.B(n_277),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_668),
.B(n_285),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_686),
.Y(n_934)
);

O2A1O1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_620),
.A2(n_509),
.B(n_422),
.C(n_423),
.Y(n_935)
);

BUFx4f_ASAP7_75t_L g936 ( 
.A(n_670),
.Y(n_936)
);

INVx4_ASAP7_75t_L g937 ( 
.A(n_680),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_674),
.A2(n_406),
.B(n_420),
.Y(n_938)
);

NAND3xp33_ASAP7_75t_L g939 ( 
.A(n_697),
.B(n_295),
.C(n_298),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_677),
.B(n_578),
.Y(n_940)
);

CKINVDCx20_ASAP7_75t_R g941 ( 
.A(n_623),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_740),
.A2(n_676),
.B1(n_668),
.B2(n_688),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_733),
.A2(n_578),
.B(n_415),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_674),
.A2(n_406),
.B(n_420),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_676),
.B(n_578),
.Y(n_945)
);

OAI21xp33_ASAP7_75t_L g946 ( 
.A1(n_688),
.A2(n_302),
.B(n_303),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_678),
.B(n_305),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_745),
.A2(n_427),
.B(n_422),
.C(n_423),
.Y(n_948)
);

O2A1O1Ixp5_ASAP7_75t_L g949 ( 
.A1(n_672),
.A2(n_427),
.B(n_423),
.C(n_424),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_621),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_696),
.A2(n_306),
.B1(n_310),
.B2(n_311),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_711),
.A2(n_578),
.B1(n_431),
.B2(n_422),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_691),
.B(n_708),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_720),
.B(n_578),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_694),
.B(n_16),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_628),
.Y(n_956)
);

O2A1O1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_620),
.A2(n_431),
.B(n_424),
.C(n_425),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_672),
.A2(n_418),
.B(n_415),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_783),
.B(n_617),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_693),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_679),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_675),
.A2(n_406),
.B(n_420),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_720),
.B(n_427),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_675),
.A2(n_406),
.B(n_420),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_680),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_696),
.A2(n_425),
.B1(n_424),
.B2(n_444),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_722),
.A2(n_406),
.B(n_420),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_695),
.A2(n_415),
.B(n_418),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_657),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_701),
.B(n_425),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_756),
.B(n_432),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_780),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_700),
.A2(n_443),
.B(n_441),
.C(n_445),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_780),
.B(n_455),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_780),
.B(n_455),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_927),
.B(n_681),
.Y(n_976)
);

CKINVDCx16_ASAP7_75t_R g977 ( 
.A(n_848),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_SL g978 ( 
.A1(n_878),
.A2(n_730),
.B(n_712),
.C(n_711),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_942),
.A2(n_670),
.B1(n_712),
.B2(n_764),
.Y(n_979)
);

AND2x2_ASAP7_75t_SL g980 ( 
.A(n_881),
.B(n_936),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_818),
.Y(n_981)
);

OAI22x1_ASAP7_75t_L g982 ( 
.A1(n_932),
.A2(n_666),
.B1(n_771),
.B2(n_625),
.Y(n_982)
);

BUFx2_ASAP7_75t_L g983 ( 
.A(n_799),
.Y(n_983)
);

BUFx8_ASAP7_75t_L g984 ( 
.A(n_849),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_950),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_R g986 ( 
.A(n_813),
.B(n_724),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_914),
.B(n_625),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_934),
.B(n_752),
.Y(n_988)
);

OAI21xp33_ASAP7_75t_L g989 ( 
.A1(n_932),
.A2(n_721),
.B(n_754),
.Y(n_989)
);

O2A1O1Ixp5_ASAP7_75t_L g990 ( 
.A1(n_795),
.A2(n_723),
.B(n_782),
.C(n_778),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_907),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_920),
.A2(n_680),
.B(n_754),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_790),
.A2(n_753),
.B(n_774),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_868),
.Y(n_994)
);

BUFx12f_ASAP7_75t_L g995 ( 
.A(n_867),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_914),
.B(n_769),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_798),
.A2(n_781),
.B(n_773),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_956),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_833),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_804),
.A2(n_760),
.B(n_748),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_955),
.A2(n_727),
.B(n_731),
.C(n_744),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_823),
.A2(n_714),
.B1(n_703),
.B2(n_663),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_960),
.B(n_661),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_924),
.B(n_17),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_857),
.B(n_900),
.Y(n_1005)
);

OAI21x1_ASAP7_75t_L g1006 ( 
.A1(n_917),
.A2(n_415),
.B(n_418),
.Y(n_1006)
);

INVxp67_ASAP7_75t_L g1007 ( 
.A(n_868),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_836),
.Y(n_1008)
);

INVxp67_ASAP7_75t_L g1009 ( 
.A(n_947),
.Y(n_1009)
);

OR2x6_ASAP7_75t_L g1010 ( 
.A(n_923),
.B(n_418),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_961),
.B(n_444),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_SL g1012 ( 
.A(n_810),
.B(n_66),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_854),
.A2(n_443),
.B1(n_441),
.B2(n_445),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_794),
.A2(n_434),
.B(n_432),
.Y(n_1014)
);

NOR2x1_ASAP7_75t_L g1015 ( 
.A(n_793),
.B(n_447),
.Y(n_1015)
);

OAI21xp33_ASAP7_75t_L g1016 ( 
.A1(n_925),
.A2(n_447),
.B(n_454),
.Y(n_1016)
);

NOR3xp33_ASAP7_75t_SL g1017 ( 
.A(n_946),
.B(n_447),
.C(n_20),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_929),
.Y(n_1018)
);

OAI21xp33_ASAP7_75t_SL g1019 ( 
.A1(n_826),
.A2(n_455),
.B(n_454),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_912),
.B(n_18),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_858),
.A2(n_455),
.B1(n_454),
.B2(n_434),
.Y(n_1021)
);

INVx2_ASAP7_75t_SL g1022 ( 
.A(n_895),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_857),
.B(n_887),
.Y(n_1023)
);

NOR3xp33_ASAP7_75t_L g1024 ( 
.A(n_929),
.B(n_455),
.C(n_454),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_933),
.B(n_434),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_941),
.Y(n_1026)
);

A2O1A1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_955),
.A2(n_454),
.B(n_434),
.C(n_432),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_797),
.A2(n_434),
.B(n_432),
.Y(n_1028)
);

BUFx8_ASAP7_75t_L g1029 ( 
.A(n_959),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_972),
.A2(n_881),
.B1(n_936),
.B2(n_830),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_907),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_969),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_802),
.A2(n_434),
.B(n_432),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_800),
.B(n_434),
.Y(n_1034)
);

O2A1O1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_791),
.A2(n_18),
.B(n_20),
.C(n_21),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_907),
.B(n_434),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_816),
.A2(n_157),
.B(n_149),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_972),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_1038)
);

INVx3_ASAP7_75t_SL g1039 ( 
.A(n_922),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_907),
.B(n_147),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_831),
.Y(n_1041)
);

AOI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_953),
.A2(n_140),
.B1(n_123),
.B2(n_122),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_925),
.B(n_26),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_820),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_838),
.A2(n_27),
.B(n_28),
.C(n_31),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_846),
.A2(n_27),
.B(n_33),
.C(n_34),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_850),
.A2(n_33),
.B(n_34),
.C(n_35),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_930),
.B(n_39),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_876),
.B(n_930),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_861),
.A2(n_59),
.B(n_114),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_836),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_836),
.B(n_117),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_867),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_788),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_796),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_787),
.B(n_110),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_801),
.B(n_39),
.Y(n_1057)
);

NAND2x1p5_ASAP7_75t_L g1058 ( 
.A(n_836),
.B(n_91),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_866),
.A2(n_87),
.B(n_85),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_787),
.B(n_801),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_871),
.A2(n_84),
.B(n_78),
.Y(n_1061)
);

AOI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_939),
.A2(n_69),
.B1(n_68),
.B2(n_43),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_843),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_805),
.A2(n_55),
.B(n_42),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_806),
.A2(n_40),
.B(n_44),
.Y(n_1065)
);

AO21x1_ASAP7_75t_L g1066 ( 
.A1(n_905),
.A2(n_40),
.B(n_46),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_884),
.B(n_47),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_832),
.A2(n_55),
.B(n_49),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_843),
.B(n_47),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_888),
.B(n_49),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_815),
.B(n_51),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_843),
.B(n_53),
.Y(n_1072)
);

O2A1O1Ixp5_ASAP7_75t_L g1073 ( 
.A1(n_847),
.A2(n_877),
.B(n_864),
.C(n_859),
.Y(n_1073)
);

OAI21xp33_ASAP7_75t_L g1074 ( 
.A1(n_951),
.A2(n_821),
.B(n_834),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_905),
.A2(n_851),
.B(n_963),
.C(n_948),
.Y(n_1075)
);

AOI21x1_ASAP7_75t_L g1076 ( 
.A1(n_898),
.A2(n_909),
.B(n_817),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_822),
.B(n_842),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_922),
.B(n_853),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_897),
.A2(n_886),
.B1(n_809),
.B2(n_908),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_789),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_937),
.A2(n_856),
.B(n_898),
.Y(n_1081)
);

BUFx2_ASAP7_75t_L g1082 ( 
.A(n_906),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_937),
.A2(n_865),
.B(n_862),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_SL g1084 ( 
.A(n_792),
.B(n_873),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_843),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_899),
.B(n_911),
.Y(n_1086)
);

OAI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_840),
.A2(n_829),
.B1(n_841),
.B2(n_855),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_860),
.A2(n_803),
.B1(n_890),
.B2(n_931),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_860),
.B(n_845),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_910),
.B(n_916),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_926),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_863),
.A2(n_839),
.B(n_837),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_860),
.Y(n_1093)
);

O2A1O1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_883),
.A2(n_918),
.B(n_827),
.C(n_970),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_860),
.B(n_845),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_873),
.B(n_792),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_814),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_873),
.A2(n_975),
.B1(n_974),
.B2(n_824),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_814),
.B(n_824),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_945),
.A2(n_943),
.B(n_869),
.C(n_940),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_L g1101 ( 
.A1(n_954),
.A2(n_909),
.B1(n_875),
.B2(n_817),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_808),
.B(n_921),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_819),
.A2(n_828),
.B(n_844),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_893),
.B(n_952),
.Y(n_1104)
);

NOR2x1_ASAP7_75t_L g1105 ( 
.A(n_808),
.B(n_913),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_R g1106 ( 
.A(n_873),
.B(n_825),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_965),
.B(n_852),
.Y(n_1107)
);

INVx4_ASAP7_75t_L g1108 ( 
.A(n_965),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_811),
.A2(n_812),
.B(n_882),
.Y(n_1109)
);

NOR3xp33_ASAP7_75t_SL g1110 ( 
.A(n_913),
.B(n_957),
.C(n_966),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_965),
.B(n_852),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_901),
.Y(n_1112)
);

O2A1O1Ixp5_ASAP7_75t_L g1113 ( 
.A1(n_971),
.A2(n_949),
.B(n_915),
.C(n_928),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_965),
.B(n_903),
.Y(n_1114)
);

AND2x6_ASAP7_75t_L g1115 ( 
.A(n_928),
.B(n_904),
.Y(n_1115)
);

OR2x2_ASAP7_75t_L g1116 ( 
.A(n_894),
.B(n_902),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_935),
.B(n_835),
.Y(n_1117)
);

INVx6_ASAP7_75t_L g1118 ( 
.A(n_896),
.Y(n_1118)
);

BUFx3_ASAP7_75t_L g1119 ( 
.A(n_967),
.Y(n_1119)
);

BUFx12f_ASAP7_75t_L g1120 ( 
.A(n_973),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_919),
.A2(n_807),
.B(n_891),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_892),
.Y(n_1122)
);

INVx4_ASAP7_75t_L g1123 ( 
.A(n_880),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_874),
.B(n_879),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_872),
.A2(n_870),
.B(n_968),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_949),
.Y(n_1126)
);

NOR3xp33_ASAP7_75t_SL g1127 ( 
.A(n_964),
.B(n_938),
.C(n_944),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1125),
.A2(n_885),
.B(n_889),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_1109),
.A2(n_962),
.B(n_958),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_992),
.A2(n_1086),
.B(n_1116),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1103),
.A2(n_1092),
.B(n_1006),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_989),
.A2(n_1083),
.B(n_1124),
.Y(n_1132)
);

CKINVDCx11_ASAP7_75t_R g1133 ( 
.A(n_995),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_1060),
.A2(n_976),
.B1(n_988),
.B2(n_979),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_1033),
.A2(n_1121),
.B(n_1081),
.Y(n_1135)
);

OAI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1087),
.A2(n_1100),
.B(n_1073),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_1049),
.B(n_1023),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_981),
.Y(n_1138)
);

AO31x2_ASAP7_75t_L g1139 ( 
.A1(n_1087),
.A2(n_1027),
.A3(n_1030),
.B(n_1088),
.Y(n_1139)
);

AO31x2_ASAP7_75t_L g1140 ( 
.A1(n_1030),
.A2(n_1088),
.A3(n_1098),
.B(n_1021),
.Y(n_1140)
);

AO31x2_ASAP7_75t_L g1141 ( 
.A1(n_1098),
.A2(n_1021),
.A3(n_1066),
.B(n_1126),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1019),
.A2(n_990),
.B(n_1094),
.Y(n_1142)
);

OAI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_987),
.A2(n_1102),
.B(n_1056),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_1043),
.A2(n_1048),
.B(n_1004),
.C(n_1012),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_976),
.B(n_988),
.Y(n_1145)
);

AOI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1114),
.A2(n_1056),
.B(n_1076),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1000),
.A2(n_997),
.B(n_1014),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_999),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_977),
.Y(n_1149)
);

INVxp67_ASAP7_75t_L g1150 ( 
.A(n_994),
.Y(n_1150)
);

BUFx4f_ASAP7_75t_L g1151 ( 
.A(n_980),
.Y(n_1151)
);

CKINVDCx20_ASAP7_75t_R g1152 ( 
.A(n_984),
.Y(n_1152)
);

AO31x2_ASAP7_75t_L g1153 ( 
.A1(n_1013),
.A2(n_1047),
.A3(n_1046),
.B(n_1002),
.Y(n_1153)
);

BUFx12f_ASAP7_75t_L g1154 ( 
.A(n_984),
.Y(n_1154)
);

AOI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1067),
.A2(n_1070),
.B(n_1025),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1028),
.A2(n_1112),
.B(n_1113),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1012),
.A2(n_1009),
.B1(n_982),
.B2(n_1074),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_983),
.Y(n_1158)
);

AOI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1078),
.A2(n_1020),
.B1(n_1082),
.B2(n_1077),
.Y(n_1159)
);

BUFx10_ASAP7_75t_L g1160 ( 
.A(n_1041),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1078),
.B(n_1018),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_1022),
.Y(n_1162)
);

A2O1A1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_1075),
.A2(n_1057),
.B(n_996),
.C(n_1001),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1002),
.A2(n_993),
.B(n_1034),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_1007),
.B(n_1005),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_993),
.A2(n_1034),
.B(n_1101),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_SL g1167 ( 
.A1(n_1053),
.A2(n_1038),
.B1(n_1039),
.B2(n_1026),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1003),
.B(n_1067),
.Y(n_1168)
);

BUFx4f_ASAP7_75t_L g1169 ( 
.A(n_991),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1071),
.B(n_1054),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1045),
.A2(n_1035),
.B(n_1038),
.C(n_978),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1070),
.A2(n_1065),
.B(n_1042),
.C(n_1104),
.Y(n_1172)
);

OA21x2_ASAP7_75t_L g1173 ( 
.A1(n_1117),
.A2(n_1122),
.B(n_1016),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1105),
.A2(n_1037),
.B(n_1079),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1090),
.B(n_1044),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_SL g1176 ( 
.A1(n_1052),
.A2(n_1040),
.B(n_1069),
.C(n_1072),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1123),
.A2(n_1084),
.B(n_1111),
.Y(n_1177)
);

O2A1O1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1017),
.A2(n_1068),
.B(n_1064),
.C(n_1091),
.Y(n_1178)
);

OR2x2_ASAP7_75t_L g1179 ( 
.A(n_1055),
.B(n_985),
.Y(n_1179)
);

AOI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1120),
.A2(n_1029),
.B1(n_1099),
.B2(n_998),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1123),
.A2(n_1084),
.B(n_1107),
.Y(n_1181)
);

NOR4xp25_ASAP7_75t_L g1182 ( 
.A(n_1013),
.B(n_1011),
.C(n_1097),
.D(n_1036),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1089),
.A2(n_1095),
.B(n_1119),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1050),
.A2(n_1061),
.B(n_1059),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_1080),
.B(n_1032),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1110),
.A2(n_1062),
.B1(n_1118),
.B2(n_1058),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1015),
.A2(n_1058),
.B(n_1063),
.Y(n_1187)
);

NOR2x1_ASAP7_75t_R g1188 ( 
.A(n_991),
.B(n_1031),
.Y(n_1188)
);

AO31x2_ASAP7_75t_L g1189 ( 
.A1(n_1115),
.A2(n_1127),
.A3(n_1108),
.B(n_1118),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_986),
.B(n_991),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1118),
.A2(n_1031),
.B1(n_1085),
.B2(n_1051),
.Y(n_1191)
);

NOR4xp25_ASAP7_75t_L g1192 ( 
.A(n_1008),
.B(n_1063),
.C(n_1024),
.D(n_1115),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1031),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1096),
.A2(n_1108),
.B(n_1008),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_SL g1195 ( 
.A1(n_1096),
.A2(n_1051),
.B(n_1085),
.Y(n_1195)
);

INVx3_ASAP7_75t_L g1196 ( 
.A(n_1085),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1093),
.B(n_1115),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1010),
.Y(n_1198)
);

OA21x2_ASAP7_75t_L g1199 ( 
.A1(n_1115),
.A2(n_1106),
.B(n_1010),
.Y(n_1199)
);

AO31x2_ASAP7_75t_L g1200 ( 
.A1(n_1010),
.A2(n_877),
.A3(n_795),
.B(n_1087),
.Y(n_1200)
);

AOI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1029),
.A2(n_920),
.B(n_1114),
.Y(n_1201)
);

OA21x2_ASAP7_75t_L g1202 ( 
.A1(n_1073),
.A2(n_1113),
.B(n_990),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1060),
.B(n_976),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_984),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1060),
.A2(n_728),
.B1(n_758),
.B2(n_685),
.Y(n_1205)
);

INVx1_ASAP7_75t_SL g1206 ( 
.A(n_994),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_SL g1207 ( 
.A1(n_1066),
.A2(n_838),
.B(n_1075),
.Y(n_1207)
);

O2A1O1Ixp33_ASAP7_75t_SL g1208 ( 
.A1(n_1046),
.A2(n_878),
.B(n_1047),
.C(n_858),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1060),
.B(n_976),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1049),
.B(n_932),
.Y(n_1210)
);

OA21x2_ASAP7_75t_L g1211 ( 
.A1(n_1073),
.A2(n_1113),
.B(n_990),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1060),
.B(n_976),
.Y(n_1212)
);

A2O1A1Ixp33_ASAP7_75t_L g1213 ( 
.A1(n_1043),
.A2(n_942),
.B(n_1048),
.C(n_1004),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1125),
.A2(n_920),
.B(n_659),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1060),
.B(n_976),
.Y(n_1215)
);

HB1xp67_ASAP7_75t_L g1216 ( 
.A(n_994),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1125),
.A2(n_920),
.B(n_659),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_1049),
.B(n_653),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1087),
.A2(n_878),
.B(n_1100),
.Y(n_1219)
);

OR2x2_ASAP7_75t_L g1220 ( 
.A(n_1022),
.B(n_642),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1109),
.A2(n_1103),
.B(n_1092),
.Y(n_1221)
);

OAI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1012),
.A2(n_942),
.B1(n_660),
.B2(n_684),
.Y(n_1222)
);

OR2x6_ASAP7_75t_L g1223 ( 
.A(n_983),
.B(n_991),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_977),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_981),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_981),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1125),
.A2(n_920),
.B(n_659),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_977),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1125),
.A2(n_920),
.B(n_659),
.Y(n_1229)
);

AOI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1043),
.A2(n_619),
.B1(n_942),
.B2(n_887),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1060),
.A2(n_728),
.B1(n_758),
.B2(n_685),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1125),
.A2(n_920),
.B(n_659),
.Y(n_1232)
);

OAI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1087),
.A2(n_878),
.B(n_1100),
.Y(n_1233)
);

AOI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1114),
.A2(n_920),
.B(n_1125),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1060),
.A2(n_728),
.B1(n_758),
.B2(n_685),
.Y(n_1235)
);

NAND3xp33_ASAP7_75t_L g1236 ( 
.A(n_1043),
.B(n_942),
.C(n_1048),
.Y(n_1236)
);

AO21x2_ASAP7_75t_L g1237 ( 
.A1(n_1125),
.A2(n_920),
.B(n_1103),
.Y(n_1237)
);

AO21x2_ASAP7_75t_L g1238 ( 
.A1(n_1125),
.A2(n_920),
.B(n_1103),
.Y(n_1238)
);

AOI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1114),
.A2(n_920),
.B(n_1125),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1109),
.A2(n_1103),
.B(n_1092),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1087),
.A2(n_877),
.A3(n_795),
.B(n_1027),
.Y(n_1241)
);

AO31x2_ASAP7_75t_L g1242 ( 
.A1(n_1087),
.A2(n_877),
.A3(n_795),
.B(n_1027),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1109),
.A2(n_1103),
.B(n_1092),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1109),
.A2(n_1103),
.B(n_1092),
.Y(n_1244)
);

NAND3x1_ASAP7_75t_L g1245 ( 
.A(n_1043),
.B(n_619),
.C(n_1048),
.Y(n_1245)
);

CKINVDCx20_ASAP7_75t_R g1246 ( 
.A(n_977),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1108),
.Y(n_1247)
);

CKINVDCx20_ASAP7_75t_R g1248 ( 
.A(n_977),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_981),
.Y(n_1249)
);

AND2x4_ASAP7_75t_L g1250 ( 
.A(n_1078),
.B(n_907),
.Y(n_1250)
);

NOR2xp67_ASAP7_75t_L g1251 ( 
.A(n_1009),
.B(n_813),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1051),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1049),
.B(n_660),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_984),
.Y(n_1254)
);

O2A1O1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1043),
.A2(n_1048),
.B(n_660),
.C(n_684),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_977),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1109),
.A2(n_1103),
.B(n_1092),
.Y(n_1257)
);

A2O1A1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1043),
.A2(n_942),
.B(n_1048),
.C(n_1004),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1049),
.B(n_932),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1060),
.B(n_626),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1109),
.A2(n_1103),
.B(n_1092),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1125),
.A2(n_920),
.B(n_659),
.Y(n_1262)
);

BUFx12f_ASAP7_75t_L g1263 ( 
.A(n_995),
.Y(n_1263)
);

AOI221x1_ASAP7_75t_L g1264 ( 
.A1(n_1043),
.A2(n_1048),
.B1(n_1047),
.B2(n_1030),
.C(n_1046),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_984),
.Y(n_1265)
);

A2O1A1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_1043),
.A2(n_942),
.B(n_1048),
.C(n_1004),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1060),
.B(n_976),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1109),
.A2(n_1103),
.B(n_1092),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1060),
.B(n_976),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1060),
.B(n_626),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1125),
.A2(n_920),
.B(n_659),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1125),
.A2(n_920),
.B(n_659),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1060),
.A2(n_728),
.B1(n_758),
.B2(n_685),
.Y(n_1273)
);

AOI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1043),
.A2(n_619),
.B1(n_942),
.B2(n_887),
.Y(n_1274)
);

OR2x2_ASAP7_75t_L g1275 ( 
.A(n_1022),
.B(n_642),
.Y(n_1275)
);

CKINVDCx11_ASAP7_75t_R g1276 ( 
.A(n_1160),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1230),
.A2(n_1274),
.B1(n_1245),
.B2(n_1144),
.Y(n_1277)
);

INVx4_ASAP7_75t_L g1278 ( 
.A(n_1169),
.Y(n_1278)
);

AOI22xp5_ASAP7_75t_SL g1279 ( 
.A1(n_1137),
.A2(n_1260),
.B1(n_1270),
.B2(n_1210),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1158),
.Y(n_1280)
);

CKINVDCx20_ASAP7_75t_R g1281 ( 
.A(n_1149),
.Y(n_1281)
);

CKINVDCx11_ASAP7_75t_R g1282 ( 
.A(n_1160),
.Y(n_1282)
);

CKINVDCx20_ASAP7_75t_R g1283 ( 
.A(n_1246),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1213),
.A2(n_1258),
.B1(n_1266),
.B2(n_1236),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1236),
.A2(n_1222),
.B1(n_1273),
.B2(n_1231),
.Y(n_1285)
);

BUFx12f_ASAP7_75t_L g1286 ( 
.A(n_1133),
.Y(n_1286)
);

INVx6_ASAP7_75t_L g1287 ( 
.A(n_1223),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_SL g1288 ( 
.A1(n_1205),
.A2(n_1231),
.B1(n_1273),
.B2(n_1235),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1138),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_1190),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_1224),
.Y(n_1291)
);

INVxp67_ASAP7_75t_SL g1292 ( 
.A(n_1145),
.Y(n_1292)
);

INVx1_ASAP7_75t_SL g1293 ( 
.A(n_1206),
.Y(n_1293)
);

AOI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1259),
.A2(n_1253),
.B1(n_1157),
.B2(n_1218),
.Y(n_1294)
);

INVx5_ASAP7_75t_L g1295 ( 
.A(n_1252),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1205),
.A2(n_1235),
.B1(n_1134),
.B2(n_1219),
.Y(n_1296)
);

NAND2x1p5_ASAP7_75t_L g1297 ( 
.A(n_1151),
.B(n_1247),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_SL g1298 ( 
.A1(n_1186),
.A2(n_1136),
.B1(n_1167),
.B2(n_1134),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1203),
.B(n_1209),
.Y(n_1299)
);

OAI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1255),
.A2(n_1163),
.B(n_1172),
.Y(n_1300)
);

BUFx8_ASAP7_75t_L g1301 ( 
.A(n_1263),
.Y(n_1301)
);

INVx6_ASAP7_75t_L g1302 ( 
.A(n_1223),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1186),
.A2(n_1219),
.B1(n_1233),
.B2(n_1220),
.Y(n_1303)
);

BUFx4f_ASAP7_75t_SL g1304 ( 
.A(n_1154),
.Y(n_1304)
);

INVx8_ASAP7_75t_L g1305 ( 
.A(n_1223),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1233),
.A2(n_1275),
.B1(n_1159),
.B2(n_1151),
.Y(n_1306)
);

INVx6_ASAP7_75t_L g1307 ( 
.A(n_1161),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1161),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1203),
.B(n_1209),
.Y(n_1309)
);

OAI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1212),
.A2(n_1269),
.B1(n_1215),
.B2(n_1267),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1212),
.A2(n_1269),
.B1(n_1215),
.B2(n_1267),
.Y(n_1311)
);

INVx6_ASAP7_75t_L g1312 ( 
.A(n_1252),
.Y(n_1312)
);

BUFx10_ASAP7_75t_L g1313 ( 
.A(n_1228),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1145),
.A2(n_1170),
.B1(n_1251),
.B2(n_1165),
.Y(n_1314)
);

NAND2x1p5_ASAP7_75t_L g1315 ( 
.A(n_1247),
.B(n_1169),
.Y(n_1315)
);

BUFx8_ASAP7_75t_SL g1316 ( 
.A(n_1248),
.Y(n_1316)
);

CKINVDCx6p67_ASAP7_75t_R g1317 ( 
.A(n_1152),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_SL g1318 ( 
.A1(n_1264),
.A2(n_1180),
.B(n_1171),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1168),
.B(n_1175),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_SL g1320 ( 
.A1(n_1136),
.A2(n_1143),
.B1(n_1207),
.B2(n_1168),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1206),
.B(n_1162),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_SL g1322 ( 
.A1(n_1256),
.A2(n_1265),
.B1(n_1204),
.B2(n_1254),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1143),
.A2(n_1249),
.B1(n_1226),
.B2(n_1225),
.Y(n_1323)
);

BUFx10_ASAP7_75t_L g1324 ( 
.A(n_1216),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1179),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1185),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1132),
.A2(n_1142),
.B1(n_1173),
.B2(n_1250),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1252),
.Y(n_1328)
);

INVx11_ASAP7_75t_L g1329 ( 
.A(n_1188),
.Y(n_1329)
);

INVx6_ASAP7_75t_L g1330 ( 
.A(n_1250),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_1193),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1196),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1142),
.A2(n_1173),
.B1(n_1130),
.B2(n_1198),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_SL g1334 ( 
.A1(n_1199),
.A2(n_1202),
.B1(n_1211),
.B2(n_1174),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1155),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1197),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_1150),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1178),
.B(n_1176),
.Y(n_1338)
);

BUFx8_ASAP7_75t_L g1339 ( 
.A(n_1195),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1197),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1191),
.A2(n_1199),
.B1(n_1181),
.B2(n_1177),
.Y(n_1341)
);

INVx6_ASAP7_75t_L g1342 ( 
.A(n_1191),
.Y(n_1342)
);

INVx1_ASAP7_75t_SL g1343 ( 
.A(n_1194),
.Y(n_1343)
);

CKINVDCx11_ASAP7_75t_R g1344 ( 
.A(n_1201),
.Y(n_1344)
);

OAI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1183),
.A2(n_1211),
.B1(n_1202),
.B2(n_1184),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_1237),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1208),
.B(n_1189),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_SL g1348 ( 
.A1(n_1166),
.A2(n_1237),
.B1(n_1238),
.B2(n_1140),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1272),
.A2(n_1217),
.B(n_1262),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1187),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1156),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1141),
.Y(n_1352)
);

BUFx10_ASAP7_75t_L g1353 ( 
.A(n_1192),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1200),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1139),
.B(n_1140),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1238),
.A2(n_1164),
.B1(n_1232),
.B2(n_1229),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1182),
.A2(n_1192),
.B1(n_1227),
.B2(n_1214),
.Y(n_1357)
);

INVx1_ASAP7_75t_SL g1358 ( 
.A(n_1128),
.Y(n_1358)
);

OAI21xp5_ASAP7_75t_SL g1359 ( 
.A1(n_1271),
.A2(n_1234),
.B(n_1239),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1182),
.B(n_1139),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_1139),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1129),
.A2(n_1221),
.B1(n_1261),
.B2(n_1257),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1200),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_1146),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1240),
.A2(n_1268),
.B1(n_1244),
.B2(n_1243),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1241),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_SL g1367 ( 
.A1(n_1153),
.A2(n_1135),
.B1(n_1147),
.B2(n_1241),
.Y(n_1367)
);

BUFx4f_ASAP7_75t_L g1368 ( 
.A(n_1153),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1153),
.B(n_1241),
.Y(n_1369)
);

OAI22x1_ASAP7_75t_L g1370 ( 
.A1(n_1242),
.A2(n_1230),
.B1(n_1274),
.B2(n_1236),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1242),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1131),
.A2(n_1236),
.B1(n_1274),
.B2(n_1230),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1242),
.Y(n_1373)
);

INVx3_ASAP7_75t_SL g1374 ( 
.A(n_1224),
.Y(n_1374)
);

BUFx4f_ASAP7_75t_SL g1375 ( 
.A(n_1263),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1230),
.A2(n_1274),
.B1(n_1245),
.B2(n_1144),
.Y(n_1376)
);

CKINVDCx10_ASAP7_75t_R g1377 ( 
.A(n_1133),
.Y(n_1377)
);

BUFx12f_ASAP7_75t_L g1378 ( 
.A(n_1133),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_SL g1379 ( 
.A1(n_1205),
.A2(n_1235),
.B1(n_1273),
.B2(n_1231),
.Y(n_1379)
);

OAI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1230),
.A2(n_1274),
.B1(n_1205),
.B2(n_1231),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_SL g1381 ( 
.A1(n_1205),
.A2(n_1235),
.B1(n_1273),
.B2(n_1231),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1247),
.Y(n_1382)
);

BUFx5_ASAP7_75t_L g1383 ( 
.A(n_1138),
.Y(n_1383)
);

OAI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1230),
.A2(n_1274),
.B1(n_1205),
.B2(n_1231),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_SL g1385 ( 
.A1(n_1205),
.A2(n_1235),
.B1(n_1273),
.B2(n_1231),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_SL g1386 ( 
.A1(n_1205),
.A2(n_1235),
.B1(n_1273),
.B2(n_1231),
.Y(n_1386)
);

CKINVDCx11_ASAP7_75t_R g1387 ( 
.A(n_1160),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1236),
.A2(n_1274),
.B1(n_1230),
.B2(n_1043),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1236),
.A2(n_1274),
.B1(n_1230),
.B2(n_1043),
.Y(n_1389)
);

INVx8_ASAP7_75t_L g1390 ( 
.A(n_1223),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1148),
.Y(n_1391)
);

CKINVDCx11_ASAP7_75t_R g1392 ( 
.A(n_1160),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1236),
.A2(n_1274),
.B1(n_1230),
.B2(n_1043),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1247),
.Y(n_1394)
);

CKINVDCx20_ASAP7_75t_R g1395 ( 
.A(n_1149),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_SL g1396 ( 
.A1(n_1205),
.A2(n_1235),
.B1(n_1273),
.B2(n_1231),
.Y(n_1396)
);

INVxp67_ASAP7_75t_L g1397 ( 
.A(n_1321),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1371),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1355),
.B(n_1288),
.Y(n_1399)
);

INVx3_ASAP7_75t_L g1400 ( 
.A(n_1369),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1288),
.B(n_1379),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1373),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1350),
.B(n_1369),
.Y(n_1403)
);

AO21x2_ASAP7_75t_L g1404 ( 
.A1(n_1345),
.A2(n_1349),
.B(n_1359),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1383),
.Y(n_1405)
);

AO32x1_ASAP7_75t_L g1406 ( 
.A1(n_1284),
.A2(n_1341),
.A3(n_1352),
.B1(n_1363),
.B2(n_1366),
.Y(n_1406)
);

OA21x2_ASAP7_75t_L g1407 ( 
.A1(n_1357),
.A2(n_1360),
.B(n_1356),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_1377),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1379),
.B(n_1381),
.Y(n_1409)
);

AOI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1338),
.A2(n_1370),
.B(n_1300),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1293),
.Y(n_1411)
);

OAI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1388),
.A2(n_1393),
.B(n_1389),
.Y(n_1412)
);

BUFx6f_ASAP7_75t_L g1413 ( 
.A(n_1342),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1365),
.A2(n_1356),
.B(n_1362),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1361),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1346),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1335),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1368),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1365),
.A2(n_1362),
.B(n_1351),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1381),
.B(n_1385),
.Y(n_1420)
);

INVxp67_ASAP7_75t_L g1421 ( 
.A(n_1337),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1354),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1316),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1333),
.A2(n_1327),
.B(n_1347),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1333),
.A2(n_1327),
.B(n_1296),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1358),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1296),
.B(n_1292),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1285),
.B(n_1303),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1289),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1336),
.A2(n_1340),
.B(n_1285),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1314),
.B(n_1385),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1386),
.B(n_1396),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1311),
.B(n_1299),
.Y(n_1433)
);

INVx2_ASAP7_75t_SL g1434 ( 
.A(n_1287),
.Y(n_1434)
);

OAI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1277),
.A2(n_1376),
.B1(n_1318),
.B2(n_1384),
.Y(n_1435)
);

AOI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1388),
.A2(n_1384),
.B1(n_1380),
.B2(n_1298),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1325),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1386),
.B(n_1396),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1353),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1353),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1320),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1320),
.Y(n_1442)
);

BUFx4f_ASAP7_75t_SL g1443 ( 
.A(n_1286),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1298),
.B(n_1372),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1302),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1348),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1290),
.B(n_1279),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1348),
.Y(n_1448)
);

BUFx6f_ASAP7_75t_L g1449 ( 
.A(n_1342),
.Y(n_1449)
);

INVxp33_ASAP7_75t_L g1450 ( 
.A(n_1308),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1342),
.Y(n_1451)
);

INVx3_ASAP7_75t_L g1452 ( 
.A(n_1343),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1323),
.A2(n_1372),
.B(n_1297),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1380),
.B(n_1310),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1334),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1334),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1367),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1367),
.Y(n_1458)
);

OA21x2_ASAP7_75t_L g1459 ( 
.A1(n_1306),
.A2(n_1319),
.B(n_1309),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1391),
.B(n_1294),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_1310),
.B(n_1326),
.Y(n_1461)
);

BUFx4f_ASAP7_75t_SL g1462 ( 
.A(n_1378),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1364),
.B(n_1332),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1344),
.Y(n_1464)
);

A2O1A1Ixp33_ASAP7_75t_L g1465 ( 
.A1(n_1305),
.A2(n_1390),
.B(n_1394),
.C(n_1382),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1307),
.B(n_1395),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1345),
.B(n_1305),
.Y(n_1467)
);

INVxp67_ASAP7_75t_L g1468 ( 
.A(n_1280),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1307),
.B(n_1281),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1297),
.Y(n_1470)
);

NAND4xp25_ASAP7_75t_L g1471 ( 
.A(n_1331),
.B(n_1278),
.C(n_1328),
.D(n_1324),
.Y(n_1471)
);

AO21x2_ASAP7_75t_L g1472 ( 
.A1(n_1339),
.A2(n_1390),
.B(n_1295),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1437),
.B(n_1324),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1412),
.A2(n_1307),
.B1(n_1322),
.B2(n_1374),
.Y(n_1474)
);

AOI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1436),
.A2(n_1283),
.B1(n_1330),
.B2(n_1291),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1463),
.B(n_1374),
.Y(n_1476)
);

AOI221xp5_ASAP7_75t_L g1477 ( 
.A1(n_1435),
.A2(n_1278),
.B1(n_1328),
.B2(n_1315),
.C(n_1295),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1416),
.B(n_1313),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_SL g1479 ( 
.A1(n_1436),
.A2(n_1472),
.B(n_1459),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1411),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1447),
.A2(n_1428),
.B1(n_1444),
.B2(n_1433),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1461),
.B(n_1339),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1399),
.B(n_1313),
.Y(n_1483)
);

AND2x2_ASAP7_75t_SL g1484 ( 
.A(n_1401),
.B(n_1276),
.Y(n_1484)
);

O2A1O1Ixp33_ASAP7_75t_SL g1485 ( 
.A1(n_1428),
.A2(n_1329),
.B(n_1315),
.C(n_1392),
.Y(n_1485)
);

O2A1O1Ixp33_ASAP7_75t_SL g1486 ( 
.A1(n_1465),
.A2(n_1282),
.B(n_1387),
.C(n_1304),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1444),
.A2(n_1317),
.B1(n_1304),
.B2(n_1375),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1399),
.B(n_1446),
.Y(n_1488)
);

OAI211xp5_ASAP7_75t_L g1489 ( 
.A1(n_1410),
.A2(n_1375),
.B(n_1301),
.C(n_1312),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1429),
.Y(n_1490)
);

O2A1O1Ixp33_ASAP7_75t_SL g1491 ( 
.A1(n_1431),
.A2(n_1301),
.B(n_1454),
.C(n_1464),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1446),
.B(n_1448),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1397),
.B(n_1459),
.Y(n_1493)
);

O2A1O1Ixp5_ASAP7_75t_L g1494 ( 
.A1(n_1410),
.A2(n_1439),
.B(n_1440),
.C(n_1454),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1459),
.B(n_1460),
.Y(n_1495)
);

AO21x2_ASAP7_75t_L g1496 ( 
.A1(n_1414),
.A2(n_1419),
.B(n_1404),
.Y(n_1496)
);

OAI211xp5_ASAP7_75t_L g1497 ( 
.A1(n_1401),
.A2(n_1438),
.B(n_1420),
.C(n_1409),
.Y(n_1497)
);

AOI221xp5_ASAP7_75t_L g1498 ( 
.A1(n_1409),
.A2(n_1432),
.B1(n_1438),
.B2(n_1420),
.C(n_1441),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_1431),
.B(n_1432),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1459),
.B(n_1460),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1464),
.A2(n_1442),
.B1(n_1441),
.B2(n_1468),
.Y(n_1501)
);

AOI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1464),
.A2(n_1442),
.B1(n_1418),
.B2(n_1469),
.Y(n_1502)
);

NOR2x1_ASAP7_75t_R g1503 ( 
.A(n_1408),
.B(n_1423),
.Y(n_1503)
);

AO32x2_ASAP7_75t_L g1504 ( 
.A1(n_1434),
.A2(n_1445),
.A3(n_1406),
.B1(n_1458),
.B2(n_1457),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1400),
.B(n_1403),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1403),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1448),
.B(n_1457),
.Y(n_1507)
);

OAI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1453),
.A2(n_1425),
.B(n_1430),
.Y(n_1508)
);

OA21x2_ASAP7_75t_L g1509 ( 
.A1(n_1414),
.A2(n_1424),
.B(n_1419),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_SL g1510 ( 
.A1(n_1434),
.A2(n_1445),
.B(n_1470),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1426),
.B(n_1452),
.Y(n_1511)
);

AO32x2_ASAP7_75t_L g1512 ( 
.A1(n_1406),
.A2(n_1407),
.A3(n_1456),
.B1(n_1455),
.B2(n_1415),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1400),
.B(n_1405),
.Y(n_1513)
);

AO22x2_ASAP7_75t_L g1514 ( 
.A1(n_1455),
.A2(n_1456),
.B1(n_1422),
.B2(n_1415),
.Y(n_1514)
);

OR2x6_ASAP7_75t_L g1515 ( 
.A(n_1453),
.B(n_1467),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1398),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1413),
.B(n_1449),
.Y(n_1517)
);

A2O1A1Ixp33_ASAP7_75t_L g1518 ( 
.A1(n_1427),
.A2(n_1424),
.B(n_1452),
.C(n_1413),
.Y(n_1518)
);

AND2x6_ASAP7_75t_L g1519 ( 
.A(n_1413),
.B(n_1449),
.Y(n_1519)
);

INVxp67_ASAP7_75t_L g1520 ( 
.A(n_1421),
.Y(n_1520)
);

AND2x4_ASAP7_75t_L g1521 ( 
.A(n_1513),
.B(n_1506),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1493),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1495),
.B(n_1407),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1516),
.Y(n_1524)
);

INVxp67_ASAP7_75t_L g1525 ( 
.A(n_1500),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1497),
.A2(n_1449),
.B1(n_1451),
.B2(n_1413),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1509),
.B(n_1404),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1509),
.B(n_1404),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1481),
.A2(n_1449),
.B1(n_1413),
.B2(n_1451),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1501),
.B(n_1450),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1500),
.B(n_1407),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_SL g1532 ( 
.A(n_1484),
.B(n_1449),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1490),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_1519),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1514),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1513),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1496),
.B(n_1405),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1496),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1518),
.B(n_1508),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1512),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1512),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1514),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1512),
.B(n_1518),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1492),
.B(n_1417),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1504),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1504),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1498),
.A2(n_1451),
.B1(n_1452),
.B2(n_1426),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1515),
.B(n_1402),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1514),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1534),
.Y(n_1550)
);

INVx5_ASAP7_75t_L g1551 ( 
.A(n_1527),
.Y(n_1551)
);

OAI33xp33_ASAP7_75t_L g1552 ( 
.A1(n_1549),
.A2(n_1546),
.A3(n_1541),
.B1(n_1540),
.B2(n_1526),
.B3(n_1547),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1529),
.A2(n_1474),
.B1(n_1487),
.B2(n_1484),
.Y(n_1553)
);

NOR2x1_ASAP7_75t_L g1554 ( 
.A(n_1534),
.B(n_1479),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1525),
.B(n_1511),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1525),
.B(n_1507),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1522),
.B(n_1507),
.Y(n_1557)
);

BUFx2_ASAP7_75t_SL g1558 ( 
.A(n_1534),
.Y(n_1558)
);

INVx1_ASAP7_75t_SL g1559 ( 
.A(n_1521),
.Y(n_1559)
);

NAND3xp33_ASAP7_75t_L g1560 ( 
.A(n_1539),
.B(n_1494),
.C(n_1502),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1522),
.B(n_1488),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1524),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1524),
.Y(n_1563)
);

AOI322xp5_ASAP7_75t_L g1564 ( 
.A1(n_1532),
.A2(n_1499),
.A3(n_1487),
.B1(n_1474),
.B2(n_1475),
.C1(n_1488),
.C2(n_1482),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1536),
.B(n_1505),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1531),
.B(n_1480),
.Y(n_1566)
);

OR2x6_ASAP7_75t_L g1567 ( 
.A(n_1539),
.B(n_1479),
.Y(n_1567)
);

OAI33xp33_ASAP7_75t_L g1568 ( 
.A1(n_1549),
.A2(n_1546),
.A3(n_1540),
.B1(n_1541),
.B2(n_1526),
.B3(n_1547),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1524),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1536),
.B(n_1505),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1531),
.B(n_1523),
.Y(n_1571)
);

AO21x2_ASAP7_75t_L g1572 ( 
.A1(n_1538),
.A2(n_1528),
.B(n_1527),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1533),
.Y(n_1573)
);

AND2x4_ASAP7_75t_SL g1574 ( 
.A(n_1529),
.B(n_1476),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1535),
.Y(n_1575)
);

AO21x2_ASAP7_75t_L g1576 ( 
.A1(n_1538),
.A2(n_1510),
.B(n_1489),
.Y(n_1576)
);

AOI211xp5_ASAP7_75t_L g1577 ( 
.A1(n_1526),
.A2(n_1482),
.B(n_1499),
.C(n_1491),
.Y(n_1577)
);

BUFx3_ASAP7_75t_L g1578 ( 
.A(n_1544),
.Y(n_1578)
);

OA211x2_ASAP7_75t_L g1579 ( 
.A1(n_1532),
.A2(n_1477),
.B(n_1520),
.C(n_1517),
.Y(n_1579)
);

NAND2x1_ASAP7_75t_L g1580 ( 
.A(n_1543),
.B(n_1519),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1566),
.B(n_1549),
.Y(n_1581)
);

INVx1_ASAP7_75t_SL g1582 ( 
.A(n_1574),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1575),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1551),
.B(n_1543),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1551),
.B(n_1543),
.Y(n_1585)
);

INVx1_ASAP7_75t_SL g1586 ( 
.A(n_1574),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1563),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1560),
.B(n_1478),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1571),
.B(n_1535),
.Y(n_1589)
);

INVx4_ASAP7_75t_L g1590 ( 
.A(n_1550),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1551),
.B(n_1543),
.Y(n_1591)
);

INVx2_ASAP7_75t_SL g1592 ( 
.A(n_1551),
.Y(n_1592)
);

INVx1_ASAP7_75t_SL g1593 ( 
.A(n_1558),
.Y(n_1593)
);

INVx3_ASAP7_75t_L g1594 ( 
.A(n_1551),
.Y(n_1594)
);

INVx3_ASAP7_75t_L g1595 ( 
.A(n_1551),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1571),
.B(n_1542),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1563),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1567),
.B(n_1545),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1569),
.Y(n_1599)
);

NAND2x1p5_ASAP7_75t_L g1600 ( 
.A(n_1554),
.B(n_1539),
.Y(n_1600)
);

AND2x4_ASAP7_75t_L g1601 ( 
.A(n_1554),
.B(n_1537),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1556),
.B(n_1542),
.Y(n_1602)
);

AND2x4_ASAP7_75t_SL g1603 ( 
.A(n_1550),
.B(n_1548),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1579),
.A2(n_1553),
.B1(n_1547),
.B2(n_1532),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1556),
.B(n_1483),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1562),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1569),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1567),
.B(n_1545),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1558),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1567),
.B(n_1545),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1573),
.Y(n_1611)
);

AND2x4_ASAP7_75t_SL g1612 ( 
.A(n_1550),
.B(n_1548),
.Y(n_1612)
);

INVx1_ASAP7_75t_SL g1613 ( 
.A(n_1557),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1573),
.Y(n_1614)
);

NAND3xp33_ASAP7_75t_L g1615 ( 
.A(n_1564),
.B(n_1539),
.C(n_1530),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1567),
.B(n_1545),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1572),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1567),
.B(n_1580),
.Y(n_1618)
);

INVx4_ASAP7_75t_L g1619 ( 
.A(n_1590),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1583),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1583),
.Y(n_1621)
);

INVx4_ASAP7_75t_L g1622 ( 
.A(n_1590),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1587),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1618),
.B(n_1565),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1587),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1606),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1597),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1606),
.Y(n_1628)
);

NAND2x1p5_ASAP7_75t_L g1629 ( 
.A(n_1593),
.B(n_1609),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1597),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1599),
.Y(n_1631)
);

AOI211xp5_ASAP7_75t_L g1632 ( 
.A1(n_1615),
.A2(n_1577),
.B(n_1491),
.C(n_1530),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1588),
.B(n_1443),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1618),
.B(n_1565),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1588),
.B(n_1578),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1602),
.B(n_1561),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1607),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1618),
.B(n_1570),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1606),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1602),
.B(n_1561),
.Y(n_1640)
);

O2A1O1Ixp33_ASAP7_75t_L g1641 ( 
.A1(n_1615),
.A2(n_1568),
.B(n_1552),
.C(n_1577),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1589),
.B(n_1596),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1611),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1614),
.Y(n_1644)
);

NOR5xp2_ASAP7_75t_L g1645 ( 
.A(n_1600),
.B(n_1546),
.C(n_1541),
.D(n_1540),
.E(n_1579),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1603),
.B(n_1570),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1605),
.B(n_1578),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1605),
.B(n_1555),
.Y(n_1648)
);

INVx1_ASAP7_75t_SL g1649 ( 
.A(n_1582),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1614),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1613),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1603),
.B(n_1612),
.Y(n_1652)
);

NOR2x1_ASAP7_75t_L g1653 ( 
.A(n_1590),
.B(n_1576),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1612),
.B(n_1559),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1612),
.B(n_1584),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1613),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1655),
.B(n_1592),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1655),
.B(n_1600),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1623),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1649),
.B(n_1582),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1652),
.B(n_1600),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1652),
.B(n_1600),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1642),
.B(n_1589),
.Y(n_1663)
);

NAND3xp33_ASAP7_75t_L g1664 ( 
.A(n_1641),
.B(n_1604),
.C(n_1564),
.Y(n_1664)
);

OAI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1632),
.A2(n_1604),
.B1(n_1586),
.B2(n_1609),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1623),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1635),
.B(n_1586),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1642),
.B(n_1596),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1651),
.B(n_1581),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1651),
.B(n_1581),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1629),
.B(n_1584),
.Y(n_1671)
);

INVxp67_ASAP7_75t_L g1672 ( 
.A(n_1629),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_SL g1673 ( 
.A(n_1633),
.B(n_1593),
.Y(n_1673)
);

NAND2x1p5_ASAP7_75t_L g1674 ( 
.A(n_1653),
.B(n_1594),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1629),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1625),
.Y(n_1676)
);

OAI21xp5_ASAP7_75t_SL g1677 ( 
.A1(n_1656),
.A2(n_1585),
.B(n_1584),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1624),
.B(n_1585),
.Y(n_1678)
);

NAND2x1p5_ASAP7_75t_L g1679 ( 
.A(n_1619),
.B(n_1622),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1656),
.B(n_1598),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1624),
.B(n_1585),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1625),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1619),
.B(n_1592),
.Y(n_1683)
);

INVx1_ASAP7_75t_SL g1684 ( 
.A(n_1647),
.Y(n_1684)
);

AOI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1648),
.A2(n_1486),
.B(n_1485),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1620),
.B(n_1598),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1620),
.A2(n_1486),
.B(n_1485),
.Y(n_1687)
);

AND2x2_ASAP7_75t_SL g1688 ( 
.A(n_1645),
.B(n_1591),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1626),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1634),
.B(n_1591),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1636),
.B(n_1462),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1621),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_SL g1693 ( 
.A(n_1664),
.B(n_1594),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1664),
.B(n_1621),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1688),
.A2(n_1591),
.B1(n_1640),
.B2(n_1636),
.Y(n_1695)
);

OAI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1665),
.A2(n_1592),
.B(n_1594),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1684),
.B(n_1640),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1688),
.A2(n_1528),
.B1(n_1527),
.B2(n_1483),
.Y(n_1698)
);

INVxp67_ASAP7_75t_L g1699 ( 
.A(n_1660),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1667),
.B(n_1691),
.Y(n_1700)
);

NAND3xp33_ASAP7_75t_L g1701 ( 
.A(n_1688),
.B(n_1622),
.C(n_1619),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1672),
.B(n_1598),
.Y(n_1702)
);

AOI21xp33_ASAP7_75t_L g1703 ( 
.A1(n_1673),
.A2(n_1622),
.B(n_1595),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1685),
.B(n_1608),
.Y(n_1704)
);

AOI221xp5_ASAP7_75t_L g1705 ( 
.A1(n_1677),
.A2(n_1669),
.B1(n_1670),
.B2(n_1680),
.C(n_1692),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1659),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1687),
.A2(n_1503),
.B(n_1594),
.Y(n_1707)
);

INVx2_ASAP7_75t_SL g1708 ( 
.A(n_1671),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1659),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1658),
.B(n_1634),
.Y(n_1710)
);

AOI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1675),
.A2(n_1595),
.B(n_1594),
.Y(n_1711)
);

AOI21xp33_ASAP7_75t_L g1712 ( 
.A1(n_1675),
.A2(n_1595),
.B(n_1627),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1671),
.Y(n_1713)
);

OAI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1674),
.A2(n_1595),
.B(n_1601),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1666),
.Y(n_1715)
);

OAI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1674),
.A2(n_1668),
.B1(n_1663),
.B2(n_1679),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1658),
.B(n_1638),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1678),
.B(n_1608),
.Y(n_1718)
);

INVx2_ASAP7_75t_SL g1719 ( 
.A(n_1708),
.Y(n_1719)
);

OAI32xp33_ASAP7_75t_L g1720 ( 
.A1(n_1695),
.A2(n_1674),
.A3(n_1679),
.B1(n_1668),
.B2(n_1663),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1699),
.B(n_1678),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1706),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1709),
.Y(n_1723)
);

A2O1A1Ixp33_ASAP7_75t_L g1724 ( 
.A1(n_1694),
.A2(n_1693),
.B(n_1696),
.C(n_1703),
.Y(n_1724)
);

OAI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1693),
.A2(n_1679),
.B(n_1662),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1697),
.B(n_1686),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1708),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1700),
.B(n_1661),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1713),
.B(n_1683),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1710),
.B(n_1661),
.Y(n_1730)
);

HB1xp67_ASAP7_75t_L g1731 ( 
.A(n_1715),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1717),
.Y(n_1732)
);

AOI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1698),
.A2(n_1662),
.B1(n_1657),
.B2(n_1681),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1705),
.B(n_1681),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1707),
.B(n_1657),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1701),
.Y(n_1736)
);

AOI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1698),
.A2(n_1657),
.B1(n_1690),
.B2(n_1683),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1731),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1731),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1727),
.Y(n_1740)
);

XNOR2xp5_ASAP7_75t_L g1741 ( 
.A(n_1732),
.B(n_1704),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1719),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1728),
.B(n_1716),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1729),
.B(n_1690),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1722),
.Y(n_1745)
);

XNOR2x2_ASAP7_75t_L g1746 ( 
.A(n_1725),
.B(n_1714),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_SL g1747 ( 
.A(n_1724),
.B(n_1716),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1723),
.Y(n_1748)
);

NOR4xp25_ASAP7_75t_L g1749 ( 
.A(n_1747),
.B(n_1736),
.C(n_1724),
.D(n_1734),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1738),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1743),
.B(n_1728),
.Y(n_1751)
);

NAND3xp33_ASAP7_75t_SL g1752 ( 
.A(n_1747),
.B(n_1737),
.C(n_1735),
.Y(n_1752)
);

INVxp67_ASAP7_75t_L g1753 ( 
.A(n_1743),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_L g1754 ( 
.A(n_1741),
.B(n_1735),
.Y(n_1754)
);

AOI221xp5_ASAP7_75t_L g1755 ( 
.A1(n_1739),
.A2(n_1720),
.B1(n_1721),
.B2(n_1729),
.C(n_1712),
.Y(n_1755)
);

NAND4xp25_ASAP7_75t_L g1756 ( 
.A(n_1742),
.B(n_1744),
.C(n_1740),
.D(n_1733),
.Y(n_1756)
);

NOR2xp33_ASAP7_75t_L g1757 ( 
.A(n_1746),
.B(n_1726),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_SL g1758 ( 
.A(n_1745),
.B(n_1730),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1748),
.Y(n_1759)
);

INVx1_ASAP7_75t_SL g1760 ( 
.A(n_1751),
.Y(n_1760)
);

O2A1O1Ixp33_ASAP7_75t_L g1761 ( 
.A1(n_1757),
.A2(n_1702),
.B(n_1711),
.C(n_1666),
.Y(n_1761)
);

OAI21xp5_ASAP7_75t_SL g1762 ( 
.A1(n_1752),
.A2(n_1657),
.B(n_1683),
.Y(n_1762)
);

AOI211xp5_ASAP7_75t_L g1763 ( 
.A1(n_1749),
.A2(n_1683),
.B(n_1718),
.C(n_1676),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1758),
.B(n_1638),
.Y(n_1764)
);

AOI221xp5_ASAP7_75t_L g1765 ( 
.A1(n_1753),
.A2(n_1682),
.B1(n_1676),
.B2(n_1689),
.C(n_1617),
.Y(n_1765)
);

A2O1A1Ixp33_ASAP7_75t_L g1766 ( 
.A1(n_1761),
.A2(n_1754),
.B(n_1755),
.C(n_1750),
.Y(n_1766)
);

AOI21xp5_ASAP7_75t_SL g1767 ( 
.A1(n_1764),
.A2(n_1759),
.B(n_1682),
.Y(n_1767)
);

OA211x2_ASAP7_75t_L g1768 ( 
.A1(n_1765),
.A2(n_1756),
.B(n_1466),
.C(n_1473),
.Y(n_1768)
);

OAI211xp5_ASAP7_75t_L g1769 ( 
.A1(n_1762),
.A2(n_1689),
.B(n_1595),
.C(n_1590),
.Y(n_1769)
);

AOI221x1_ASAP7_75t_SL g1770 ( 
.A1(n_1763),
.A2(n_1627),
.B1(n_1650),
.B2(n_1644),
.C(n_1643),
.Y(n_1770)
);

AOI211xp5_ASAP7_75t_L g1771 ( 
.A1(n_1760),
.A2(n_1601),
.B(n_1608),
.C(n_1610),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1767),
.Y(n_1772)
);

XNOR2x1_ASAP7_75t_L g1773 ( 
.A(n_1768),
.B(n_1601),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1770),
.B(n_1630),
.Y(n_1774)
);

OR3x2_ASAP7_75t_L g1775 ( 
.A(n_1766),
.B(n_1471),
.C(n_1630),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1771),
.B(n_1646),
.Y(n_1776)
);

NAND2x1p5_ASAP7_75t_L g1777 ( 
.A(n_1772),
.B(n_1769),
.Y(n_1777)
);

NAND3xp33_ASAP7_75t_SL g1778 ( 
.A(n_1774),
.B(n_1590),
.C(n_1654),
.Y(n_1778)
);

AOI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1776),
.A2(n_1601),
.B1(n_1616),
.B2(n_1610),
.Y(n_1779)
);

INVx3_ASAP7_75t_L g1780 ( 
.A(n_1777),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1780),
.Y(n_1781)
);

OAI22x1_ASAP7_75t_L g1782 ( 
.A1(n_1781),
.A2(n_1780),
.B1(n_1774),
.B2(n_1779),
.Y(n_1782)
);

OAI22x1_ASAP7_75t_L g1783 ( 
.A1(n_1781),
.A2(n_1775),
.B1(n_1778),
.B2(n_1773),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1783),
.Y(n_1784)
);

CKINVDCx20_ASAP7_75t_R g1785 ( 
.A(n_1782),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1784),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1785),
.A2(n_1628),
.B1(n_1626),
.B2(n_1639),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1786),
.Y(n_1788)
);

OAI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1788),
.A2(n_1787),
.B(n_1639),
.Y(n_1789)
);

HB1xp67_ASAP7_75t_L g1790 ( 
.A(n_1789),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1790),
.A2(n_1628),
.B1(n_1617),
.B2(n_1631),
.Y(n_1791)
);

AOI211xp5_ASAP7_75t_L g1792 ( 
.A1(n_1791),
.A2(n_1643),
.B(n_1637),
.C(n_1631),
.Y(n_1792)
);


endmodule