module fake_aes_8754_n_33 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_33);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_30;
wire n_13;
wire n_26;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx16_ASAP7_75t_R g10 ( .A(n_7), .Y(n_10) );
BUFx2_ASAP7_75t_L g11 ( .A(n_6), .Y(n_11) );
HB1xp67_ASAP7_75t_L g12 ( .A(n_2), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_5), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_5), .B(n_4), .Y(n_14) );
BUFx2_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_15), .B(n_11), .Y(n_16) );
NAND3xp33_ASAP7_75t_SL g17 ( .A(n_15), .B(n_0), .C(n_2), .Y(n_17) );
AND2x4_ASAP7_75t_L g18 ( .A(n_11), .B(n_0), .Y(n_18) );
OAI22x1_ASAP7_75t_L g19 ( .A1(n_12), .A2(n_3), .B1(n_4), .B2(n_8), .Y(n_19) );
NAND2xp5_ASAP7_75t_SL g20 ( .A(n_10), .B(n_3), .Y(n_20) );
NOR2xp33_ASAP7_75t_R g21 ( .A(n_16), .B(n_14), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_18), .Y(n_22) );
NAND3xp33_ASAP7_75t_L g23 ( .A(n_18), .B(n_13), .C(n_14), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_20), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_22), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_23), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g27 ( .A(n_21), .B(n_17), .Y(n_27) );
INVx3_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
AND3x1_ASAP7_75t_L g29 ( .A(n_27), .B(n_24), .C(n_17), .Y(n_29) );
INVx1_ASAP7_75t_SL g30 ( .A(n_28), .Y(n_30) );
OA22x2_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_19), .B1(n_26), .B2(n_28), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_31), .Y(n_32) );
AOI22xp33_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_25), .B1(n_29), .B2(n_9), .Y(n_33) );
endmodule