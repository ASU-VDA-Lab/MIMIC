module fake_jpeg_16961_n_359 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_359);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_359;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx6_ASAP7_75t_SL g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_9),
.B(n_7),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_SL g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_40),
.B(n_44),
.Y(n_114)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_22),
.Y(n_49)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_49),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_51),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_55),
.Y(n_79)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_59),
.Y(n_81)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_63),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_61),
.Y(n_124)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_67),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_68),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_70),
.Y(n_87)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_72),
.Y(n_96)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_38),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_39),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_76),
.B(n_77),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_39),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_39),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_83),
.B(n_90),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_43),
.A2(n_17),
.B1(n_25),
.B2(n_30),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_86),
.A2(n_112),
.B1(n_117),
.B2(n_3),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_41),
.A2(n_25),
.B1(n_34),
.B2(n_27),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_88),
.A2(n_92),
.B1(n_95),
.B2(n_109),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_30),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_30),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_91),
.B(n_93),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_17),
.B1(n_21),
.B2(n_25),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_21),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_21),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_94),
.B(n_103),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_42),
.A2(n_17),
.B1(n_34),
.B2(n_24),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_97),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_23),
.Y(n_98)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_23),
.Y(n_100)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_24),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_62),
.A2(n_38),
.B1(n_37),
.B2(n_35),
.Y(n_104)
);

OAI32xp33_ASAP7_75t_L g170 ( 
.A1(n_104),
.A2(n_84),
.A3(n_79),
.B1(n_87),
.B2(n_99),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_37),
.Y(n_105)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_105),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_35),
.C(n_33),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_108),
.B(n_109),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_66),
.A2(n_33),
.B1(n_32),
.B2(n_15),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_57),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_58),
.B(n_32),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_113),
.B(n_9),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_49),
.A2(n_15),
.B1(n_12),
.B2(n_10),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_60),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_9),
.B1(n_69),
.B2(n_50),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_54),
.B(n_10),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_121),
.B(n_123),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_73),
.B(n_0),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_68),
.B(n_2),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_125),
.B(n_4),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_126),
.A2(n_133),
.B1(n_168),
.B2(n_158),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_51),
.Y(n_127)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_127),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_119),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_130),
.B(n_145),
.Y(n_187)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_131),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_132),
.B(n_172),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_82),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_135),
.A2(n_152),
.B1(n_161),
.B2(n_170),
.Y(n_179)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_7),
.C(n_8),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_137),
.A2(n_124),
.B(n_101),
.C(n_118),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_77),
.A2(n_45),
.B(n_47),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_139),
.A2(n_173),
.B(n_174),
.Y(n_203)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_141),
.Y(n_193)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_143),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_144),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_107),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_146),
.B(n_156),
.Y(n_215)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_114),
.B(n_8),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_148),
.B(n_154),
.Y(n_200)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_150),
.Y(n_208)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_151),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_85),
.B(n_9),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_155),
.B(n_163),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_78),
.Y(n_157)
);

INVxp67_ASAP7_75t_SL g185 ( 
.A(n_157),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_158),
.B(n_160),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_120),
.A2(n_104),
.B1(n_125),
.B2(n_95),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_75),
.A2(n_106),
.B1(n_102),
.B2(n_122),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_108),
.B(n_113),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_74),
.Y(n_164)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_111),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_165),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_111),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_166),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_102),
.A2(n_122),
.B1(n_81),
.B2(n_104),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_167),
.A2(n_152),
.B1(n_159),
.B2(n_141),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_92),
.A2(n_104),
.B1(n_93),
.B2(n_94),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_83),
.B(n_90),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_171),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_80),
.B(n_74),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_80),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_75),
.A2(n_106),
.B1(n_124),
.B2(n_101),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_124),
.A2(n_36),
.B1(n_19),
.B2(n_43),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g227 ( 
.A(n_176),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_118),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_178),
.B(n_181),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_155),
.C(n_169),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_131),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_183),
.B(n_184),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_138),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_138),
.B(n_136),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_189),
.B(n_206),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_190),
.A2(n_176),
.B1(n_186),
.B2(n_194),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_153),
.B(n_129),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_197),
.B(n_199),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_198),
.A2(n_179),
.B1(n_209),
.B2(n_206),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_136),
.B(n_160),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_139),
.B(n_142),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_201),
.B(n_207),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_143),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_147),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_170),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_142),
.B(n_171),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_128),
.B(n_134),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_211),
.A2(n_213),
.B(n_215),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_146),
.A2(n_175),
.B1(n_162),
.B2(n_149),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_150),
.B(n_156),
.Y(n_214)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_214),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_151),
.B(n_164),
.Y(n_216)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_216),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_216),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_217),
.B(n_245),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_219),
.A2(n_224),
.B1(n_247),
.B2(n_246),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_220),
.Y(n_271)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_223),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_177),
.A2(n_157),
.B(n_144),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_247),
.Y(n_258)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_225),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_178),
.B(n_165),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_226),
.A2(n_228),
.B1(n_243),
.B2(n_251),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_177),
.A2(n_166),
.B(n_201),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_228),
.Y(n_270)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_192),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_232),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_230),
.A2(n_235),
.B1(n_238),
.B2(n_240),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_204),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_241),
.Y(n_252)
);

INVxp33_ASAP7_75t_L g232 ( 
.A(n_187),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_193),
.B(n_207),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_248),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_198),
.A2(n_209),
.B1(n_190),
.B2(n_210),
.Y(n_235)
);

BUFx24_ASAP7_75t_L g236 ( 
.A(n_185),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_236),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_209),
.A2(n_182),
.B1(n_184),
.B2(n_183),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_203),
.A2(n_182),
.B1(n_189),
.B2(n_181),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_200),
.B(n_213),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_195),
.B(n_212),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_244),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_203),
.A2(n_211),
.B1(n_180),
.B2(n_186),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_243),
.A2(n_246),
.B1(n_226),
.B2(n_217),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_202),
.B(n_192),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_180),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_211),
.A2(n_205),
.B(n_208),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_191),
.B(n_194),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_188),
.B(n_187),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_251),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_188),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_229),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_253),
.B(n_269),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_222),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_222),
.Y(n_282)
);

A2O1A1Ixp33_ASAP7_75t_L g256 ( 
.A1(n_239),
.A2(n_227),
.B(n_241),
.C(n_230),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_256),
.B(n_264),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_259),
.A2(n_276),
.B(n_226),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_261),
.A2(n_258),
.B1(n_279),
.B2(n_264),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_218),
.B(n_225),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_218),
.B(n_234),
.Y(n_266)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_266),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_221),
.B(n_237),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_267),
.B(n_266),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_221),
.Y(n_268)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_268),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_231),
.B(n_220),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_238),
.B(n_250),
.Y(n_272)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_220),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_223),
.B(n_242),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_277),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_237),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_219),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_240),
.B(n_235),
.Y(n_280)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_282),
.B(n_285),
.C(n_275),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_284),
.A2(n_290),
.B1(n_292),
.B2(n_295),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_254),
.B(n_239),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_286),
.B(n_294),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_270),
.A2(n_236),
.B1(n_280),
.B2(n_261),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_270),
.A2(n_236),
.B1(n_279),
.B2(n_276),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_265),
.B(n_255),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_293),
.Y(n_305)
);

NOR3xp33_ASAP7_75t_L g294 ( 
.A(n_252),
.B(n_236),
.C(n_257),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_275),
.A2(n_271),
.B1(n_262),
.B2(n_253),
.Y(n_296)
);

INVx13_ASAP7_75t_L g309 ( 
.A(n_296),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_267),
.B(n_252),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_300),
.Y(n_312)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_263),
.Y(n_299)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_299),
.Y(n_306)
);

NAND3xp33_ASAP7_75t_L g301 ( 
.A(n_257),
.B(n_255),
.C(n_256),
.Y(n_301)
);

OA21x2_ASAP7_75t_SL g315 ( 
.A1(n_301),
.A2(n_298),
.B(n_303),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_268),
.A2(n_272),
.B1(n_274),
.B2(n_262),
.Y(n_302)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_260),
.B(n_265),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_303),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_274),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_317),
.C(n_319),
.Y(n_323)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_299),
.Y(n_308)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_308),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_258),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_311),
.B(n_314),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_284),
.B(n_260),
.Y(n_314)
);

HAxp5_ASAP7_75t_SL g327 ( 
.A(n_315),
.B(n_287),
.CON(n_327),
.SN(n_327)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_281),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_318),
.A2(n_283),
.B(n_288),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_289),
.B(n_271),
.C(n_273),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_297),
.Y(n_320)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_320),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_300),
.Y(n_321)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_321),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_305),
.B(n_291),
.Y(n_324)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_324),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_304),
.B(n_302),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_326),
.B(n_334),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_327),
.B(n_330),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_318),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_328),
.B(n_329),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_312),
.B(n_283),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_308),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_331),
.A2(n_332),
.B1(n_313),
.B2(n_320),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_316),
.A2(n_297),
.B1(n_288),
.B2(n_289),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_307),
.A2(n_292),
.B(n_290),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_323),
.B(n_317),
.C(n_319),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_338),
.B(n_339),
.C(n_340),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_323),
.B(n_314),
.Y(n_340)
);

BUFx24_ASAP7_75t_SL g342 ( 
.A(n_333),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_342),
.B(n_305),
.Y(n_350)
);

AOI322xp5_ASAP7_75t_L g343 ( 
.A1(n_334),
.A2(n_309),
.A3(n_315),
.B1(n_287),
.B2(n_313),
.C1(n_306),
.C2(n_311),
.Y(n_343)
);

AOI21xp33_ASAP7_75t_L g349 ( 
.A1(n_343),
.A2(n_337),
.B(n_335),
.Y(n_349)
);

AOI31xp67_ASAP7_75t_SL g345 ( 
.A1(n_341),
.A2(n_330),
.A3(n_310),
.B(n_306),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_345),
.B(n_347),
.Y(n_353)
);

NAND3xp33_ASAP7_75t_L g347 ( 
.A(n_344),
.B(n_310),
.C(n_329),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_338),
.B(n_333),
.C(n_326),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_348),
.A2(n_349),
.B1(n_350),
.B2(n_321),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_346),
.A2(n_309),
.B1(n_331),
.B2(n_325),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_351),
.A2(n_322),
.B1(n_325),
.B2(n_332),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_352),
.B(n_340),
.C(n_336),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_354),
.B(n_355),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_356),
.B(n_353),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_357),
.A2(n_351),
.B1(n_355),
.B2(n_322),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_358),
.B(n_336),
.Y(n_359)
);


endmodule