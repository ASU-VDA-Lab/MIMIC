module fake_jpeg_29046_n_305 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_305);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_305;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_11),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_34),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_36),
.Y(n_48)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_23),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_19),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_19),
.B1(n_31),
.B2(n_27),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_45),
.A2(n_54),
.B1(n_56),
.B2(n_36),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_52),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_19),
.B1(n_31),
.B2(n_27),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_30),
.B1(n_41),
.B2(n_27),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_30),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_29),
.B1(n_16),
.B2(n_22),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_21),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_31),
.B1(n_27),
.B2(n_29),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_30),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_41),
.C(n_36),
.Y(n_90)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_54),
.A2(n_22),
.B1(n_16),
.B2(n_28),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_62),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_77),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_60),
.A2(n_22),
.B1(n_16),
.B2(n_28),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_66),
.A2(n_99),
.B(n_36),
.Y(n_123)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_41),
.B(n_40),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_68),
.A2(n_36),
.B(n_37),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_57),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_69),
.B(n_71),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_48),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_78),
.A2(n_39),
.B1(n_38),
.B2(n_37),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_20),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_85),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_51),
.A2(n_41),
.B1(n_28),
.B2(n_32),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_80),
.A2(n_84),
.B1(n_36),
.B2(n_37),
.Y(n_113)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_83),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_53),
.B(n_20),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_87),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_56),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_89),
.Y(n_119)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_98),
.C(n_36),
.Y(n_106)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_95),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_49),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_93),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_49),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_94),
.B(n_100),
.Y(n_120)
);

INVx4_ASAP7_75t_SL g95 ( 
.A(n_59),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_97),
.Y(n_109)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_46),
.B(n_42),
.C(n_26),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_54),
.A2(n_32),
.B1(n_18),
.B2(n_42),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_60),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_103),
.A2(n_90),
.B(n_76),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_124),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_78),
.B1(n_77),
.B2(n_81),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_69),
.B(n_33),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_24),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_87),
.A2(n_42),
.B1(n_37),
.B2(n_38),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_122),
.A2(n_126),
.B1(n_128),
.B2(n_38),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_123),
.A2(n_93),
.B(n_96),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_63),
.B(n_21),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_91),
.A2(n_42),
.B1(n_32),
.B2(n_38),
.Y(n_128)
);

INVxp33_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_155),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_68),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_133),
.B(n_136),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_137),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_114),
.B(n_63),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_138),
.A2(n_146),
.B1(n_156),
.B2(n_144),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_118),
.Y(n_139)
);

NAND2xp33_ASAP7_75t_SL g169 ( 
.A(n_139),
.B(n_143),
.Y(n_169)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

AO22x1_ASAP7_75t_SL g142 ( 
.A1(n_113),
.A2(n_63),
.B1(n_75),
.B2(n_83),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_142),
.B(n_145),
.Y(n_184)
);

AOI22x1_ASAP7_75t_SL g143 ( 
.A1(n_107),
.A2(n_21),
.B1(n_98),
.B2(n_92),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_144),
.Y(n_190)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_105),
.A2(n_75),
.B1(n_61),
.B2(n_73),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_111),
.B1(n_127),
.B2(n_129),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_120),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_148),
.B(n_149),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_120),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_102),
.B(n_67),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_151),
.B(n_153),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_86),
.B1(n_95),
.B2(n_88),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_152),
.A2(n_158),
.B1(n_159),
.B2(n_127),
.Y(n_167)
);

NAND2x1_ASAP7_75t_L g153 ( 
.A(n_103),
.B(n_70),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_119),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_154),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_121),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_128),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_147),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_106),
.B(n_89),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_160),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_126),
.A2(n_64),
.B1(n_74),
.B2(n_97),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_122),
.A2(n_39),
.B1(n_38),
.B2(n_82),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_124),
.A2(n_33),
.B(n_25),
.C(n_24),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_161),
.A2(n_167),
.B1(n_146),
.B2(n_139),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_162),
.A2(n_158),
.B1(n_145),
.B2(n_150),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_143),
.A2(n_104),
.B1(n_123),
.B2(n_129),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_163),
.A2(n_18),
.B1(n_35),
.B2(n_8),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_115),
.C(n_117),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_174),
.C(n_177),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_135),
.A2(n_115),
.B1(n_117),
.B2(n_111),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_171),
.A2(n_179),
.B1(n_187),
.B2(n_159),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_108),
.C(n_110),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_132),
.B(n_108),
.C(n_110),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_133),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_154),
.A2(n_112),
.B1(n_116),
.B2(n_18),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_136),
.B(n_133),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_186),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_134),
.B(n_25),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_6),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_116),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_151),
.A2(n_116),
.B1(n_112),
.B2(n_39),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_151),
.B(n_112),
.C(n_39),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_191),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_152),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_18),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_153),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_210),
.C(n_211),
.Y(n_227)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_178),
.Y(n_195)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_195),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_196),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_197),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_229)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_190),
.Y(n_198)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_173),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_199),
.B(n_206),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_200),
.A2(n_201),
.B1(n_214),
.B2(n_183),
.Y(n_234)
);

OAI32xp33_ASAP7_75t_L g202 ( 
.A1(n_184),
.A2(n_153),
.A3(n_18),
.B1(n_38),
.B2(n_39),
.Y(n_202)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_186),
.A2(n_39),
.B1(n_9),
.B2(n_10),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_167),
.A2(n_35),
.B1(n_6),
.B2(n_10),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_172),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_209),
.B(n_212),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_35),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_35),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_175),
.B(n_15),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_168),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_174),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_162),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_166),
.A2(n_179),
.B(n_164),
.Y(n_215)
);

AO21x1_ASAP7_75t_L g235 ( 
.A1(n_215),
.A2(n_218),
.B(n_169),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_187),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_216),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_165),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_217),
.Y(n_236)
);

AO21x1_ASAP7_75t_L g218 ( 
.A1(n_166),
.A2(n_35),
.B(n_14),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_180),
.Y(n_219)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_168),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_194),
.Y(n_240)
);

XNOR2x1_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_177),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_239),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_183),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_230),
.Y(n_248)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_202),
.Y(n_230)
);

BUFx4f_ASAP7_75t_SL g232 ( 
.A(n_218),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_232),
.Y(n_253)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_203),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_238),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_234),
.A2(n_12),
.B1(n_11),
.B2(n_2),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_14),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_170),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_219),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_233),
.A2(n_207),
.B1(n_197),
.B2(n_192),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_241),
.A2(n_242),
.B1(n_231),
.B2(n_234),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_229),
.A2(n_207),
.B1(n_192),
.B2(n_191),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_208),
.C(n_213),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_250),
.C(n_251),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_236),
.B(n_208),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_247),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_188),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_171),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_254),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_215),
.C(n_164),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_211),
.C(n_210),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_252),
.B(n_255),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_238),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_0),
.C(n_1),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_220),
.C(n_226),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_271),
.Y(n_276)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_260),
.Y(n_275)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_248),
.Y(n_261)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_253),
.A2(n_224),
.B1(n_230),
.B2(n_231),
.Y(n_262)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_262),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_267),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_265),
.B(n_257),
.Y(n_272)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_244),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_220),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_235),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_224),
.C(n_225),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_245),
.C(n_251),
.Y(n_273)
);

AO21x1_ASAP7_75t_L g271 ( 
.A1(n_250),
.A2(n_232),
.B(n_228),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_274),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_267),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_256),
.C(n_229),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_280),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_232),
.C(n_1),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_288),
.C(n_287),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_280),
.A2(n_271),
.B(n_263),
.Y(n_284)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_284),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_276),
.A2(n_268),
.B(n_269),
.Y(n_285)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_285),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_277),
.B(n_265),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_286),
.A2(n_289),
.B(n_281),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_264),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_279),
.A2(n_270),
.B(n_262),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_275),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_291),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_292),
.B(n_276),
.C(n_286),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_297),
.Y(n_298)
);

NOR2xp67_ASAP7_75t_SL g297 ( 
.A(n_294),
.B(n_0),
.Y(n_297)
);

AOI21xp33_ASAP7_75t_L g299 ( 
.A1(n_296),
.A2(n_293),
.B(n_290),
.Y(n_299)
);

A2O1A1O1Ixp25_ASAP7_75t_L g300 ( 
.A1(n_299),
.A2(n_1),
.B(n_2),
.C(n_3),
.D(n_4),
.Y(n_300)
);

AOI321xp33_ASAP7_75t_L g301 ( 
.A1(n_300),
.A2(n_298),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C(n_2),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_2),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_302),
.A2(n_3),
.B(n_4),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_303),
.B(n_3),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_4),
.Y(n_305)
);


endmodule