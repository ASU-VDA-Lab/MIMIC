module fake_jpeg_19097_n_310 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_310);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_310;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_26),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_18),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_0),
.Y(n_27)
);

AOI21xp33_ASAP7_75t_L g35 ( 
.A1(n_27),
.A2(n_20),
.B(n_12),
.Y(n_35)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_35),
.B(n_27),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_32),
.A2(n_13),
.B1(n_11),
.B2(n_20),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_25),
.C(n_26),
.Y(n_60)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_27),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_47),
.B(n_55),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_25),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_36),
.Y(n_64)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_50),
.Y(n_79)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_52),
.Y(n_67)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_53),
.A2(n_39),
.B1(n_38),
.B2(n_28),
.Y(n_70)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_32),
.B1(n_26),
.B2(n_25),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_56),
.A2(n_37),
.B1(n_43),
.B2(n_32),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_57),
.Y(n_69)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_36),
.B1(n_28),
.B2(n_41),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_61),
.A2(n_74),
.B1(n_39),
.B2(n_58),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_66),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_37),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_30),
.C(n_24),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_78),
.C(n_30),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_38),
.B1(n_45),
.B2(n_54),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_72),
.A2(n_39),
.B1(n_28),
.B2(n_53),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_36),
.B1(n_28),
.B2(n_43),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_31),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_24),
.C(n_29),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_31),
.Y(n_117)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_77),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_62),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_84),
.B(n_86),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_64),
.B(n_41),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_88),
.A2(n_70),
.B1(n_72),
.B2(n_69),
.Y(n_111)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_41),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_93),
.B(n_95),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_66),
.A2(n_31),
.B(n_43),
.C(n_50),
.Y(n_94)
);

AO22x1_ASAP7_75t_L g120 ( 
.A1(n_94),
.A2(n_99),
.B1(n_31),
.B2(n_24),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_52),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_49),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_96),
.B(n_98),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_75),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_43),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_12),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_100),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_91),
.A2(n_76),
.B(n_65),
.Y(n_103)
);

HAxp5_ASAP7_75t_SL g150 ( 
.A(n_103),
.B(n_108),
.CON(n_150),
.SN(n_150)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_76),
.B(n_71),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_111),
.A2(n_119),
.B1(n_99),
.B2(n_84),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_86),
.A2(n_71),
.B(n_78),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_78),
.C(n_74),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_117),
.C(n_125),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_96),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_118),
.Y(n_127)
);

BUFx24_ASAP7_75t_SL g118 ( 
.A(n_100),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_89),
.A2(n_39),
.B1(n_80),
.B2(n_67),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_126),
.Y(n_128)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_85),
.A2(n_73),
.B(n_67),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_87),
.Y(n_124)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_68),
.C(n_75),
.Y(n_126)
);

NOR2x1_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_94),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_159),
.Y(n_164)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_93),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_137),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_134),
.B(n_135),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_102),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_110),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_138),
.B(n_149),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_105),
.A2(n_90),
.B1(n_98),
.B2(n_99),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_144),
.B1(n_80),
.B2(n_63),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_102),
.B(n_94),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_141),
.B(n_142),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_84),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_143),
.A2(n_120),
.B1(n_80),
.B2(n_13),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_105),
.A2(n_97),
.B1(n_88),
.B2(n_83),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_101),
.B(n_92),
.Y(n_145)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_145),
.Y(n_188)
);

XNOR2x2_ASAP7_75t_SL g147 ( 
.A(n_103),
.B(n_97),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_112),
.B(n_117),
.C(n_107),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_75),
.Y(n_148)
);

AO22x1_ASAP7_75t_L g177 ( 
.A1(n_148),
.A2(n_142),
.B1(n_137),
.B2(n_132),
.Y(n_177)
);

AND2x6_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_68),
.Y(n_149)
);

OAI22x1_ASAP7_75t_L g151 ( 
.A1(n_111),
.A2(n_63),
.B1(n_83),
.B2(n_69),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_152),
.B1(n_157),
.B2(n_31),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_119),
.Y(n_152)
);

OAI21xp33_ASAP7_75t_L g153 ( 
.A1(n_121),
.A2(n_31),
.B(n_83),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_153),
.A2(n_158),
.B(n_33),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_77),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_154),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_106),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_126),
.B(n_63),
.Y(n_157)
);

A2O1A1Ixp33_ASAP7_75t_SL g158 ( 
.A1(n_120),
.A2(n_122),
.B(n_106),
.C(n_108),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_115),
.B(n_63),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_161),
.B(n_168),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_163),
.A2(n_172),
.B1(n_189),
.B2(n_129),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_167),
.A2(n_171),
.B1(n_176),
.B2(n_180),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_31),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_169),
.B(n_33),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_51),
.C(n_57),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_173),
.C(n_185),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_139),
.A2(n_0),
.B1(n_13),
.B2(n_2),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_59),
.B1(n_46),
.B2(n_19),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_128),
.B(n_51),
.C(n_57),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_160),
.A2(n_46),
.B(n_57),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_177),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_22),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_136),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_178),
.A2(n_182),
.B(n_186),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_40),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_181),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_144),
.A2(n_156),
.B1(n_130),
.B2(n_160),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_128),
.B(n_40),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_30),
.C(n_29),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_158),
.A2(n_59),
.B1(n_14),
.B2(n_21),
.Y(n_189)
);

XNOR2x1_ASAP7_75t_SL g190 ( 
.A(n_164),
.B(n_150),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_190),
.B(n_171),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_184),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_191),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_187),
.A2(n_127),
.B1(n_146),
.B2(n_129),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_195),
.A2(n_208),
.B1(n_178),
.B2(n_172),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_148),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_207),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_138),
.Y(n_197)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_150),
.C(n_147),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_201),
.C(n_210),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_163),
.A2(n_131),
.B1(n_158),
.B2(n_134),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_200),
.A2(n_205),
.B1(n_176),
.B2(n_174),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_158),
.C(n_133),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_162),
.B(n_188),
.Y(n_203)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_209),
.Y(n_229)
);

AOI21xp33_ASAP7_75t_L g205 ( 
.A1(n_178),
.A2(n_158),
.B(n_22),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_33),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_162),
.B(n_22),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_30),
.C(n_29),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_164),
.B(n_29),
.C(n_24),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_212),
.C(n_189),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_177),
.C(n_180),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_33),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_213),
.B(n_182),
.C(n_167),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_191),
.B(n_175),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_214),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_217),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_220),
.C(n_224),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_186),
.C(n_165),
.Y(n_220)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_183),
.C(n_161),
.Y(n_224)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_175),
.C(n_17),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_230),
.C(n_232),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_17),
.C(n_16),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_192),
.B(n_15),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_233),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_202),
.B(n_22),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_206),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_198),
.B(n_15),
.C(n_17),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_207),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_201),
.B(n_17),
.C(n_15),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_210),
.C(n_193),
.Y(n_241)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

OAI321xp33_ASAP7_75t_L g239 ( 
.A1(n_228),
.A2(n_190),
.A3(n_213),
.B1(n_211),
.B2(n_208),
.C(n_193),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_239),
.A2(n_235),
.B1(n_230),
.B2(n_3),
.Y(n_261)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_223),
.A2(n_23),
.B(n_1),
.Y(n_242)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_17),
.C(n_15),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_248),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_17),
.C(n_15),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_229),
.A2(n_7),
.B(n_1),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_249),
.A2(n_251),
.B(n_9),
.Y(n_259)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_250),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_222),
.A2(n_7),
.B(n_1),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_219),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_218),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_243),
.B(n_218),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_260),
.Y(n_274)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_225),
.B1(n_226),
.B2(n_232),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_256),
.A2(n_262),
.B1(n_240),
.B2(n_23),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_227),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_259),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_241),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_261),
.A2(n_7),
.B1(n_2),
.B2(n_3),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_246),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_237),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_260),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_258),
.A2(n_248),
.B(n_245),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_267),
.A2(n_271),
.B(n_7),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_254),
.A2(n_244),
.B(n_249),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_268),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_264),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_279),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_263),
.A2(n_251),
.B(n_240),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_275),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_273),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_23),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_21),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_277),
.B(n_278),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_21),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_271),
.A2(n_265),
.B1(n_259),
.B2(n_21),
.Y(n_280)
);

NOR2xp67_ASAP7_75t_SL g294 ( 
.A(n_280),
.B(n_4),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_283),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_19),
.C(n_14),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_272),
.B(n_276),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_4),
.Y(n_298)
);

NOR2xp67_ASAP7_75t_SL g289 ( 
.A(n_270),
.B(n_19),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_289),
.A2(n_0),
.B(n_4),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_269),
.A2(n_19),
.B(n_14),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_290),
.A2(n_4),
.B(n_5),
.Y(n_295)
);

OA21x2_ASAP7_75t_SL g291 ( 
.A1(n_270),
.A2(n_4),
.B(n_5),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_5),
.C(n_6),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_293),
.C(n_294),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_0),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_295),
.A2(n_298),
.B(n_5),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_282),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_296),
.A2(n_285),
.B(n_280),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_286),
.C(n_288),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_300),
.A2(n_285),
.B(n_298),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_302),
.A2(n_303),
.B(n_297),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_304),
.B(n_305),
.Y(n_306)
);

AOI322xp5_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_6),
.A3(n_7),
.B1(n_9),
.B2(n_10),
.C1(n_301),
.C2(n_304),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_6),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_9),
.Y(n_309)
);

OAI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_309),
.A2(n_9),
.B1(n_10),
.B2(n_265),
.Y(n_310)
);


endmodule