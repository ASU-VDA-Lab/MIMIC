module real_aes_13887_n_3 (n_0, n_2, n_1, n_3);
input n_0;
input n_2;
input n_1;
output n_3;
wire n_4;
wire n_5;
wire n_7;
wire n_9;
wire n_6;
wire n_8;
INVx3_ASAP7_75t_L g8 ( .A(n_0), .Y(n_8) );
AOI22xp33_ASAP7_75t_L g3 ( .A1(n_1), .A2(n_2), .B1(n_4), .B2(n_9), .Y(n_3) );
INVx3_ASAP7_75t_L g4 ( .A(n_5), .Y(n_4) );
BUFx6f_ASAP7_75t_L g9 ( .A(n_5), .Y(n_9) );
INVx2_ASAP7_75t_L g5 ( .A(n_6), .Y(n_5) );
INVx2_ASAP7_75t_L g6 ( .A(n_7), .Y(n_6) );
INVx2_ASAP7_75t_L g7 ( .A(n_8), .Y(n_7) );
endmodule