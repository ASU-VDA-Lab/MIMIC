module fake_jpeg_3028_n_120 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_120);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_120;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_21),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_45),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_47),
.Y(n_58)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_49),
.Y(n_56)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

CKINVDCx12_ASAP7_75t_R g60 ( 
.A(n_50),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_49),
.A2(n_42),
.B1(n_40),
.B2(n_33),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_51),
.A2(n_38),
.B1(n_15),
.B2(n_16),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_33),
.B1(n_39),
.B2(n_34),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_59),
.B1(n_38),
.B2(n_14),
.Y(n_64)
);

AO22x1_ASAP7_75t_SL g55 ( 
.A1(n_47),
.A2(n_37),
.B1(n_36),
.B2(n_35),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_57),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_37),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_43),
.B1(n_39),
.B2(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_62),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_56),
.A2(n_43),
.B(n_35),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_3),
.B(n_4),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_54),
.B1(n_4),
.B2(n_5),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_68),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_67),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_2),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_71),
.Y(n_79)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_3),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_38),
.C(n_17),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_6),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_85),
.B1(n_7),
.B2(n_8),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_66),
.A2(n_54),
.B(n_60),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_83),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_10),
.B(n_11),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_6),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_73),
.A2(n_70),
.B1(n_72),
.B2(n_9),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_91),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_20),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_92),
.C(n_95),
.Y(n_98)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_23),
.C(n_28),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_97),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_24),
.C(n_27),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_79),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_76),
.C(n_82),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_102),
.C(n_32),
.Y(n_111)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_101),
.Y(n_107)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_103),
.A2(n_105),
.B(n_87),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_87),
.B(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_110),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_SL g110 ( 
.A1(n_100),
.A2(n_92),
.B(n_75),
.C(n_89),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_98),
.C(n_104),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_113),
.Y(n_115)
);

XNOR2x1_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_106),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_114),
.B(n_98),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_116),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_115),
.B(n_108),
.Y(n_118)
);

A2O1A1O1Ixp25_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_107),
.B(n_19),
.C(n_25),
.D(n_26),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_12),
.Y(n_120)
);


endmodule