module fake_jpeg_6771_n_222 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_222);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_222;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_SL g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_33),
.Y(n_45)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_34),
.Y(n_52)
);

AOI21xp33_ASAP7_75t_L g35 ( 
.A1(n_25),
.A2(n_0),
.B(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_1),
.Y(n_42)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx5_ASAP7_75t_SL g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_38),
.Y(n_50)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_15),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_15),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_42),
.B(n_31),
.Y(n_80)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_54),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_38),
.A2(n_40),
.B1(n_21),
.B2(n_27),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_44),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_21),
.B1(n_27),
.B2(n_20),
.Y(n_46)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_19),
.B1(n_28),
.B2(n_16),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_21),
.B1(n_20),
.B2(n_15),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_33),
.A2(n_20),
.B1(n_27),
.B2(n_17),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_51),
.A2(n_56),
.B1(n_57),
.B2(n_26),
.Y(n_74)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_23),
.B1(n_29),
.B2(n_17),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_18),
.B1(n_29),
.B2(n_23),
.Y(n_57)
);

CKINVDCx6p67_ASAP7_75t_R g58 ( 
.A(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_58),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_26),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_18),
.Y(n_68)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_31),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_63),
.B(n_76),
.Y(n_97)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_70),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_30),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_67),
.B(n_68),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_50),
.Y(n_70)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_74),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_30),
.Y(n_72)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_34),
.C(n_30),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_77),
.C(n_53),
.Y(n_93)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_79),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_28),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_45),
.C(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_25),
.Y(n_78)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_50),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_51),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_62),
.A2(n_47),
.B1(n_48),
.B2(n_44),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_76),
.B1(n_62),
.B2(n_77),
.Y(n_102)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_87),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_70),
.A2(n_53),
.B1(n_43),
.B2(n_47),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_46),
.B1(n_53),
.B2(n_79),
.Y(n_103)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_90),
.Y(n_104)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_92),
.B(n_101),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_77),
.C(n_73),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_57),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_74),
.Y(n_110)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_95),
.Y(n_106)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_100),
.B(n_74),
.Y(n_109)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_105),
.B1(n_112),
.B2(n_107),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_103),
.B(n_110),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_120),
.C(n_45),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_94),
.B(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_112),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_109),
.B(n_76),
.Y(n_140)
);

OA21x2_ASAP7_75t_L g111 ( 
.A1(n_85),
.A2(n_83),
.B(n_97),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_117),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_68),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_68),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_115),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_68),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_97),
.A2(n_76),
.B1(n_56),
.B2(n_59),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_72),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_67),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_65),
.C(n_52),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_86),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_118),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_122),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_110),
.A2(n_109),
.B(n_111),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_138),
.B1(n_115),
.B2(n_117),
.Y(n_149)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_106),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_126),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_127),
.B(n_103),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_114),
.B(n_96),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_128),
.B(n_130),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_106),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_102),
.B(n_91),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_136),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_119),
.A2(n_84),
.B(n_81),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_134),
.A2(n_135),
.B(n_113),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_111),
.A2(n_81),
.B(n_84),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_140),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_61),
.B(n_88),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_58),
.C(n_49),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_136),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_104),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_141),
.B(n_104),
.Y(n_150)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_151),
.C(n_155),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_145),
.A2(n_143),
.B(n_142),
.Y(n_169)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_146),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_134),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_132),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_149),
.A2(n_157),
.B1(n_158),
.B2(n_133),
.Y(n_162)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_127),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_135),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_153),
.Y(n_165)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_124),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_144),
.C(n_154),
.Y(n_176)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

AOI221xp5_ASAP7_75t_L g164 ( 
.A1(n_155),
.A2(n_138),
.B1(n_131),
.B2(n_143),
.C(n_140),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_164),
.A2(n_167),
.B(n_168),
.Y(n_178)
);

NOR2x1_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_133),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_167),
.B(n_170),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_173),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_152),
.A2(n_139),
.B1(n_121),
.B2(n_131),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_171),
.B(n_146),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_147),
.B(n_141),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_172),
.B(n_159),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_116),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_145),
.A2(n_158),
.B(n_157),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_78),
.B(n_49),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_178),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_185),
.Y(n_190)
);

BUFx12_ASAP7_75t_L g179 ( 
.A(n_172),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_183),
.Y(n_188)
);

INVxp33_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_182),
.A2(n_186),
.B(n_28),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_166),
.B(n_156),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_130),
.C(n_126),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_108),
.C(n_58),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_175),
.A2(n_165),
.B1(n_163),
.B2(n_171),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_189),
.A2(n_193),
.B(n_194),
.Y(n_203)
);

FAx1_ASAP7_75t_SL g191 ( 
.A(n_177),
.B(n_169),
.CI(n_174),
.CON(n_191),
.SN(n_191)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_180),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_181),
.A2(n_160),
.B1(n_173),
.B2(n_54),
.Y(n_192)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_192),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_108),
.C(n_95),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_87),
.C(n_98),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_195),
.B(n_196),
.Y(n_197)
);

AND2x6_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_180),
.Y(n_198)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_200),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_179),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_182),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_191),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_188),
.B(n_179),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_187),
.C(n_12),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_210),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_195),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_201),
.A2(n_194),
.B1(n_187),
.B2(n_59),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_208),
.A2(n_203),
.B1(n_197),
.B2(n_28),
.Y(n_212)
);

AOI322xp5_ASAP7_75t_L g215 ( 
.A1(n_212),
.A2(n_206),
.A3(n_209),
.B1(n_14),
.B2(n_16),
.C1(n_7),
.C2(n_9),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_92),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_214),
.A2(n_28),
.B(n_92),
.Y(n_216)
);

AOI322xp5_ASAP7_75t_L g218 ( 
.A1(n_215),
.A2(n_216),
.A3(n_217),
.B1(n_1),
.B2(n_2),
.C1(n_3),
.C2(n_6),
.Y(n_218)
);

AOI322xp5_ASAP7_75t_L g217 ( 
.A1(n_213),
.A2(n_211),
.A3(n_16),
.B1(n_3),
.B2(n_6),
.C1(n_7),
.C2(n_9),
.Y(n_217)
);

AOI221xp5_ASAP7_75t_SL g220 ( 
.A1(n_218),
.A2(n_219),
.B1(n_6),
.B2(n_9),
.C(n_10),
.Y(n_220)
);

AOI322xp5_ASAP7_75t_L g219 ( 
.A1(n_215),
.A2(n_211),
.A3(n_16),
.B1(n_59),
.B2(n_10),
.C1(n_11),
.C2(n_7),
.Y(n_219)
);

AOI221xp5_ASAP7_75t_L g221 ( 
.A1(n_220),
.A2(n_11),
.B1(n_75),
.B2(n_101),
.C(n_198),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_11),
.Y(n_222)
);


endmodule