module real_jpeg_31016_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_15),
.B1(n_20),
.B2(n_22),
.Y(n_19)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_1),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_1),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_2),
.A2(n_127),
.B1(n_129),
.B2(n_130),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_2),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_2),
.A2(n_129),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

OAI22x1_ASAP7_75t_SL g252 ( 
.A1(n_2),
.A2(n_129),
.B1(n_253),
.B2(n_260),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_2),
.A2(n_129),
.B1(n_396),
.B2(n_398),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_3),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_4),
.B(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_4),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_4),
.B(n_142),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g419 ( 
.A1(n_4),
.A2(n_273),
.B1(n_420),
.B2(n_422),
.Y(n_419)
);

OAI21xp33_ASAP7_75t_L g493 ( 
.A1(n_4),
.A2(n_230),
.B(n_444),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_5),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_5),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_5),
.A2(n_128),
.B1(n_214),
.B2(n_310),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_5),
.A2(n_214),
.B1(n_340),
.B2(n_344),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_6),
.A2(n_136),
.B1(n_137),
.B2(n_140),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_6),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_6),
.A2(n_136),
.B1(n_241),
.B2(n_247),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g410 ( 
.A1(n_6),
.A2(n_136),
.B1(n_411),
.B2(n_415),
.Y(n_410)
);

AOI22xp33_ASAP7_75t_L g452 ( 
.A1(n_6),
.A2(n_136),
.B1(n_453),
.B2(n_454),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_7),
.A2(n_224),
.B1(n_227),
.B2(n_229),
.Y(n_223)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_7),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_8),
.A2(n_40),
.B1(n_50),
.B2(n_54),
.Y(n_49)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_8),
.A2(n_54),
.B1(n_174),
.B2(n_178),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_9),
.A2(n_115),
.B1(n_119),
.B2(n_120),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_9),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_9),
.A2(n_119),
.B1(n_315),
.B2(n_319),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_9),
.A2(n_119),
.B1(n_369),
.B2(n_373),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_L g438 ( 
.A1(n_9),
.A2(n_119),
.B1(n_439),
.B2(n_442),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_10),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_10),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_11),
.Y(n_95)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_11),
.Y(n_101)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_12),
.Y(n_188)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_12),
.Y(n_466)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_13),
.Y(n_192)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_13),
.Y(n_196)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_13),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_14),
.A2(n_34),
.B1(n_35),
.B2(n_40),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_14),
.A2(n_34),
.B1(n_285),
.B2(n_289),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_16),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_16),
.Y(n_297)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_17),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_17),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_17),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_17),
.Y(n_259)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_18),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_18),
.Y(n_246)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_322),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_275),
.Y(n_23)
);

MAJx2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_171),
.C(n_232),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_26),
.B(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_85),
.Y(n_26)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_27),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_55),
.Y(n_27)
);

XNOR2x2_ASAP7_75t_SL g332 ( 
.A(n_28),
.B(n_56),
.Y(n_332)
);

AO22x1_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_33),
.B1(n_43),
.B2(n_48),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_32),
.Y(n_503)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_33),
.Y(n_231)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_39),
.Y(n_346)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_39),
.Y(n_401)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_42),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_42),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_42),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_43),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_43),
.B(n_395),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_43),
.A2(n_451),
.B1(n_455),
.B2(n_458),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_46),
.Y(n_43)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_44),
.Y(n_302)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g393 ( 
.A(n_45),
.Y(n_393)
);

INVx8_ASAP7_75t_L g446 ( 
.A(n_45),
.Y(n_446)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_46),
.Y(n_441)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22x1_ASAP7_75t_L g338 ( 
.A1(n_49),
.A2(n_230),
.B1(n_339),
.B2(n_347),
.Y(n_338)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_52),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_67),
.B1(n_73),
.B2(n_80),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_63),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_62),
.Y(n_272)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_66),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_66),
.Y(n_151)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_66),
.Y(n_160)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx2_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

NAND2xp33_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_77),
.Y(n_149)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVxp33_ASAP7_75t_L g274 ( 
.A(n_80),
.Y(n_274)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_84),
.Y(n_170)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_84),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_84),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_133),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_86),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_114),
.B(n_124),
.Y(n_86)
);

OAI22x1_ASAP7_75t_L g306 ( 
.A1(n_87),
.A2(n_238),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_87),
.A2(n_124),
.B(n_419),
.Y(n_418)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_88),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_88),
.B(n_126),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_102),
.Y(n_88)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_93),
.B1(n_96),
.B2(n_99),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_91),
.Y(n_217)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_92),
.Y(n_182)
);

INVx5_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_95),
.Y(n_391)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_98),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_98),
.Y(n_292)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_98),
.Y(n_372)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_105),
.B1(n_108),
.B2(n_112),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_114),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_115),
.A2(n_380),
.B1(n_383),
.B2(n_387),
.Y(n_379)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_116),
.B(n_388),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_125),
.Y(n_238)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_126),
.Y(n_307)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_133),
.B(n_279),
.C(n_280),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_152),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_142),
.Y(n_134)
);

AO22x1_ASAP7_75t_L g313 ( 
.A1(n_135),
.A2(n_142),
.B1(n_153),
.B2(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_139),
.A2(n_155),
.B1(n_159),
.B2(n_161),
.Y(n_154)
);

INVxp67_ASAP7_75t_SL g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_142),
.B(n_165),
.Y(n_266)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_146),
.B1(n_148),
.B2(n_150),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_147),
.Y(n_424)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_165),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_153),
.Y(n_268)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_167),
.Y(n_166)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_171),
.B(n_233),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_218),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_172),
.B(n_218),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_183),
.B1(n_197),
.B2(n_211),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_173),
.A2(n_183),
.B1(n_197),
.B2(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_176),
.Y(n_213)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

INVx5_ASAP7_75t_L g288 ( 
.A(n_182),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_183),
.A2(n_197),
.B1(n_368),
.B2(n_410),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_183),
.B(n_273),
.Y(n_498)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

AOI22x1_ASAP7_75t_L g251 ( 
.A1(n_184),
.A2(n_252),
.B1(n_263),
.B2(n_264),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_184),
.B(n_252),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_184),
.B(n_433),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_189),
.B1(n_193),
.B2(n_194),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx6_ASAP7_75t_L g301 ( 
.A(n_188),
.Y(n_301)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_188),
.Y(n_443)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_196),
.Y(n_201)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_197),
.Y(n_263)
);

OAI21xp33_ASAP7_75t_SL g367 ( 
.A1(n_197),
.A2(n_368),
.B(n_377),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_202),
.B1(n_205),
.B2(n_207),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_201),
.Y(n_479)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_204),
.Y(n_417)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_204),
.Y(n_490)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_211),
.Y(n_264)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_223),
.B1(n_230),
.B2(n_231),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_222),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_223),
.A2(n_230),
.B(n_294),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_224),
.Y(n_453)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx2_ASAP7_75t_SL g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_230),
.A2(n_438),
.B(n_444),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_250),
.C(n_265),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_235),
.B(n_251),
.Y(n_331)
);

AOI21x1_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B(n_239),
.Y(n_235)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI21xp33_ASAP7_75t_SL g335 ( 
.A1(n_238),
.A2(n_336),
.B(n_337),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_238),
.B(n_273),
.Y(n_435)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_240),
.Y(n_336)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_245),
.Y(n_249)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_245),
.Y(n_312)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_245),
.Y(n_421)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_252),
.B(n_263),
.Y(n_431)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx3_ASAP7_75t_SL g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_259),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_259),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_259),
.Y(n_414)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_263),
.B(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_265),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_273),
.B(n_274),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_273),
.B(n_381),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_273),
.B(n_384),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_273),
.B(n_481),
.Y(n_480)
);

OAI21xp33_ASAP7_75t_SL g487 ( 
.A1(n_273),
.A2(n_480),
.B(n_488),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_273),
.B(n_446),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_281),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_303),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_293),
.Y(n_282)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_288),
.Y(n_376)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_288),
.Y(n_386)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_302),
.Y(n_294)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_298),
.Y(n_496)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_301),
.Y(n_343)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_301),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_313),
.Y(n_305)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

OAI21xp33_ASAP7_75t_SL g322 ( 
.A1(n_323),
.A2(n_353),
.B(n_525),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_328),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_326),
.B(n_328),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_332),
.C(n_333),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_329),
.B(n_358),
.Y(n_357)
);

AND2x2_ASAP7_75t_SL g361 ( 
.A(n_329),
.B(n_358),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_332),
.A2(n_333),
.B1(n_334),
.B2(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_332),
.Y(n_359)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_338),
.C(n_351),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_335),
.B(n_365),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_338),
.B(n_352),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_339),
.A2(n_393),
.B(n_394),
.Y(n_392)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_344),
.Y(n_454)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

OAI21x1_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_402),
.B(n_523),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_360),
.B(n_362),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_357),
.B(n_361),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_362),
.B(n_524),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_366),
.C(n_378),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_363),
.A2(n_364),
.B1(n_518),
.B2(n_519),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_366),
.A2(n_367),
.B1(n_378),
.B2(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_372),
.Y(n_484)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

BUFx2_ASAP7_75t_L g469 ( 
.A(n_375),
.Y(n_469)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_377),
.B(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_378),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_392),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_379),
.B(n_392),
.Y(n_407)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

OAI21xp33_ASAP7_75t_L g499 ( 
.A1(n_394),
.A2(n_452),
.B(n_500),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_395),
.B(n_445),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx4_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

AOI21x1_ASAP7_75t_L g402 ( 
.A1(n_403),
.A2(n_514),
.B(n_521),
.Y(n_402)
);

OAI21x1_ASAP7_75t_L g403 ( 
.A1(n_404),
.A2(n_447),
.B(n_512),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_425),
.B(n_427),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_406),
.B(n_426),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_408),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_407),
.B(n_408),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_407),
.B(n_409),
.C(n_418),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_SL g408 ( 
.A(n_409),
.B(n_418),
.Y(n_408)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_410),
.Y(n_433)
);

INVx4_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx3_ASAP7_75t_SL g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_427),
.B(n_513),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_434),
.C(n_436),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_430),
.B(n_435),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_432),
.Y(n_430)
);

INVxp33_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_436),
.A2(n_437),
.B1(n_509),
.B2(n_510),
.Y(n_508)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_438),
.Y(n_458)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx5_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

AOI21x1_ASAP7_75t_L g447 ( 
.A1(n_448),
.A2(n_506),
.B(n_511),
.Y(n_447)
);

AO21x1_ASAP7_75t_SL g448 ( 
.A1(n_449),
.A2(n_491),
.B(n_505),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_459),
.Y(n_449)
);

NOR2xp67_ASAP7_75t_L g505 ( 
.A(n_450),
.B(n_459),
.Y(n_505)
);

INVxp33_ASAP7_75t_SL g451 ( 
.A(n_452),
.Y(n_451)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx5_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_485),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_R g507 ( 
.A(n_460),
.B(n_485),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_461),
.A2(n_467),
.B(n_475),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_463),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_470),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

AOI21xp33_ASAP7_75t_L g475 ( 
.A1(n_476),
.A2(n_478),
.B(n_480),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

BUFx4f_ASAP7_75t_SL g488 ( 
.A(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_492),
.A2(n_497),
.B(n_504),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_493),
.B(n_494),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_495),
.B(n_496),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_499),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_498),
.B(n_499),
.Y(n_504)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_503),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_508),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_507),
.B(n_508),
.Y(n_511)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_516),
.Y(n_514)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_515),
.Y(n_522)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

AND2x2_ASAP7_75t_SL g521 ( 
.A(n_517),
.B(n_522),
.Y(n_521)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);


endmodule