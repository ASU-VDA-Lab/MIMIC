module real_aes_2930_n_383 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_383);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_383;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_577;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_1014;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_974;
wire n_919;
wire n_857;
wire n_461;
wire n_1016;
wire n_908;
wire n_571;
wire n_549;
wire n_694;
wire n_491;
wire n_923;
wire n_894;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_742;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_963;
wire n_865;
wire n_666;
wire n_537;
wire n_884;
wire n_551;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_889;
wire n_955;
wire n_696;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_958;
wire n_677;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_994;
wire n_528;
wire n_578;
wire n_495;
wire n_892;
wire n_744;
wire n_384;
wire n_938;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_981;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_680;
wire n_595;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_529;
wire n_504;
wire n_725;
wire n_455;
wire n_960;
wire n_671;
wire n_973;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_817;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_885;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_1013;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_867;
wire n_745;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_488;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_727;
wire n_397;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_845;
wire n_850;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_637;
wire n_526;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_698;
wire n_541;
wire n_839;
wire n_639;
wire n_587;
wire n_546;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_988;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_842;
wire n_849;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_0), .A2(n_372), .B1(n_639), .B2(n_640), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g798 ( .A1(n_1), .A2(n_86), .B1(n_587), .B2(n_589), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_2), .A2(n_272), .B1(n_615), .B2(n_687), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_3), .A2(n_326), .B1(n_636), .B2(n_637), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_4), .A2(n_60), .B1(n_469), .B2(n_889), .Y(n_888) );
AOI22xp5_ASAP7_75t_L g922 ( .A1(n_5), .A2(n_107), .B1(n_469), .B2(n_923), .Y(n_922) );
AOI22xp5_ASAP7_75t_L g1003 ( .A1(n_6), .A2(n_151), .B1(n_525), .B2(n_527), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_7), .A2(n_274), .B1(n_670), .B2(n_776), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_8), .A2(n_38), .B1(n_452), .B2(n_486), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_9), .A2(n_347), .B1(n_435), .B2(n_650), .Y(n_766) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_10), .A2(n_29), .B1(n_497), .B2(n_730), .Y(n_835) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_11), .A2(n_317), .B1(n_564), .B2(n_653), .Y(n_671) );
XOR2x2_ASAP7_75t_L g521 ( .A(n_12), .B(n_522), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_13), .A2(n_88), .B1(n_525), .B2(n_616), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_14), .A2(n_111), .B1(n_447), .B2(n_530), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g857 ( .A1(n_15), .A2(n_76), .B1(n_645), .B2(n_673), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_16), .A2(n_98), .B1(n_539), .B2(n_540), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g880 ( .A(n_17), .Y(n_880) );
AOI22xp33_ASAP7_75t_SL g818 ( .A1(n_18), .A2(n_379), .B1(n_632), .B2(n_782), .Y(n_818) );
AOI22xp33_ASAP7_75t_SL g665 ( .A1(n_19), .A2(n_260), .B1(n_666), .B2(n_667), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_20), .A2(n_211), .B1(n_414), .B2(n_561), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_21), .A2(n_49), .B1(n_424), .B2(n_953), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_22), .A2(n_187), .B1(n_434), .B2(n_566), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_23), .A2(n_126), .B1(n_640), .B2(n_662), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_24), .A2(n_130), .B1(n_504), .B2(n_527), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_25), .A2(n_370), .B1(n_513), .B2(n_559), .Y(n_767) );
AO22x2_ASAP7_75t_L g546 ( .A1(n_26), .A2(n_547), .B1(n_567), .B2(n_568), .Y(n_546) );
INVx1_ASAP7_75t_L g567 ( .A(n_26), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_27), .A2(n_189), .B1(n_650), .B2(n_651), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_28), .A2(n_237), .B1(n_540), .B2(n_561), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_30), .A2(n_174), .B1(n_587), .B2(n_589), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_31), .B(n_465), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_32), .A2(n_127), .B1(n_504), .B2(n_527), .Y(n_799) );
INVx1_ASAP7_75t_SL g411 ( .A(n_33), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g980 ( .A(n_33), .B(n_46), .Y(n_980) );
INVx1_ASAP7_75t_L g942 ( .A(n_34), .Y(n_942) );
AOI222xp33_ASAP7_75t_L g542 ( .A1(n_35), .A2(n_322), .B1(n_374), .B2(n_543), .C1(n_544), .C2(n_545), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_36), .A2(n_233), .B1(n_539), .B2(n_540), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_37), .A2(n_51), .B1(n_647), .B2(n_867), .Y(n_892) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_39), .A2(n_331), .B1(n_459), .B2(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_40), .B(n_465), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_41), .A2(n_197), .B1(n_639), .B2(n_640), .Y(n_908) );
AOI22xp5_ASAP7_75t_L g853 ( .A1(n_42), .A2(n_84), .B1(n_636), .B2(n_637), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_43), .B(n_580), .Y(n_874) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_44), .A2(n_229), .B1(n_669), .B2(n_670), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_45), .B(n_629), .Y(n_852) );
AO22x2_ASAP7_75t_L g406 ( .A1(n_46), .A2(n_360), .B1(n_400), .B2(n_407), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_47), .A2(n_204), .B1(n_584), .B2(n_712), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_48), .B(n_629), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_50), .B(n_465), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_52), .A2(n_120), .B1(n_504), .B2(n_505), .Y(n_503) );
AO22x1_ASAP7_75t_L g436 ( .A1(n_53), .A2(n_357), .B1(n_437), .B2(n_440), .Y(n_436) );
INVx1_ASAP7_75t_L g412 ( .A(n_54), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_55), .A2(n_236), .B1(n_540), .B2(n_561), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_56), .A2(n_100), .B1(n_564), .B2(n_667), .Y(n_915) );
OAI22xp5_ASAP7_75t_L g1010 ( .A1(n_57), .A2(n_1011), .B1(n_1012), .B2(n_1013), .Y(n_1010) );
CKINVDCx20_ASAP7_75t_R g1011 ( .A(n_57), .Y(n_1011) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_58), .A2(n_212), .B1(n_447), .B2(n_550), .Y(n_549) );
AOI22xp33_ASAP7_75t_SL g756 ( .A1(n_59), .A2(n_333), .B1(n_554), .B2(n_704), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_61), .A2(n_191), .B1(n_589), .B2(n_870), .Y(n_869) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_62), .A2(n_137), .B1(n_513), .B2(n_559), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_63), .A2(n_368), .B1(n_517), .B2(n_584), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g957 ( .A1(n_64), .A2(n_290), .B1(n_434), .B2(n_958), .Y(n_957) );
XNOR2x1_ASAP7_75t_L g918 ( .A(n_65), .B(n_919), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g933 ( .A1(n_65), .A2(n_919), .B1(n_934), .B2(n_935), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_65), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_66), .A2(n_350), .B1(n_536), .B2(n_802), .Y(n_1001) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_67), .A2(n_245), .B1(n_645), .B2(n_673), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_68), .A2(n_170), .B1(n_636), .B2(n_817), .Y(n_816) );
AOI21xp5_ASAP7_75t_SL g445 ( .A1(n_69), .A2(n_446), .B(n_449), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_70), .A2(n_171), .B1(n_515), .B2(n_517), .Y(n_514) );
AO22x2_ASAP7_75t_L g399 ( .A1(n_71), .A2(n_181), .B1(n_400), .B2(n_401), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_72), .A2(n_354), .B1(n_424), .B2(n_714), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_73), .A2(n_146), .B1(n_536), .B2(n_537), .Y(n_620) );
AOI22xp33_ASAP7_75t_SL g643 ( .A1(n_74), .A2(n_136), .B1(n_644), .B2(n_645), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_75), .A2(n_153), .B1(n_505), .B2(n_594), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_77), .A2(n_149), .B1(n_419), .B2(n_764), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_78), .A2(n_230), .B1(n_434), .B2(n_566), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_79), .A2(n_336), .B1(n_632), .B2(n_633), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g836 ( .A1(n_80), .A2(n_223), .B1(n_470), .B2(n_492), .Y(n_836) );
AOI222xp33_ASAP7_75t_L g815 ( .A1(n_81), .A2(n_92), .B1(n_193), .B2(n_629), .C1(n_639), .C2(n_784), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_82), .A2(n_283), .B1(n_564), .B2(n_653), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_83), .A2(n_195), .B1(n_653), .B2(n_670), .Y(n_914) );
AOI22xp5_ASAP7_75t_L g837 ( .A1(n_85), .A2(n_380), .B1(n_639), .B2(n_784), .Y(n_837) );
AOI22xp33_ASAP7_75t_SL g875 ( .A1(n_87), .A2(n_239), .B1(n_472), .B2(n_876), .Y(n_875) );
AO222x2_ASAP7_75t_SL g609 ( .A1(n_89), .A2(n_288), .B1(n_343), .B2(n_492), .C1(n_610), .C2(n_611), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_90), .A2(n_168), .B1(n_457), .B2(n_947), .Y(n_946) );
AOI22xp5_ASAP7_75t_L g831 ( .A1(n_91), .A2(n_140), .B1(n_413), .B2(n_644), .Y(n_831) );
AOI22xp5_ASAP7_75t_L g822 ( .A1(n_93), .A2(n_118), .B1(n_645), .B2(n_673), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g860 ( .A1(n_94), .A2(n_210), .B1(n_564), .B2(n_667), .Y(n_860) );
OA22x2_ASAP7_75t_L g810 ( .A1(n_95), .A2(n_811), .B1(n_812), .B2(n_813), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_95), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_96), .A2(n_207), .B1(n_539), .B2(n_589), .Y(n_1002) );
AOI22xp5_ASAP7_75t_L g823 ( .A1(n_97), .A2(n_104), .B1(n_667), .B2(n_670), .Y(n_823) );
AOI22xp5_ASAP7_75t_L g859 ( .A1(n_99), .A2(n_294), .B1(n_653), .B2(n_670), .Y(n_859) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_101), .A2(n_133), .B1(n_513), .B2(n_647), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_102), .A2(n_221), .B1(n_505), .B2(n_650), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_103), .A2(n_361), .B1(n_645), .B2(n_673), .Y(n_774) );
AO22x1_ASAP7_75t_L g429 ( .A1(n_105), .A2(n_359), .B1(n_430), .B2(n_434), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_106), .A2(n_232), .B1(n_564), .B2(n_653), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_108), .A2(n_258), .B1(n_460), .B2(n_706), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_109), .A2(n_340), .B1(n_532), .B2(n_806), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_110), .A2(n_257), .B1(n_761), .B2(n_762), .Y(n_760) );
AOI22xp5_ASAP7_75t_L g873 ( .A1(n_112), .A2(n_143), .B1(n_446), .B2(n_499), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_113), .A2(n_363), .B1(n_442), .B2(n_653), .Y(n_829) );
AOI22xp5_ASAP7_75t_L g904 ( .A1(n_114), .A2(n_215), .B1(n_632), .B2(n_633), .Y(n_904) );
AO22x2_ASAP7_75t_L g403 ( .A1(n_115), .A2(n_287), .B1(n_400), .B2(n_404), .Y(n_403) );
AOI222xp33_ASAP7_75t_SL g928 ( .A1(n_116), .A2(n_275), .B1(n_353), .B2(n_456), .C1(n_465), .C2(n_806), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_117), .A2(n_219), .B1(n_615), .B2(n_616), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_119), .A2(n_352), .B1(n_456), .B2(n_459), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_121), .A2(n_226), .B1(n_532), .B2(n_533), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_122), .A2(n_301), .B1(n_394), .B2(n_413), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_123), .A2(n_289), .B1(n_559), .B2(n_764), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_124), .A2(n_335), .B1(n_510), .B2(n_591), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g1004 ( .A1(n_125), .A2(n_342), .B1(n_504), .B2(n_512), .Y(n_1004) );
AOI22xp5_ASAP7_75t_L g858 ( .A1(n_128), .A2(n_164), .B1(n_666), .B2(n_776), .Y(n_858) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_129), .A2(n_323), .B1(n_563), .B2(n_564), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_131), .A2(n_205), .B1(n_587), .B2(n_589), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_132), .A2(n_209), .B1(n_533), .B2(n_553), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_134), .A2(n_366), .B1(n_456), .B2(n_725), .Y(n_887) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_135), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_138), .A2(n_206), .B1(n_505), .B2(n_525), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_139), .A2(n_277), .B1(n_647), .B2(n_712), .Y(n_871) );
AOI22xp33_ASAP7_75t_SL g635 ( .A1(n_141), .A2(n_172), .B1(n_636), .B2(n_637), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_142), .A2(n_306), .B1(n_666), .B2(n_669), .Y(n_830) );
INVx1_ASAP7_75t_L g989 ( .A(n_144), .Y(n_989) );
AO22x1_ASAP7_75t_L g418 ( .A1(n_145), .A2(n_238), .B1(n_419), .B2(n_424), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g996 ( .A1(n_147), .A2(n_303), .B1(n_447), .B2(n_607), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_148), .A2(n_244), .B1(n_459), .B2(n_575), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_150), .A2(n_327), .B1(n_470), .B2(n_474), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_152), .B(n_580), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_154), .A2(n_346), .B1(n_645), .B2(n_673), .Y(n_911) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_155), .A2(n_270), .B1(n_632), .B2(n_782), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_156), .B(n_543), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_157), .A2(n_203), .B1(n_553), .B2(n_554), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_158), .A2(n_316), .B1(n_632), .B2(n_633), .Y(n_660) );
AO21x2_ASAP7_75t_L g721 ( .A1(n_159), .A2(n_722), .B(n_745), .Y(n_721) );
INVx1_ASAP7_75t_L g747 ( .A(n_159), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_160), .A2(n_253), .B1(n_536), .B2(n_802), .Y(n_801) );
AO22x2_ASAP7_75t_L g770 ( .A1(n_161), .A2(n_771), .B1(n_786), .B2(n_787), .Y(n_770) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_161), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_162), .A2(n_324), .B1(n_587), .B2(n_744), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_163), .B(n_692), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_165), .A2(n_182), .B1(n_587), .B2(n_589), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_166), .B(n_483), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_167), .A2(n_351), .B1(n_495), .B2(n_499), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_169), .A2(n_304), .B1(n_632), .B2(n_633), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_173), .A2(n_278), .B1(n_662), .B2(n_784), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_175), .A2(n_325), .B1(n_470), .B2(n_924), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_176), .A2(n_213), .B1(n_497), .B2(n_607), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_177), .A2(n_224), .B1(n_489), .B2(n_492), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_178), .A2(n_199), .B1(n_447), .B2(n_530), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_179), .A2(n_281), .B1(n_430), .B2(n_740), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_180), .A2(n_235), .B1(n_640), .B2(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g979 ( .A(n_181), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g997 ( .A1(n_183), .A2(n_328), .B1(n_457), .B2(n_806), .Y(n_997) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_184), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_185), .A2(n_297), .B1(n_495), .B2(n_499), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_186), .A2(n_284), .B1(n_575), .B2(n_729), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_188), .A2(n_337), .B1(n_510), .B2(n_512), .Y(n_800) );
AO222x2_ASAP7_75t_SL g724 ( .A1(n_190), .A2(n_282), .B1(n_344), .B2(n_465), .C1(n_486), .C2(n_725), .Y(n_724) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_192), .A2(n_299), .B1(n_666), .B2(n_776), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_194), .A2(n_381), .B1(n_564), .B2(n_653), .Y(n_652) );
OA22x2_ASAP7_75t_L g389 ( .A1(n_196), .A2(n_390), .B1(n_391), .B2(n_477), .Y(n_389) );
INVx1_ASAP7_75t_L g477 ( .A(n_196), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_198), .A2(n_255), .B1(n_564), .B2(n_647), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_200), .A2(n_252), .B1(n_636), .B2(n_637), .Y(n_785) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_201), .A2(n_320), .B1(n_711), .B2(n_712), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_202), .B(n_629), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_208), .A2(n_285), .B1(n_544), .B2(n_545), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_214), .A2(n_218), .B1(n_486), .B2(n_487), .Y(n_485) );
XOR2x2_ASAP7_75t_L g656 ( .A(n_216), .B(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_217), .B(n_580), .Y(n_579) );
XNOR2x1_ASAP7_75t_L g679 ( .A(n_220), .B(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g986 ( .A(n_222), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_225), .A2(n_307), .B1(n_550), .B2(n_706), .Y(n_705) );
XOR2x2_ASAP7_75t_L g993 ( .A(n_227), .B(n_994), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_227), .A2(n_1009), .B1(n_1010), .B2(n_1014), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_228), .A2(n_296), .B1(n_725), .B2(n_878), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_231), .A2(n_382), .B1(n_650), .B2(n_740), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_234), .A2(n_377), .B1(n_533), .B2(n_553), .Y(n_608) );
AOI22xp33_ASAP7_75t_SL g949 ( .A1(n_240), .A2(n_365), .B1(n_730), .B2(n_950), .Y(n_949) );
CKINVDCx20_ASAP7_75t_R g630 ( .A(n_241), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_242), .A2(n_250), .B1(n_544), .B2(n_545), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_243), .A2(n_341), .B1(n_584), .B2(n_712), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_246), .B(n_780), .Y(n_779) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_247), .A2(n_293), .B1(n_533), .B2(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g479 ( .A(n_248), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_249), .A2(n_314), .B1(n_489), .B2(n_545), .Y(n_695) );
XNOR2x1_ASAP7_75t_L g849 ( .A(n_251), .B(n_850), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_254), .A2(n_286), .B1(n_645), .B2(n_673), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_256), .A2(n_295), .B1(n_866), .B2(n_867), .Y(n_865) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_259), .Y(n_734) );
XOR2x2_ASAP7_75t_L g571 ( .A(n_261), .B(n_572), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_262), .A2(n_378), .B1(n_470), .B2(n_492), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_263), .A2(n_334), .B1(n_459), .B2(n_497), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_264), .A2(n_373), .B1(n_684), .B2(n_711), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_265), .A2(n_371), .B1(n_594), .B2(n_740), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_266), .A2(n_271), .B1(n_413), .B2(n_507), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_267), .A2(n_311), .B1(n_536), .B2(n_537), .Y(n_535) );
XNOR2x1_ASAP7_75t_L g698 ( .A(n_268), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g654 ( .A(n_269), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_273), .A2(n_348), .B1(n_474), .B2(n_611), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_276), .A2(n_291), .B1(n_512), .B2(n_525), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_279), .A2(n_319), .B1(n_666), .B2(n_669), .Y(n_912) );
OA22x2_ASAP7_75t_L g824 ( .A1(n_280), .A2(n_825), .B1(n_826), .B2(n_838), .Y(n_824) );
INVx1_ASAP7_75t_L g838 ( .A(n_280), .Y(n_838) );
NOR2xp33_ASAP7_75t_L g977 ( .A(n_287), .B(n_978), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_292), .A2(n_356), .B1(n_566), .B2(n_955), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_298), .A2(n_318), .B1(n_544), .B2(n_545), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_300), .A2(n_330), .B1(n_437), .B2(n_666), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_302), .A2(n_339), .B1(n_474), .B2(n_491), .Y(n_754) );
AOI22xp5_ASAP7_75t_L g468 ( .A1(n_305), .A2(n_338), .B1(n_469), .B2(n_472), .Y(n_468) );
INVx3_ASAP7_75t_L g400 ( .A(n_308), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_309), .A2(n_329), .B1(n_536), .B2(n_684), .Y(n_683) );
XOR2x1_ASAP7_75t_L g883 ( .A(n_310), .B(n_884), .Y(n_883) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_312), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_313), .A2(n_345), .B1(n_510), .B2(n_512), .Y(n_509) );
OA22x2_ASAP7_75t_L g793 ( .A1(n_315), .A2(n_794), .B1(n_795), .B2(n_796), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_315), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_321), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_332), .B(n_465), .Y(n_834) );
AO22x2_ASAP7_75t_L g603 ( .A1(n_349), .A2(n_604), .B1(n_621), .B2(n_622), .Y(n_603) );
INVx1_ASAP7_75t_L g622 ( .A(n_349), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g907 ( .A1(n_355), .A2(n_364), .B1(n_636), .B2(n_817), .Y(n_907) );
INVx1_ASAP7_75t_L g916 ( .A(n_358), .Y(n_916) );
NAND2xp5_ASAP7_75t_SL g999 ( .A(n_362), .B(n_483), .Y(n_999) );
INVx1_ASAP7_75t_L g974 ( .A(n_367), .Y(n_974) );
AND2x4_ASAP7_75t_L g988 ( .A(n_367), .B(n_975), .Y(n_988) );
AO21x1_ASAP7_75t_L g1015 ( .A1(n_367), .A2(n_984), .B(n_1016), .Y(n_1015) );
INVx1_ASAP7_75t_L g975 ( .A(n_369), .Y(n_975) );
AND2x2_ASAP7_75t_R g1009 ( .A(n_369), .B(n_974), .Y(n_1009) );
INVxp67_ASAP7_75t_L g985 ( .A(n_375), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g948 ( .A(n_376), .B(n_780), .Y(n_948) );
O2A1O1Ixp33_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_716), .B(n_970), .C(n_981), .Y(n_383) );
AOI21xp33_ASAP7_75t_L g970 ( .A1(n_384), .A2(n_716), .B(n_971), .Y(n_970) );
XOR2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_598), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B1(n_519), .B2(n_597), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AOI22xp33_ASAP7_75t_R g387 ( .A1(n_388), .A2(n_389), .B1(n_478), .B2(n_518), .Y(n_387) );
INVx2_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NOR2xp67_ASAP7_75t_L g391 ( .A(n_392), .B(n_444), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_417), .Y(n_392) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g508 ( .A(n_395), .Y(n_508) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_395), .Y(n_539) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g588 ( .A(n_396), .Y(n_588) );
INVx1_ASAP7_75t_L g761 ( .A(n_396), .Y(n_761) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_397), .Y(n_561) );
BUFx3_ASAP7_75t_L g644 ( .A(n_397), .Y(n_644) );
AND2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_405), .Y(n_397) );
AND2x4_ASAP7_75t_L g426 ( .A(n_398), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g448 ( .A(n_398), .B(n_433), .Y(n_448) );
AND2x6_ASAP7_75t_L g564 ( .A(n_398), .B(n_427), .Y(n_564) );
AND2x4_ASAP7_75t_L g636 ( .A(n_398), .B(n_433), .Y(n_636) );
AND2x2_ASAP7_75t_L g673 ( .A(n_398), .B(n_405), .Y(n_673) );
AND2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_402), .Y(n_398) );
AND2x2_ASAP7_75t_L g416 ( .A(n_399), .B(n_403), .Y(n_416) );
INVx2_ASAP7_75t_L g423 ( .A(n_399), .Y(n_423) );
INVx1_ASAP7_75t_L g401 ( .A(n_400), .Y(n_401) );
INVx2_ASAP7_75t_L g404 ( .A(n_400), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_400), .Y(n_407) );
OAI22x1_ASAP7_75t_L g409 ( .A1(n_400), .A2(n_410), .B1(n_411), .B2(n_412), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_400), .Y(n_410) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_402), .Y(n_463) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g422 ( .A(n_403), .Y(n_422) );
AND2x4_ASAP7_75t_L g443 ( .A(n_403), .B(n_423), .Y(n_443) );
AND2x2_ASAP7_75t_L g420 ( .A(n_405), .B(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g458 ( .A(n_405), .B(n_443), .Y(n_458) );
AND2x2_ASAP7_75t_L g639 ( .A(n_405), .B(n_443), .Y(n_639) );
AND2x6_ASAP7_75t_L g653 ( .A(n_405), .B(n_421), .Y(n_653) );
AND2x2_ASAP7_75t_L g662 ( .A(n_405), .B(n_443), .Y(n_662) );
AND2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_408), .Y(n_405) );
BUFx2_ASAP7_75t_L g415 ( .A(n_406), .Y(n_415) );
INVx2_ASAP7_75t_L g428 ( .A(n_406), .Y(n_428) );
AND2x2_ASAP7_75t_L g454 ( .A(n_406), .B(n_409), .Y(n_454) );
AND2x4_ASAP7_75t_L g427 ( .A(n_408), .B(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g433 ( .A(n_409), .B(n_428), .Y(n_433) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_409), .Y(n_476) );
BUFx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx5_ASAP7_75t_SL g541 ( .A(n_414), .Y(n_541) );
AND2x4_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
AND2x4_ASAP7_75t_L g645 ( .A(n_415), .B(n_416), .Y(n_645) );
AND2x4_ASAP7_75t_L g435 ( .A(n_416), .B(n_427), .Y(n_435) );
AND2x2_ASAP7_75t_L g475 ( .A(n_416), .B(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_SL g633 ( .A(n_416), .B(n_476), .Y(n_633) );
AND2x4_ASAP7_75t_L g666 ( .A(n_416), .B(n_427), .Y(n_666) );
AND2x2_ASAP7_75t_SL g782 ( .A(n_416), .B(n_476), .Y(n_782) );
NOR3xp33_ASAP7_75t_L g417 ( .A(n_418), .B(n_429), .C(n_436), .Y(n_417) );
BUFx3_ASAP7_75t_L g866 ( .A(n_419), .Y(n_866) );
BUFx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx3_ASAP7_75t_L g516 ( .A(n_420), .Y(n_516) );
BUFx2_ASAP7_75t_L g563 ( .A(n_420), .Y(n_563) );
AND2x4_ASAP7_75t_L g432 ( .A(n_421), .B(n_433), .Y(n_432) );
AND2x4_ASAP7_75t_L g439 ( .A(n_421), .B(n_427), .Y(n_439) );
AND2x2_ASAP7_75t_L g467 ( .A(n_421), .B(n_454), .Y(n_467) );
AND2x4_ASAP7_75t_L g629 ( .A(n_421), .B(n_454), .Y(n_629) );
AND2x2_ASAP7_75t_L g667 ( .A(n_421), .B(n_427), .Y(n_667) );
AND2x2_ASAP7_75t_L g669 ( .A(n_421), .B(n_433), .Y(n_669) );
AND2x2_ASAP7_75t_L g776 ( .A(n_421), .B(n_433), .Y(n_776) );
AND2x4_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
INVxp67_ASAP7_75t_L g453 ( .A(n_423), .Y(n_453) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g517 ( .A(n_425), .Y(n_517) );
INVx1_ASAP7_75t_SL g537 ( .A(n_425), .Y(n_537) );
INVx2_ASAP7_75t_SL g684 ( .A(n_425), .Y(n_684) );
INVx2_ASAP7_75t_L g764 ( .A(n_425), .Y(n_764) );
INVx2_ASAP7_75t_L g802 ( .A(n_425), .Y(n_802) );
INVx2_ASAP7_75t_SL g867 ( .A(n_425), .Y(n_867) );
INVx8_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND2x4_ASAP7_75t_L g442 ( .A(n_427), .B(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g670 ( .A(n_427), .B(n_443), .Y(n_670) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g504 ( .A(n_431), .Y(n_504) );
INVx1_ASAP7_75t_SL g594 ( .A(n_431), .Y(n_594) );
INVx2_ASAP7_75t_L g615 ( .A(n_431), .Y(n_615) );
INVx6_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx3_ASAP7_75t_L g566 ( .A(n_432), .Y(n_566) );
BUFx3_ASAP7_75t_L g650 ( .A(n_432), .Y(n_650) );
AND2x2_ASAP7_75t_L g471 ( .A(n_433), .B(n_443), .Y(n_471) );
AND2x4_ASAP7_75t_L g632 ( .A(n_433), .B(n_443), .Y(n_632) );
BUFx3_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx2_ASAP7_75t_SL g505 ( .A(n_435), .Y(n_505) );
BUFx2_ASAP7_75t_SL g527 ( .A(n_435), .Y(n_527) );
BUFx3_ASAP7_75t_L g651 ( .A(n_435), .Y(n_651) );
INVx2_ASAP7_75t_L g688 ( .A(n_435), .Y(n_688) );
INVx2_ASAP7_75t_L g511 ( .A(n_437), .Y(n_511) );
BUFx6f_ASAP7_75t_L g525 ( .A(n_437), .Y(n_525) );
INVx4_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g559 ( .A(n_438), .Y(n_559) );
INVx3_ASAP7_75t_SL g647 ( .A(n_438), .Y(n_647) );
INVx3_ASAP7_75t_L g714 ( .A(n_438), .Y(n_714) );
INVx2_ASAP7_75t_SL g958 ( .A(n_438), .Y(n_958) );
INVx8_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g616 ( .A(n_441), .Y(n_616) );
INVx1_ASAP7_75t_L g712 ( .A(n_441), .Y(n_712) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_442), .Y(n_513) );
BUFx3_ASAP7_75t_L g737 ( .A(n_442), .Y(n_737) );
BUFx6f_ASAP7_75t_L g955 ( .A(n_442), .Y(n_955) );
NAND4xp25_ASAP7_75t_L g444 ( .A(n_445), .B(n_455), .C(n_464), .D(n_468), .Y(n_444) );
BUFx6f_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx3_ASAP7_75t_L g498 ( .A(n_448), .Y(n_498) );
BUFx6f_ASAP7_75t_L g706 ( .A(n_448), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
INVx2_ASAP7_75t_L g487 ( .A(n_451), .Y(n_487) );
INVx2_ASAP7_75t_SL g533 ( .A(n_451), .Y(n_533) );
INVx2_ASAP7_75t_L g554 ( .A(n_451), .Y(n_554) );
INVx2_ASAP7_75t_L g725 ( .A(n_451), .Y(n_725) );
INVx2_ASAP7_75t_L g806 ( .A(n_451), .Y(n_806) );
INVx1_ASAP7_75t_L g947 ( .A(n_451), .Y(n_947) );
INVx6_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
AND2x2_ASAP7_75t_L g640 ( .A(n_453), .B(n_454), .Y(n_640) );
AND2x2_ASAP7_75t_L g784 ( .A(n_453), .B(n_454), .Y(n_784) );
AND2x4_ASAP7_75t_L g461 ( .A(n_454), .B(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g637 ( .A(n_454), .B(n_462), .Y(n_637) );
AND2x2_ASAP7_75t_L g817 ( .A(n_454), .B(n_462), .Y(n_817) );
BUFx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx2_ASAP7_75t_L g486 ( .A(n_457), .Y(n_486) );
BUFx4f_ASAP7_75t_SL g532 ( .A(n_457), .Y(n_532) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx3_ASAP7_75t_L g553 ( .A(n_458), .Y(n_553) );
BUFx2_ASAP7_75t_L g704 ( .A(n_458), .Y(n_704) );
BUFx6f_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
BUFx3_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g501 ( .A(n_461), .Y(n_501) );
BUFx4f_ASAP7_75t_L g530 ( .A(n_461), .Y(n_530) );
INVx1_ASAP7_75t_L g551 ( .A(n_461), .Y(n_551) );
BUFx6f_ASAP7_75t_SL g730 ( .A(n_461), .Y(n_730) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx3_ASAP7_75t_SL g484 ( .A(n_466), .Y(n_484) );
INVx4_ASAP7_75t_SL g543 ( .A(n_466), .Y(n_543) );
INVx3_ASAP7_75t_L g610 ( .A(n_466), .Y(n_610) );
BUFx2_ASAP7_75t_L g693 ( .A(n_466), .Y(n_693) );
INVx4_ASAP7_75t_SL g780 ( .A(n_466), .Y(n_780) );
INVx6_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx3_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx3_ASAP7_75t_L g491 ( .A(n_471), .Y(n_491) );
INVx2_ASAP7_75t_L g612 ( .A(n_471), .Y(n_612) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx3_ASAP7_75t_L g889 ( .A(n_474), .Y(n_889) );
BUFx12f_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx3_ASAP7_75t_L g493 ( .A(n_475), .Y(n_493) );
INVx2_ASAP7_75t_L g518 ( .A(n_478), .Y(n_518) );
XNOR2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
NOR2x1_ASAP7_75t_L g480 ( .A(n_481), .B(n_502), .Y(n_480) );
NAND4xp25_ASAP7_75t_SL g481 ( .A(n_482), .B(n_485), .C(n_488), .D(n_494), .Y(n_481) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g581 ( .A(n_484), .Y(n_581) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx6f_ASAP7_75t_SL g544 ( .A(n_491), .Y(n_544) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_492), .Y(n_545) );
INVx3_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g924 ( .A(n_493), .Y(n_924) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
INVx4_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g576 ( .A(n_498), .Y(n_576) );
INVx2_ASAP7_75t_L g950 ( .A(n_498), .Y(n_950) );
INVx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g607 ( .A(n_501), .Y(n_607) );
NAND4xp25_ASAP7_75t_L g502 ( .A(n_503), .B(n_506), .C(n_509), .D(n_514), .Y(n_502) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx6f_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g592 ( .A(n_513), .Y(n_592) );
INVx2_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_SL g536 ( .A(n_516), .Y(n_536) );
INVx3_ASAP7_75t_L g711 ( .A(n_516), .Y(n_711) );
INVx2_ASAP7_75t_L g953 ( .A(n_516), .Y(n_953) );
INVxp67_ASAP7_75t_L g597 ( .A(n_519), .Y(n_597) );
AOI22x1_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_571), .B1(n_595), .B2(n_596), .Y(n_519) );
INVx2_ASAP7_75t_SL g596 ( .A(n_520), .Y(n_596) );
OA22x2_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_546), .B1(n_569), .B2(n_570), .Y(n_520) );
INVx2_ASAP7_75t_SL g569 ( .A(n_521), .Y(n_569) );
NAND4xp75_ASAP7_75t_SL g522 ( .A(n_523), .B(n_528), .C(n_534), .D(n_542), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_526), .Y(n_523) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .Y(n_528) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_538), .Y(n_534) );
INVx3_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g589 ( .A(n_541), .Y(n_589) );
INVx2_ASAP7_75t_L g744 ( .A(n_541), .Y(n_744) );
INVx2_ASAP7_75t_L g762 ( .A(n_541), .Y(n_762) );
INVx2_ASAP7_75t_L g570 ( .A(n_546), .Y(n_570) );
INVx1_ASAP7_75t_L g568 ( .A(n_547), .Y(n_568) );
NOR2x1_ASAP7_75t_L g547 ( .A(n_548), .B(n_557), .Y(n_547) );
NAND4xp25_ASAP7_75t_L g548 ( .A(n_549), .B(n_552), .C(n_555), .D(n_556), .Y(n_548) );
INVx2_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g879 ( .A(n_553), .Y(n_879) );
NAND4xp25_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .C(n_562), .D(n_565), .Y(n_557) );
INVx1_ASAP7_75t_L g733 ( .A(n_559), .Y(n_733) );
INVx2_ASAP7_75t_L g585 ( .A(n_563), .Y(n_585) );
INVx1_ASAP7_75t_L g595 ( .A(n_571), .Y(n_595) );
NOR2x1_ASAP7_75t_L g572 ( .A(n_573), .B(n_582), .Y(n_572) );
NAND4xp25_ASAP7_75t_L g573 ( .A(n_574), .B(n_577), .C(n_578), .D(n_579), .Y(n_573) );
BUFx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OAI21xp33_ASAP7_75t_SL g752 ( .A1(n_581), .A2(n_753), .B(n_754), .Y(n_752) );
NAND4xp25_ASAP7_75t_L g582 ( .A(n_583), .B(n_586), .C(n_590), .D(n_593), .Y(n_582) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_601), .B1(n_676), .B2(n_715), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_603), .B1(n_623), .B2(n_675), .Y(n_601) );
INVx2_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_SL g621 ( .A(n_604), .Y(n_621) );
NOR4xp75_ASAP7_75t_L g604 ( .A(n_605), .B(n_609), .C(n_613), .D(n_618), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g876 ( .A(n_612), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_617), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
INVx2_ASAP7_75t_L g675 ( .A(n_623), .Y(n_675) );
OA22x2_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_655), .B1(n_656), .B2(n_674), .Y(n_623) );
INVx1_ASAP7_75t_L g674 ( .A(n_624), .Y(n_674) );
XOR2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_654), .Y(n_624) );
NAND2x1_ASAP7_75t_L g625 ( .A(n_626), .B(n_641), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_627), .B(n_634), .Y(n_626) );
OAI21xp5_ASAP7_75t_SL g627 ( .A1(n_628), .A2(n_630), .B(n_631), .Y(n_627) );
INVx2_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_638), .Y(n_634) );
NOR2x1_ASAP7_75t_L g641 ( .A(n_642), .B(n_648), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_646), .Y(n_642) );
BUFx2_ASAP7_75t_L g870 ( .A(n_644), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_652), .Y(n_648) );
BUFx6f_ASAP7_75t_L g740 ( .A(n_651), .Y(n_740) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NOR2x1_ASAP7_75t_L g657 ( .A(n_658), .B(n_664), .Y(n_657) );
NAND4xp25_ASAP7_75t_SL g658 ( .A(n_659), .B(n_660), .C(n_661), .D(n_663), .Y(n_658) );
NAND4xp25_ASAP7_75t_L g664 ( .A(n_665), .B(n_668), .C(n_671), .D(n_672), .Y(n_664) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OA22x2_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B1(n_696), .B2(n_697), .Y(n_677) );
XOR2x2_ASAP7_75t_L g715 ( .A(n_678), .B(n_696), .Y(n_715) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NOR2x1_ASAP7_75t_L g680 ( .A(n_681), .B(n_689), .Y(n_680) );
NAND4xp25_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .C(n_685), .D(n_686), .Y(n_681) );
INVx2_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
NAND4xp25_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .C(n_694), .D(n_695), .Y(n_689) );
INVx2_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OR2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_707), .Y(n_699) );
NAND4xp25_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .C(n_703), .D(n_705), .Y(n_700) );
NAND4xp25_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .C(n_710), .D(n_713), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_896), .B1(n_965), .B2(n_966), .Y(n_716) );
INVxp67_ASAP7_75t_L g965 ( .A(n_717), .Y(n_965) );
AOI22x1_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_719), .B1(n_844), .B2(n_845), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
OA22x2_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_791), .B1(n_792), .B2(n_843), .Y(n_719) );
INVx1_ASAP7_75t_L g843 ( .A(n_720), .Y(n_843) );
AOI22xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_748), .B1(n_789), .B2(n_790), .Y(n_720) );
INVx1_ASAP7_75t_L g789 ( .A(n_721), .Y(n_789) );
NAND3xp33_ASAP7_75t_L g722 ( .A(n_723), .B(n_731), .C(n_741), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_724), .B(n_726), .Y(n_723) );
NOR4xp25_ASAP7_75t_L g745 ( .A(n_724), .B(n_726), .C(n_732), .D(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
BUFx2_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
INVxp67_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
OAI221xp5_ASAP7_75t_SL g732 ( .A1(n_733), .A2(n_734), .B1(n_735), .B2(n_738), .C(n_739), .Y(n_732) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
BUFx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g746 ( .A(n_741), .B(n_747), .Y(n_746) );
AND2x2_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .Y(n_741) );
INVx1_ASAP7_75t_L g790 ( .A(n_748), .Y(n_790) );
OAI22x1_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_769), .B1(n_770), .B2(n_788), .Y(n_748) );
INVx2_ASAP7_75t_L g788 ( .A(n_749), .Y(n_788) );
XNOR2x1_ASAP7_75t_L g749 ( .A(n_750), .B(n_768), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_751), .B(n_758), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_755), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_759), .B(n_765), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_760), .B(n_763), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
OA22x2_ASAP7_75t_L g937 ( .A1(n_769), .A2(n_938), .B1(n_939), .B2(n_960), .Y(n_937) );
INVxp67_ASAP7_75t_L g960 ( .A(n_769), .Y(n_960) );
OA22x2_ASAP7_75t_L g964 ( .A1(n_769), .A2(n_938), .B1(n_939), .B2(n_960), .Y(n_964) );
INVx3_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g787 ( .A(n_771), .Y(n_787) );
NOR2xp67_ASAP7_75t_L g771 ( .A(n_772), .B(n_778), .Y(n_771) );
NAND4xp25_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .C(n_775), .D(n_777), .Y(n_772) );
NAND4xp25_ASAP7_75t_SL g778 ( .A(n_779), .B(n_781), .C(n_783), .D(n_785), .Y(n_778) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_809), .B1(n_841), .B2(n_842), .Y(n_792) );
INVx2_ASAP7_75t_SL g842 ( .A(n_793), .Y(n_842) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
NOR2x1_ASAP7_75t_L g796 ( .A(n_797), .B(n_803), .Y(n_796) );
NAND4xp25_ASAP7_75t_L g797 ( .A(n_798), .B(n_799), .C(n_800), .D(n_801), .Y(n_797) );
NAND4xp25_ASAP7_75t_SL g803 ( .A(n_804), .B(n_805), .C(n_807), .D(n_808), .Y(n_803) );
INVx1_ASAP7_75t_L g841 ( .A(n_809), .Y(n_841) );
OAI22xp33_ASAP7_75t_SL g809 ( .A1(n_810), .A2(n_824), .B1(n_839), .B2(n_840), .Y(n_809) );
INVx1_ASAP7_75t_L g839 ( .A(n_810), .Y(n_839) );
AO22x2_ASAP7_75t_L g848 ( .A1(n_810), .A2(n_839), .B1(n_849), .B2(n_861), .Y(n_848) );
INVx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
NOR2x1_ASAP7_75t_L g813 ( .A(n_814), .B(n_819), .Y(n_813) );
NAND3xp33_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .C(n_818), .Y(n_814) );
NAND4xp25_ASAP7_75t_L g819 ( .A(n_820), .B(n_821), .C(n_822), .D(n_823), .Y(n_819) );
INVx2_ASAP7_75t_L g840 ( .A(n_824), .Y(n_840) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
NOR2xp67_ASAP7_75t_L g826 ( .A(n_827), .B(n_833), .Y(n_826) );
NAND3xp33_ASAP7_75t_L g827 ( .A(n_828), .B(n_831), .C(n_832), .Y(n_827) );
AND2x2_ASAP7_75t_L g828 ( .A(n_829), .B(n_830), .Y(n_828) );
NAND4xp25_ASAP7_75t_L g833 ( .A(n_834), .B(n_835), .C(n_836), .D(n_837), .Y(n_833) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
XOR2x1_ASAP7_75t_SL g845 ( .A(n_846), .B(n_882), .Y(n_845) );
AO22x2_ASAP7_75t_L g846 ( .A1(n_847), .A2(n_848), .B1(n_862), .B2(n_881), .Y(n_846) );
INVx2_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g861 ( .A(n_849), .Y(n_861) );
OR2x2_ASAP7_75t_L g850 ( .A(n_851), .B(n_856), .Y(n_850) );
NAND4xp25_ASAP7_75t_SL g851 ( .A(n_852), .B(n_853), .C(n_854), .D(n_855), .Y(n_851) );
NAND4xp25_ASAP7_75t_SL g856 ( .A(n_857), .B(n_858), .C(n_859), .D(n_860), .Y(n_856) );
INVx1_ASAP7_75t_L g881 ( .A(n_862), .Y(n_881) );
XOR2x2_ASAP7_75t_L g862 ( .A(n_863), .B(n_880), .Y(n_862) );
NOR2x1_ASAP7_75t_L g863 ( .A(n_864), .B(n_872), .Y(n_863) );
NAND4xp25_ASAP7_75t_L g864 ( .A(n_865), .B(n_868), .C(n_869), .D(n_871), .Y(n_864) );
NAND4xp25_ASAP7_75t_L g872 ( .A(n_873), .B(n_874), .C(n_875), .D(n_877), .Y(n_872) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx1_ASAP7_75t_SL g882 ( .A(n_883), .Y(n_882) );
OR2x2_ASAP7_75t_L g884 ( .A(n_885), .B(n_891), .Y(n_884) );
NAND4xp25_ASAP7_75t_L g885 ( .A(n_886), .B(n_887), .C(n_888), .D(n_890), .Y(n_885) );
NAND4xp25_ASAP7_75t_L g891 ( .A(n_892), .B(n_893), .C(n_894), .D(n_895), .Y(n_891) );
OAI21xp5_ASAP7_75t_L g896 ( .A1(n_897), .A2(n_936), .B(n_961), .Y(n_896) );
INVx2_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
AOI21xp5_ASAP7_75t_L g966 ( .A1(n_898), .A2(n_967), .B(n_968), .Y(n_966) );
BUFx3_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx2_ASAP7_75t_L g962 ( .A(n_899), .Y(n_962) );
OA21x2_ASAP7_75t_L g899 ( .A1(n_900), .A2(n_917), .B(n_932), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_900), .B(n_933), .Y(n_932) );
OA22x2_ASAP7_75t_L g939 ( .A1(n_900), .A2(n_940), .B1(n_941), .B2(n_959), .Y(n_939) );
INVx3_ASAP7_75t_SL g959 ( .A(n_900), .Y(n_959) );
XOR2x2_ASAP7_75t_L g900 ( .A(n_901), .B(n_916), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_902), .B(n_909), .Y(n_901) );
NOR2xp33_ASAP7_75t_L g902 ( .A(n_903), .B(n_906), .Y(n_902) );
NAND2xp5_ASAP7_75t_SL g903 ( .A(n_904), .B(n_905), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_907), .B(n_908), .Y(n_906) );
NOR2xp33_ASAP7_75t_L g909 ( .A(n_910), .B(n_913), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_911), .B(n_912), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_914), .B(n_915), .Y(n_913) );
INVxp67_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
INVx2_ASAP7_75t_L g935 ( .A(n_919), .Y(n_935) );
NAND4xp75_ASAP7_75t_L g919 ( .A(n_920), .B(n_925), .C(n_928), .D(n_929), .Y(n_919) );
AND2x2_ASAP7_75t_L g920 ( .A(n_921), .B(n_922), .Y(n_920) );
BUFx2_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
AND2x2_ASAP7_75t_L g925 ( .A(n_926), .B(n_927), .Y(n_925) );
AND2x2_ASAP7_75t_SL g929 ( .A(n_930), .B(n_931), .Y(n_929) );
INVx1_ASAP7_75t_L g967 ( .A(n_936), .Y(n_967) );
INVx2_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
INVx2_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
INVx1_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
XNOR2x2_ASAP7_75t_SL g941 ( .A(n_942), .B(n_943), .Y(n_941) );
OR2x2_ASAP7_75t_L g943 ( .A(n_944), .B(n_951), .Y(n_943) );
NAND4xp25_ASAP7_75t_L g944 ( .A(n_945), .B(n_946), .C(n_948), .D(n_949), .Y(n_944) );
NAND4xp25_ASAP7_75t_L g951 ( .A(n_952), .B(n_954), .C(n_956), .D(n_957), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g961 ( .A(n_962), .B(n_963), .Y(n_961) );
INVx2_ASAP7_75t_L g969 ( .A(n_962), .Y(n_969) );
INVx1_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
NOR2xp33_ASAP7_75t_L g968 ( .A(n_964), .B(n_969), .Y(n_968) );
INVx2_ASAP7_75t_SL g971 ( .A(n_972), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_973), .B(n_976), .Y(n_972) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_973), .B(n_977), .Y(n_1007) );
NOR2xp33_ASAP7_75t_L g973 ( .A(n_974), .B(n_975), .Y(n_973) );
INVx1_ASAP7_75t_L g1016 ( .A(n_975), .Y(n_1016) );
INVx1_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
NAND2xp5_ASAP7_75t_L g978 ( .A(n_979), .B(n_980), .Y(n_978) );
OAI221xp5_ASAP7_75t_L g981 ( .A1(n_982), .A2(n_989), .B1(n_990), .B2(n_1005), .C(n_1008), .Y(n_981) );
OR2x2_ASAP7_75t_L g982 ( .A(n_983), .B(n_987), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
NOR2xp33_ASAP7_75t_L g984 ( .A(n_985), .B(n_986), .Y(n_984) );
INVxp67_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
INVxp67_ASAP7_75t_SL g990 ( .A(n_991), .Y(n_990) );
INVx2_ASAP7_75t_SL g991 ( .A(n_992), .Y(n_991) );
BUFx3_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
HB1xp67_ASAP7_75t_L g1013 ( .A(n_994), .Y(n_1013) );
NOR2xp67_ASAP7_75t_L g994 ( .A(n_995), .B(n_1000), .Y(n_994) );
NAND4xp25_ASAP7_75t_L g995 ( .A(n_996), .B(n_997), .C(n_998), .D(n_999), .Y(n_995) );
NAND4xp25_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1002), .C(n_1003), .D(n_1004), .Y(n_1000) );
INVx1_ASAP7_75t_SL g1005 ( .A(n_1006), .Y(n_1005) );
CKINVDCx6p67_ASAP7_75t_R g1006 ( .A(n_1007), .Y(n_1006) );
CKINVDCx20_ASAP7_75t_R g1012 ( .A(n_1013), .Y(n_1012) );
CKINVDCx20_ASAP7_75t_R g1014 ( .A(n_1015), .Y(n_1014) );
endmodule