module fake_jpeg_24448_n_60 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_60);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_60;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

INVx8_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_0),
.B(n_6),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_2),
.B(n_8),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx8_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_18),
.B(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_0),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_20),
.B(n_12),
.Y(n_31)
);

AOI21xp33_ASAP7_75t_L g21 ( 
.A1(n_11),
.A2(n_1),
.B(n_2),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_13),
.C(n_17),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_1),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_24),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_23),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_31),
.Y(n_34)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_28),
.B(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_38),
.C(n_39),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_30),
.A2(n_9),
.B1(n_15),
.B2(n_12),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_9),
.B1(n_13),
.B2(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_43),
.Y(n_50)
);

MAJx2_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_16),
.C(n_14),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_45),
.C(n_16),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_16),
.B(n_14),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_46),
.B(n_49),
.Y(n_53)
);

NAND3xp33_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_33),
.C(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_42),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_9),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_16),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_47),
.Y(n_54)
);

A2O1A1O1Ixp25_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_53),
.B(n_51),
.C(n_6),
.D(n_5),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_14),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_57),
.B(n_3),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_58),
.Y(n_59)
);

NAND4xp25_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_55),
.C(n_5),
.D(n_14),
.Y(n_60)
);


endmodule