module fake_jpeg_9651_n_253 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_253);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_253;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_38),
.Y(n_44)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_21),
.Y(n_37)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_42),
.Y(n_46)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_20),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_49),
.Y(n_87)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_51),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_54),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_20),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_23),
.Y(n_67)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_25),
.B1(n_31),
.B2(n_17),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_64),
.B1(n_15),
.B2(n_28),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_25),
.B1(n_30),
.B2(n_29),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_56),
.A2(n_58),
.B1(n_17),
.B2(n_19),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_32),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_57),
.B(n_63),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_34),
.A2(n_30),
.B1(n_29),
.B2(n_16),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_36),
.A2(n_26),
.B1(n_16),
.B2(n_19),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_22),
.B1(n_27),
.B2(n_21),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_32),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_34),
.A2(n_31),
.B1(n_17),
.B2(n_26),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_31),
.Y(n_66)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_74),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_66),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_70),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_0),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_71),
.A2(n_83),
.B(n_28),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_75),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_37),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_34),
.B1(n_33),
.B2(n_23),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_76),
.A2(n_81),
.B1(n_50),
.B2(n_52),
.Y(n_95)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_46),
.A2(n_15),
.B(n_21),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_58),
.C(n_63),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_78),
.Y(n_90)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_46),
.A2(n_27),
.B1(n_23),
.B2(n_40),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_60),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_47),
.Y(n_92)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_96),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_105),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_85),
.B1(n_75),
.B2(n_50),
.Y(n_120)
);

INVx6_ASAP7_75t_SL g96 ( 
.A(n_68),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_102),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_51),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_76),
.B(n_77),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_43),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_101),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_43),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_80),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_86),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_57),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_107),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_70),
.Y(n_107)
);

BUFx24_ASAP7_75t_SL g108 ( 
.A(n_69),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_109),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_86),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_74),
.C(n_67),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_116),
.C(n_119),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_73),
.C(n_80),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_117),
.A2(n_126),
.B(n_32),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_72),
.C(n_81),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_120),
.A2(n_91),
.B1(n_90),
.B2(n_110),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_96),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_122),
.Y(n_139)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_91),
.A2(n_68),
.B1(n_62),
.B2(n_72),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_124),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_88),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_54),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_129),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_65),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_131),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_102),
.B(n_78),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_90),
.A2(n_62),
.B1(n_79),
.B2(n_65),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_133),
.A2(n_91),
.B1(n_95),
.B2(n_79),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_105),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_136),
.B(n_138),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_118),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_137),
.B(n_142),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_107),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_101),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_153),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_141),
.A2(n_148),
.B(n_151),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_125),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_144),
.A2(n_131),
.B1(n_135),
.B2(n_134),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_133),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_145),
.B(n_146),
.Y(n_165)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_120),
.A2(n_106),
.B1(n_109),
.B2(n_104),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_147),
.A2(n_113),
.B1(n_119),
.B2(n_116),
.Y(n_168)
);

NAND2x1_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_98),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_94),
.B(n_97),
.Y(n_151)
);

OAI211xp5_ASAP7_75t_SL g152 ( 
.A1(n_112),
.A2(n_93),
.B(n_35),
.C(n_40),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_65),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_93),
.C(n_61),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_154),
.A2(n_134),
.B(n_149),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_48),
.Y(n_155)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_115),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_114),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_139),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_166),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_159),
.A2(n_171),
.B1(n_173),
.B2(n_177),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_122),
.Y(n_161)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_154),
.B(n_152),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_147),
.B(n_126),
.Y(n_166)
);

NOR2x1_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_123),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_167),
.B(n_169),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_168),
.A2(n_138),
.B1(n_140),
.B2(n_128),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_135),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_143),
.A2(n_114),
.B1(n_113),
.B2(n_121),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_172),
.A2(n_174),
.B1(n_149),
.B2(n_148),
.Y(n_180)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_151),
.A2(n_121),
.B1(n_129),
.B2(n_68),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_129),
.Y(n_176)
);

AOI21xp33_ASAP7_75t_L g192 ( 
.A1(n_176),
.A2(n_28),
.B(n_35),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_136),
.C(n_150),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_183),
.C(n_186),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_180),
.A2(n_181),
.B(n_189),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_175),
.C(n_150),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_159),
.Y(n_203)
);

A2O1A1O1Ixp25_ASAP7_75t_L g185 ( 
.A1(n_167),
.A2(n_61),
.B(n_32),
.C(n_35),
.D(n_60),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_193),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_32),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_157),
.C(n_163),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_161),
.C(n_162),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_174),
.B(n_173),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_28),
.B(n_60),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_191),
.A2(n_158),
.B(n_172),
.Y(n_200)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_192),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_165),
.A2(n_103),
.B1(n_48),
.B2(n_0),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_194),
.A2(n_103),
.B1(n_177),
.B2(n_4),
.Y(n_206)
);

BUFx12_ASAP7_75t_L g198 ( 
.A(n_190),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_204),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_203),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_166),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_205),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_162),
.C(n_164),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_206),
.A2(n_185),
.B1(n_4),
.B2(n_5),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_178),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_207),
.A2(n_209),
.B(n_210),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_28),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_1),
.Y(n_219)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_195),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_191),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_196),
.B(n_189),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_196),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_214),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_209),
.B(n_180),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_200),
.A2(n_188),
.B1(n_181),
.B2(n_184),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_216),
.A2(n_221),
.B1(n_206),
.B2(n_197),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_205),
.B(n_186),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_218),
.B(n_219),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_220),
.B(n_2),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_210),
.A2(n_183),
.B1(n_4),
.B2(n_5),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_222),
.A2(n_199),
.B(n_197),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_223),
.A2(n_225),
.B(n_2),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_204),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_226),
.B(n_228),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_198),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_217),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_231),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_201),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_237),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_227),
.A2(n_212),
.B(n_215),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_235),
.C(n_236),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_224),
.A2(n_201),
.B(n_221),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_228),
.A2(n_203),
.B1(n_5),
.B2(n_6),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_238),
.B(n_226),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_240),
.B(n_243),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_231),
.Y(n_242)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_242),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_2),
.Y(n_243)
);

AOI31xp67_ASAP7_75t_SL g245 ( 
.A1(n_239),
.A2(n_7),
.A3(n_8),
.B(n_9),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_245),
.A2(n_247),
.B(n_11),
.Y(n_249)
);

O2A1O1Ixp33_ASAP7_75t_SL g247 ( 
.A1(n_241),
.A2(n_7),
.B(n_9),
.C(n_10),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_10),
.C(n_11),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_248),
.A2(n_12),
.B(n_13),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_SL g250 ( 
.A1(n_249),
.A2(n_244),
.B(n_13),
.C(n_14),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_250),
.A2(n_251),
.B1(n_12),
.B2(n_13),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_12),
.C(n_14),
.Y(n_253)
);


endmodule