module fake_jpeg_12276_n_119 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_119);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_119;

wire n_117;
wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_12),
.B(n_1),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_30),
.B(n_31),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_12),
.B(n_5),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_10),
.A2(n_5),
.B1(n_2),
.B2(n_3),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_32),
.A2(n_42),
.B1(n_50),
.B2(n_54),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_2),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_33),
.B(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_10),
.B(n_3),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_41),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_3),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_34),
.C(n_52),
.Y(n_62)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_15),
.A2(n_21),
.B1(n_23),
.B2(n_22),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_11),
.A2(n_27),
.B1(n_26),
.B2(n_20),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_47),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_16),
.A2(n_21),
.B(n_23),
.C(n_22),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_19),
.B(n_20),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_27),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_26),
.A2(n_27),
.B1(n_14),
.B2(n_13),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_52),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_28),
.B(n_15),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_28),
.B(n_14),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_49),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_10),
.A2(n_18),
.B1(n_25),
.B2(n_26),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_59),
.B(n_64),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_62),
.B(n_76),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_37),
.Y(n_67)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_46),
.B(n_40),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_39),
.B(n_38),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_90),
.C(n_61),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_66),
.B1(n_60),
.B2(n_71),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_79),
.B(n_91),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_60),
.A2(n_73),
.B1(n_68),
.B2(n_66),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_72),
.B(n_55),
.Y(n_98)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_57),
.B(n_58),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_83),
.A2(n_72),
.B(n_61),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_87),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_57),
.A2(n_62),
.B1(n_69),
.B2(n_74),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_57),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_88),
.B(n_72),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_63),
.B(n_68),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_55),
.A2(n_70),
.B1(n_66),
.B2(n_60),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_93),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_85),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_96),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_98),
.A2(n_88),
.B1(n_83),
.B2(n_78),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_101),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_95),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_107),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_105),
.A2(n_100),
.B1(n_101),
.B2(n_87),
.Y(n_112)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_108),
.B(n_100),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_99),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_111),
.Y(n_114)
);

A2O1A1O1Ixp25_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_104),
.B(n_100),
.C(n_106),
.D(n_108),
.Y(n_113)
);

NOR3xp33_ASAP7_75t_SL g115 ( 
.A(n_113),
.B(n_82),
.C(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_116),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_117),
.B(n_114),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_109),
.Y(n_119)
);


endmodule