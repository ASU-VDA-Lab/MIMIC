module fake_jpeg_15592_n_327 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_327);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx5p33_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_39),
.B(n_40),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_41),
.B(n_42),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_21),
.B(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_21),
.B(n_8),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_20),
.A2(n_8),
.B1(n_2),
.B2(n_3),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_52),
.A2(n_13),
.B1(n_31),
.B2(n_33),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_8),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_65),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_57),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_60),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_22),
.B(n_1),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_61),
.B(n_2),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_64),
.Y(n_90)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_22),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_20),
.B(n_1),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_33),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_70),
.B(n_99),
.Y(n_153)
);

BUFx4f_ASAP7_75t_SL g72 ( 
.A(n_63),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_72),
.Y(n_146)
);

AO22x2_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_17),
.B1(n_18),
.B2(n_15),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_74),
.A2(n_76),
.B1(n_96),
.B2(n_106),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_32),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_75),
.B(n_77),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_19),
.B1(n_20),
.B2(n_32),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_25),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_79),
.B(n_84),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_115),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_42),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_51),
.A2(n_19),
.B1(n_38),
.B2(n_55),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_86),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_130)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_65),
.B(n_31),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_87),
.A2(n_17),
.B(n_26),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_41),
.B(n_27),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_89),
.B(n_95),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_30),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_60),
.A2(n_19),
.B1(n_13),
.B2(n_30),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_67),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

CKINVDCx6p67_ASAP7_75t_R g102 ( 
.A(n_57),
.Y(n_102)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_57),
.A2(n_13),
.B1(n_15),
.B2(n_3),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_44),
.A2(n_29),
.B1(n_27),
.B2(n_15),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_44),
.A2(n_29),
.B1(n_34),
.B2(n_5),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_46),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_62),
.B(n_24),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_24),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_111),
.B(n_6),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_46),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_112),
.A2(n_103),
.B1(n_98),
.B2(n_93),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_114),
.Y(n_147)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_50),
.A2(n_17),
.B1(n_26),
.B2(n_24),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_116),
.Y(n_185)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_53),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_119),
.B(n_133),
.Y(n_162)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_121),
.Y(n_174)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_131),
.Y(n_166)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_124),
.A2(n_149),
.B1(n_128),
.B2(n_117),
.Y(n_196)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_125),
.Y(n_190)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_126),
.Y(n_179)
);

AO22x2_ASAP7_75t_L g127 ( 
.A1(n_74),
.A2(n_115),
.B1(n_106),
.B2(n_109),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_127),
.A2(n_107),
.B1(n_105),
.B2(n_102),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_90),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_141),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_132),
.Y(n_167)
);

A2O1A1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_75),
.B(n_80),
.C(n_83),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_50),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_71),
.Y(n_177)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_135),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_17),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_136),
.B(n_137),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_88),
.B(n_17),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_L g139 ( 
.A1(n_74),
.A2(n_53),
.B(n_7),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_139),
.A2(n_102),
.B(n_81),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

BUFx16f_ASAP7_75t_L g142 ( 
.A(n_72),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_144),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_82),
.B(n_26),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_145),
.B(n_151),
.Y(n_164)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_148),
.B(n_160),
.Y(n_183)
);

INVx11_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_73),
.B(n_66),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_69),
.B(n_66),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_152),
.B(n_156),
.Y(n_191)
);

AND2x4_ASAP7_75t_L g154 ( 
.A(n_74),
.B(n_66),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_81),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_93),
.B(n_101),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_159),
.B1(n_130),
.B2(n_86),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_101),
.B(n_115),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_158),
.B(n_154),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_112),
.A2(n_103),
.B1(n_98),
.B2(n_108),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_101),
.Y(n_160)
);

BUFx8_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_163),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_165),
.A2(n_194),
.B1(n_121),
.B2(n_120),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_168),
.A2(n_176),
.B(n_180),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_72),
.C(n_71),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_198),
.C(n_138),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_172),
.A2(n_189),
.B1(n_192),
.B2(n_195),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_119),
.B(n_104),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_182),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_104),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_178),
.B(n_184),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_134),
.B(n_114),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_146),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_146),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_143),
.B(n_155),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_188),
.B(n_193),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_127),
.A2(n_118),
.B1(n_148),
.B2(n_154),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_127),
.A2(n_154),
.B1(n_118),
.B2(n_150),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_127),
.B(n_122),
.Y(n_194)
);

OA21x2_ASAP7_75t_L g195 ( 
.A1(n_127),
.A2(n_123),
.B(n_118),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_196),
.Y(n_211)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_120),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_197),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_150),
.B(n_133),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_135),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_200),
.A2(n_212),
.B(n_168),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_143),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_202),
.B(n_215),
.C(n_230),
.Y(n_249)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_203),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_L g204 ( 
.A1(n_162),
.A2(n_138),
.B(n_142),
.Y(n_204)
);

AOI221xp5_ASAP7_75t_L g241 ( 
.A1(n_204),
.A2(n_220),
.B1(n_180),
.B2(n_166),
.C(n_161),
.Y(n_241)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_205),
.Y(n_231)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_207),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_147),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_208),
.B(n_209),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_147),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_140),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_194),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_218),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_166),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_162),
.B(n_128),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_217),
.A2(n_169),
.B1(n_174),
.B2(n_171),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_126),
.Y(n_218)
);

AND2x6_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_144),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_173),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_221),
.B(n_223),
.Y(n_239)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_179),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_124),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_229),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_185),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_225),
.Y(n_236)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_169),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_226),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_164),
.B(n_141),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_227),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_181),
.B(n_149),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_181),
.B(n_116),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_170),
.B(n_116),
.C(n_140),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_206),
.B(n_195),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_215),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_210),
.A2(n_172),
.B1(n_168),
.B2(n_166),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_235),
.A2(n_256),
.B1(n_230),
.B2(n_218),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_237),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_241),
.A2(n_246),
.B(n_247),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_257),
.C(n_223),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_206),
.A2(n_183),
.B(n_176),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_200),
.A2(n_176),
.B(n_190),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_207),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_250),
.B(n_205),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_200),
.A2(n_190),
.B(n_191),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_213),
.A2(n_167),
.B(n_175),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_201),
.B(n_174),
.Y(n_254)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_254),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_212),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_199),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_224),
.A2(n_171),
.B1(n_116),
.B2(n_185),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_202),
.B(n_163),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_233),
.A2(n_211),
.B1(n_212),
.B2(n_217),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_258),
.A2(n_255),
.B1(n_247),
.B2(n_252),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_259),
.A2(n_274),
.B1(n_244),
.B2(n_243),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_260),
.B(n_269),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_201),
.Y(n_261)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_214),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_249),
.C(n_245),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_236),
.Y(n_263)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_263),
.Y(n_287)
);

AOI322xp5_ASAP7_75t_SL g264 ( 
.A1(n_234),
.A2(n_219),
.A3(n_222),
.B1(n_220),
.B2(n_216),
.C1(n_163),
.C2(n_226),
.Y(n_264)
);

AOI322xp5_ASAP7_75t_SL g283 ( 
.A1(n_264),
.A2(n_277),
.A3(n_253),
.B1(n_238),
.B2(n_251),
.C1(n_235),
.C2(n_244),
.Y(n_283)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_265),
.A2(n_266),
.B(n_267),
.Y(n_280)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_231),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_199),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_270),
.A2(n_271),
.B(n_273),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_231),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_232),
.B(n_216),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_239),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_240),
.C(n_256),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_234),
.B(n_236),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_249),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_281),
.C(n_285),
.Y(n_300)
);

NAND3xp33_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_268),
.C(n_275),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_246),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_240),
.C(n_237),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_293),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_290),
.A2(n_278),
.B1(n_261),
.B2(n_271),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_263),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_292),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_289),
.A2(n_258),
.B(n_268),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_294),
.A2(n_303),
.B1(n_304),
.B2(n_298),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_290),
.B(n_274),
.Y(n_296)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_296),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_299),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_280),
.A2(n_278),
.B(n_269),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_298),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_265),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_288),
.Y(n_306)
);

O2A1O1Ixp33_ASAP7_75t_SL g303 ( 
.A1(n_284),
.A2(n_242),
.B(n_266),
.C(n_267),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_289),
.A2(n_225),
.B1(n_293),
.B2(n_287),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_291),
.B(n_285),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_305),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_300),
.C(n_301),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_302),
.A2(n_282),
.B1(n_292),
.B2(n_288),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_307),
.A2(n_308),
.B1(n_314),
.B2(n_312),
.Y(n_317)
);

OAI21xp33_ASAP7_75t_L g308 ( 
.A1(n_294),
.A2(n_279),
.B(n_281),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_313),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_303),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_300),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_317),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_319),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_297),
.Y(n_319)
);

FAx1_ASAP7_75t_SL g322 ( 
.A(n_315),
.B(n_310),
.CI(n_306),
.CON(n_322),
.SN(n_322)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_322),
.B(n_318),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_323),
.B(n_324),
.C(n_320),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_321),
.A2(n_308),
.B(n_307),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_322),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_322),
.Y(n_327)
);


endmodule