module fake_jpeg_13584_n_142 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_142);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx6_ASAP7_75t_SL g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_37),
.Y(n_38)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_52),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_23),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_16),
.Y(n_56)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx2_ASAP7_75t_SL g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_13),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_49),
.B(n_50),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_13),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_30),
.A2(n_20),
.B1(n_27),
.B2(n_15),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_31),
.B1(n_29),
.B2(n_20),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_33),
.B1(n_36),
.B2(n_34),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_14),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_54),
.B(n_58),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_34),
.B1(n_30),
.B2(n_27),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_55),
.A2(n_69),
.B1(n_18),
.B2(n_21),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_24),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_38),
.Y(n_58)
);

A2O1A1O1Ixp25_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_14),
.B(n_25),
.C(n_24),
.D(n_23),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_41),
.B(n_47),
.C(n_22),
.Y(n_75)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_39),
.B(n_25),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_19),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_52),
.Y(n_72)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

OAI22x1_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_41),
.B1(n_21),
.B2(n_17),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_42),
.A2(n_20),
.B1(n_48),
.B2(n_16),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_48),
.B1(n_42),
.B2(n_46),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_71),
.A2(n_78),
.B1(n_79),
.B2(n_82),
.Y(n_93)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

NAND3xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_75),
.C(n_81),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_55),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_57),
.A2(n_42),
.B1(n_46),
.B2(n_44),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_68),
.A2(n_20),
.B1(n_26),
.B2(n_22),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_83),
.A2(n_61),
.B1(n_67),
.B2(n_53),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_26),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_63),
.C(n_53),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_90),
.C(n_45),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_75),
.B(n_65),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_92),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_66),
.Y(n_90)
);

AO21x1_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_53),
.B(n_62),
.Y(n_91)
);

NOR3xp33_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_98),
.C(n_77),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_94),
.B(n_96),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_80),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_62),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_97),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_59),
.B(n_17),
.Y(n_98)
);

OAI22x1_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_60),
.B1(n_69),
.B2(n_17),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_21),
.Y(n_111)
);

AOI322xp5_ASAP7_75t_SL g102 ( 
.A1(n_89),
.A2(n_73),
.A3(n_74),
.B1(n_78),
.B2(n_11),
.C1(n_71),
.C2(n_19),
.Y(n_102)
);

OAI322xp33_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_108),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_9),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_104),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_95),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_109),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_82),
.B1(n_79),
.B2(n_45),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_106),
.A2(n_93),
.B1(n_2),
.B2(n_3),
.Y(n_117)
);

AOI322xp5_ASAP7_75t_SL g108 ( 
.A1(n_87),
.A2(n_21),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_26),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_90),
.C(n_94),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_111),
.A2(n_88),
.B1(n_99),
.B2(n_92),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_116),
.C(n_118),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_119),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_98),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_1),
.C(n_4),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_6),
.B(n_7),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_7),
.Y(n_126)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_122),
.Y(n_128)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_126),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_118),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_130),
.B(n_132),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_105),
.Y(n_131)
);

OAI21x1_ASAP7_75t_L g134 ( 
.A1(n_131),
.A2(n_111),
.B(n_106),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_113),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_131),
.A2(n_125),
.B1(n_100),
.B2(n_123),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_133),
.B(n_136),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_134),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_128),
.A2(n_116),
.B(n_101),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_129),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_138),
.A2(n_101),
.B(n_139),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_137),
.A2(n_101),
.B(n_9),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_140),
.B(n_141),
.Y(n_142)
);


endmodule