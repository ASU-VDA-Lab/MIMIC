module fake_jpeg_29622_n_117 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_117);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_117;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_22),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

AND2x2_ASAP7_75t_SL g44 ( 
.A(n_30),
.B(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_43),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_53),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_48),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_58),
.B(n_1),
.Y(n_67)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_59),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_15),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_2),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_19),
.B1(n_35),
.B2(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_62),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_46),
.C(n_50),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_59),
.B(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_64),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_68),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_55),
.B(n_39),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_3),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_71),
.B(n_3),
.Y(n_83)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_53),
.B1(n_41),
.B2(n_49),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_73),
.A2(n_75),
.B1(n_81),
.B2(n_74),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_41),
.B1(n_49),
.B2(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_70),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_84),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_45),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_80),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_40),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_42),
.B1(n_21),
.B2(n_24),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_85),
.B1(n_5),
.B2(n_6),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_4),
.Y(n_90)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_67),
.A2(n_42),
.B1(n_14),
.B2(n_25),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_86),
.B(n_27),
.Y(n_96)
);

NOR3xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_4),
.C(n_5),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_90),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_94),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_28),
.B1(n_32),
.B2(n_13),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_7),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_98),
.B(n_9),
.Y(n_104)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_72),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_99),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_8),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_76),
.B(n_8),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_105),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_26),
.C(n_31),
.Y(n_107)
);

A2O1A1O1Ixp25_ASAP7_75t_L g110 ( 
.A1(n_107),
.A2(n_95),
.B(n_88),
.C(n_94),
.D(n_11),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_103),
.Y(n_109)
);

BUFx24_ASAP7_75t_SL g112 ( 
.A(n_109),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_107),
.C(n_101),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_108),
.Y(n_113)
);

OAI21x1_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_112),
.B(n_102),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_114),
.Y(n_115)
);

AOI322xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_106),
.A3(n_92),
.B1(n_100),
.B2(n_37),
.C1(n_91),
.C2(n_11),
.Y(n_116)
);

NOR2xp67_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_9),
.Y(n_117)
);


endmodule