module fake_jpeg_18273_n_125 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_125);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx10_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_25),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx11_ASAP7_75t_SL g50 ( 
.A(n_29),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_13),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_24),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_60),
.Y(n_75)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_0),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_63),
.Y(n_65)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_1),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_64),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_59),
.A2(n_44),
.B1(n_46),
.B2(n_36),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_67),
.A2(n_69),
.B1(n_41),
.B2(n_75),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_46),
.B1(n_50),
.B2(n_57),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_74),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_35),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_35),
.Y(n_87)
);

INVx5_ASAP7_75t_SL g74 ( 
.A(n_59),
.Y(n_74)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_77),
.Y(n_93)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_72),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_39),
.Y(n_80)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_55),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_83),
.B(n_84),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_54),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_78),
.B1(n_81),
.B2(n_86),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_51),
.B(n_43),
.Y(n_86)
);

NOR2x1_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_3),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_87),
.B(n_56),
.Y(n_92)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_2),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_79),
.A2(n_49),
.B1(n_40),
.B2(n_52),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_92),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_37),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_91),
.B(n_102),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_94),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_88),
.A2(n_48),
.B1(n_22),
.B2(n_23),
.Y(n_95)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_88),
.B(n_1),
.Y(n_96)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_5),
.Y(n_101)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_8),
.C(n_14),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_105),
.B(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_98),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_113),
.C(n_114),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_106),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_93),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_116),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_100),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_108),
.B1(n_104),
.B2(n_110),
.Y(n_119)
);

FAx1_ASAP7_75t_SL g120 ( 
.A(n_119),
.B(n_115),
.CI(n_89),
.CON(n_120),
.SN(n_120)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_103),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_121),
.A2(n_109),
.B(n_107),
.Y(n_122)
);

AO221x1_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.C(n_19),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_20),
.B(n_21),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);


endmodule