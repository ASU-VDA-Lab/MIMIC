module real_aes_8200_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_754;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g541 ( .A1(n_0), .A2(n_188), .B(n_542), .C(n_545), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_1), .B(n_530), .Y(n_546) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_2), .B(n_111), .C(n_112), .Y(n_110) );
INVx1_ASAP7_75t_L g433 ( .A(n_2), .Y(n_433) );
OAI22xp5_ASAP7_75t_SL g750 ( .A1(n_3), .A2(n_751), .B1(n_754), .B2(n_755), .Y(n_750) );
INVx1_ASAP7_75t_L g755 ( .A(n_3), .Y(n_755) );
INVx1_ASAP7_75t_L g206 ( .A(n_4), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_5), .B(n_177), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_6), .A2(n_445), .B(n_524), .Y(n_523) );
AO21x2_ASAP7_75t_L g491 ( .A1(n_7), .A2(n_153), .B(n_492), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g187 ( .A1(n_8), .A2(n_36), .B1(n_133), .B2(n_142), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_9), .B(n_153), .Y(n_217) );
AND2x6_ASAP7_75t_L g151 ( .A(n_10), .B(n_152), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_11), .A2(n_151), .B(n_448), .C(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g108 ( .A(n_12), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_12), .B(n_37), .Y(n_434) );
INVx1_ASAP7_75t_L g149 ( .A(n_13), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_14), .B(n_140), .Y(n_160) );
INVx1_ASAP7_75t_L g198 ( .A(n_15), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_16), .B(n_177), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_17), .B(n_154), .Y(n_222) );
AO32x2_ASAP7_75t_L g185 ( .A1(n_18), .A2(n_150), .A3(n_153), .B1(n_186), .B2(n_190), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_19), .B(n_142), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_20), .B(n_154), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g189 ( .A1(n_21), .A2(n_52), .B1(n_133), .B2(n_142), .Y(n_189) );
AOI22xp33_ASAP7_75t_SL g139 ( .A1(n_22), .A2(n_81), .B1(n_140), .B2(n_142), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_23), .B(n_142), .Y(n_179) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_24), .A2(n_150), .B(n_448), .C(n_450), .Y(n_447) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_25), .A2(n_150), .B(n_448), .C(n_495), .Y(n_494) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_26), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_27), .B(n_145), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_28), .A2(n_445), .B(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_29), .B(n_145), .Y(n_183) );
INVx2_ASAP7_75t_L g135 ( .A(n_30), .Y(n_135) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_31), .A2(n_469), .B(n_478), .C(n_480), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_32), .B(n_142), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_33), .B(n_145), .Y(n_167) );
OAI22xp5_ASAP7_75t_L g117 ( .A1(n_34), .A2(n_73), .B1(n_118), .B2(n_119), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_34), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_35), .B(n_162), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_37), .B(n_108), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_38), .B(n_444), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_39), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_40), .B(n_177), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_41), .B(n_445), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_42), .A2(n_469), .B(n_478), .C(n_515), .Y(n_514) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_43), .A2(n_123), .B1(n_427), .B2(n_428), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_43), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_43), .A2(n_79), .B1(n_427), .B2(n_753), .Y(n_752) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_44), .B(n_142), .Y(n_212) );
INVx1_ASAP7_75t_L g543 ( .A(n_45), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g132 ( .A1(n_46), .A2(n_89), .B1(n_133), .B2(n_136), .Y(n_132) );
INVx1_ASAP7_75t_L g516 ( .A(n_47), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_48), .B(n_142), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_49), .B(n_142), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_50), .B(n_445), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_51), .B(n_204), .Y(n_216) );
AOI22xp33_ASAP7_75t_SL g226 ( .A1(n_53), .A2(n_58), .B1(n_140), .B2(n_142), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_54), .Y(n_457) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_55), .B(n_142), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_56), .B(n_142), .Y(n_241) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_57), .Y(n_759) );
INVx1_ASAP7_75t_L g152 ( .A(n_59), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_60), .B(n_445), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_61), .B(n_530), .Y(n_529) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_62), .A2(n_201), .B(n_204), .C(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_63), .B(n_142), .Y(n_207) );
INVx1_ASAP7_75t_L g148 ( .A(n_64), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_65), .Y(n_746) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_66), .B(n_177), .Y(n_482) );
AO32x2_ASAP7_75t_L g130 ( .A1(n_67), .A2(n_131), .A3(n_144), .B1(n_150), .B2(n_153), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_68), .B(n_143), .Y(n_506) );
INVx1_ASAP7_75t_L g240 ( .A(n_69), .Y(n_240) );
INVx1_ASAP7_75t_L g175 ( .A(n_70), .Y(n_175) );
CKINVDCx16_ASAP7_75t_R g540 ( .A(n_71), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_72), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g119 ( .A(n_73), .Y(n_119) );
A2O1A1Ixp33_ASAP7_75t_L g464 ( .A1(n_74), .A2(n_448), .B(n_465), .C(n_469), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_75), .B(n_140), .Y(n_176) );
CKINVDCx16_ASAP7_75t_R g525 ( .A(n_76), .Y(n_525) );
INVx1_ASAP7_75t_L g114 ( .A(n_77), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_78), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_79), .Y(n_753) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_80), .B(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_82), .B(n_133), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_83), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_84), .B(n_140), .Y(n_180) );
INVx2_ASAP7_75t_L g146 ( .A(n_85), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_86), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_87), .B(n_137), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_88), .B(n_140), .Y(n_213) );
INVx2_ASAP7_75t_L g111 ( .A(n_90), .Y(n_111) );
OR2x2_ASAP7_75t_L g431 ( .A(n_90), .B(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g749 ( .A(n_90), .B(n_743), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_91), .A2(n_101), .B1(n_140), .B2(n_141), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_92), .B(n_445), .Y(n_476) );
INVx1_ASAP7_75t_L g481 ( .A(n_93), .Y(n_481) );
INVxp67_ASAP7_75t_L g528 ( .A(n_94), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_95), .A2(n_103), .B1(n_115), .B2(n_762), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_96), .B(n_140), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_97), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g466 ( .A(n_98), .Y(n_466) );
INVx1_ASAP7_75t_L g502 ( .A(n_99), .Y(n_502) );
AND2x2_ASAP7_75t_L g518 ( .A(n_100), .B(n_145), .Y(n_518) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g762 ( .A(n_105), .Y(n_762) );
AND2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_109), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g730 ( .A(n_111), .B(n_432), .Y(n_730) );
NOR2x2_ASAP7_75t_L g742 ( .A(n_111), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
AO221x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_744), .B1(n_747), .B2(n_756), .C(n_758), .Y(n_115) );
OAI222xp33_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_120), .B1(n_731), .B2(n_732), .C1(n_738), .C2(n_739), .Y(n_116) );
INVx1_ASAP7_75t_L g731 ( .A(n_117), .Y(n_731) );
INVxp67_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_429), .B1(n_435), .B2(n_728), .Y(n_121) );
INVx1_ASAP7_75t_L g734 ( .A(n_122), .Y(n_734) );
INVx2_ASAP7_75t_L g428 ( .A(n_123), .Y(n_428) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
XOR2x2_ASAP7_75t_L g751 ( .A(n_124), .B(n_752), .Y(n_751) );
AND3x1_ASAP7_75t_L g124 ( .A(n_125), .B(n_347), .C(n_395), .Y(n_124) );
NOR4xp25_ASAP7_75t_L g125 ( .A(n_126), .B(n_275), .C(n_320), .D(n_334), .Y(n_125) );
OAI311xp33_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_191), .A3(n_218), .B1(n_228), .C1(n_243), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_155), .Y(n_127) );
OAI21xp33_ASAP7_75t_L g228 ( .A1(n_128), .A2(n_229), .B(n_231), .Y(n_228) );
AND2x2_ASAP7_75t_L g336 ( .A(n_128), .B(n_263), .Y(n_336) );
AND2x2_ASAP7_75t_L g393 ( .A(n_128), .B(n_279), .Y(n_393) );
BUFx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g286 ( .A(n_129), .B(n_184), .Y(n_286) );
AND2x2_ASAP7_75t_L g343 ( .A(n_129), .B(n_291), .Y(n_343) );
INVx1_ASAP7_75t_L g384 ( .A(n_129), .Y(n_384) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_130), .Y(n_252) );
AND2x2_ASAP7_75t_L g293 ( .A(n_130), .B(n_184), .Y(n_293) );
AND2x2_ASAP7_75t_L g297 ( .A(n_130), .B(n_185), .Y(n_297) );
INVx1_ASAP7_75t_L g309 ( .A(n_130), .Y(n_309) );
OAI22xp5_ASAP7_75t_SL g131 ( .A1(n_132), .A2(n_137), .B1(n_139), .B2(n_143), .Y(n_131) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
BUFx3_ASAP7_75t_L g136 ( .A(n_134), .Y(n_136) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_134), .Y(n_142) );
AND2x6_ASAP7_75t_L g448 ( .A(n_134), .B(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g141 ( .A(n_135), .Y(n_141) );
INVx1_ASAP7_75t_L g205 ( .A(n_135), .Y(n_205) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_136), .Y(n_483) );
INVx2_ASAP7_75t_L g545 ( .A(n_136), .Y(n_545) );
INVx2_ASAP7_75t_L g166 ( .A(n_137), .Y(n_166) );
OAI22xp5_ASAP7_75t_L g186 ( .A1(n_137), .A2(n_187), .B1(n_188), .B2(n_189), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g224 ( .A1(n_137), .A2(n_188), .B1(n_225), .B2(n_226), .Y(n_224) );
INVx4_ASAP7_75t_L g544 ( .A(n_137), .Y(n_544) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx3_ASAP7_75t_L g143 ( .A(n_138), .Y(n_143) );
INVx1_ASAP7_75t_L g162 ( .A(n_138), .Y(n_162) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_138), .Y(n_182) );
AND2x2_ASAP7_75t_L g446 ( .A(n_138), .B(n_205), .Y(n_446) );
INVx1_ASAP7_75t_L g449 ( .A(n_138), .Y(n_449) );
INVx2_ASAP7_75t_L g199 ( .A(n_140), .Y(n_199) );
INVx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx3_ASAP7_75t_L g174 ( .A(n_142), .Y(n_174) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_142), .Y(n_468) );
INVx5_ASAP7_75t_L g177 ( .A(n_143), .Y(n_177) );
INVx1_ASAP7_75t_L g455 ( .A(n_144), .Y(n_455) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_145), .A2(n_157), .B(n_167), .Y(n_156) );
OA21x2_ASAP7_75t_L g171 ( .A1(n_145), .A2(n_172), .B(n_183), .Y(n_171) );
INVx1_ASAP7_75t_L g458 ( .A(n_145), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_145), .A2(n_476), .B(n_477), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_145), .A2(n_513), .B(n_514), .Y(n_512) );
AND2x2_ASAP7_75t_SL g145 ( .A(n_146), .B(n_147), .Y(n_145) );
AND2x2_ASAP7_75t_L g154 ( .A(n_146), .B(n_147), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
NAND3xp33_ASAP7_75t_L g223 ( .A(n_150), .B(n_224), .C(n_227), .Y(n_223) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_150), .A2(n_236), .B(n_239), .Y(n_235) );
BUFx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
OAI21xp5_ASAP7_75t_L g157 ( .A1(n_151), .A2(n_158), .B(n_163), .Y(n_157) );
OAI21xp5_ASAP7_75t_L g172 ( .A1(n_151), .A2(n_173), .B(n_178), .Y(n_172) );
OAI21xp5_ASAP7_75t_L g196 ( .A1(n_151), .A2(n_197), .B(n_202), .Y(n_196) );
OAI21xp5_ASAP7_75t_L g210 ( .A1(n_151), .A2(n_211), .B(n_214), .Y(n_210) );
AND2x4_ASAP7_75t_L g445 ( .A(n_151), .B(n_446), .Y(n_445) );
INVx4_ASAP7_75t_SL g470 ( .A(n_151), .Y(n_470) );
NAND2x1p5_ASAP7_75t_L g503 ( .A(n_151), .B(n_446), .Y(n_503) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_153), .A2(n_210), .B(n_217), .Y(n_209) );
INVx4_ASAP7_75t_L g227 ( .A(n_153), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_153), .A2(n_493), .B(n_494), .Y(n_492) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_153), .Y(n_522) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g190 ( .A(n_154), .Y(n_190) );
AND2x2_ASAP7_75t_L g155 ( .A(n_156), .B(n_168), .Y(n_155) );
AND2x2_ASAP7_75t_L g230 ( .A(n_156), .B(n_184), .Y(n_230) );
INVx2_ASAP7_75t_L g264 ( .A(n_156), .Y(n_264) );
AND2x2_ASAP7_75t_L g279 ( .A(n_156), .B(n_185), .Y(n_279) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_156), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_156), .B(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g299 ( .A(n_156), .B(n_262), .Y(n_299) );
INVx1_ASAP7_75t_L g311 ( .A(n_156), .Y(n_311) );
INVx1_ASAP7_75t_L g352 ( .A(n_156), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_156), .B(n_252), .Y(n_405) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_161), .Y(n_158) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_165), .B(n_166), .Y(n_163) );
O2A1O1Ixp5_ASAP7_75t_L g239 ( .A1(n_166), .A2(n_203), .B(n_240), .C(n_241), .Y(n_239) );
NOR2xp67_ASAP7_75t_L g168 ( .A(n_169), .B(n_184), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g229 ( .A(n_170), .B(n_230), .Y(n_229) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_170), .Y(n_257) );
AND2x2_ASAP7_75t_SL g310 ( .A(n_170), .B(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g314 ( .A(n_170), .B(n_184), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_170), .B(n_309), .Y(n_372) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g262 ( .A(n_171), .Y(n_262) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_171), .Y(n_278) );
OR2x2_ASAP7_75t_L g351 ( .A(n_171), .B(n_352), .Y(n_351) );
O2A1O1Ixp5_ASAP7_75t_SL g173 ( .A1(n_174), .A2(n_175), .B(n_176), .C(n_177), .Y(n_173) );
INVx2_ASAP7_75t_L g188 ( .A(n_177), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_177), .A2(n_212), .B(n_213), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_177), .A2(n_237), .B(n_238), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_177), .B(n_528), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_181), .Y(n_178) );
INVx1_ASAP7_75t_L g201 ( .A(n_181), .Y(n_201) );
INVx4_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g452 ( .A(n_182), .Y(n_452) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
BUFx2_ASAP7_75t_L g258 ( .A(n_185), .Y(n_258) );
AND2x2_ASAP7_75t_L g263 ( .A(n_185), .B(n_264), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_188), .A2(n_203), .B(n_206), .C(n_207), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_188), .A2(n_215), .B(n_216), .Y(n_214) );
INVx2_ASAP7_75t_L g195 ( .A(n_190), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_190), .B(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_191), .B(n_246), .Y(n_409) );
INVx1_ASAP7_75t_SL g191 ( .A(n_192), .Y(n_191) );
OR2x2_ASAP7_75t_L g379 ( .A(n_192), .B(n_220), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_193), .B(n_209), .Y(n_192) );
AND2x2_ASAP7_75t_L g255 ( .A(n_193), .B(n_246), .Y(n_255) );
INVx2_ASAP7_75t_L g267 ( .A(n_193), .Y(n_267) );
AND2x2_ASAP7_75t_L g301 ( .A(n_193), .B(n_249), .Y(n_301) );
AND2x2_ASAP7_75t_L g368 ( .A(n_193), .B(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_194), .B(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g248 ( .A(n_194), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g288 ( .A(n_194), .B(n_209), .Y(n_288) );
AND2x2_ASAP7_75t_L g305 ( .A(n_194), .B(n_306), .Y(n_305) );
OA21x2_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B(n_208), .Y(n_194) );
OA21x2_ASAP7_75t_L g234 ( .A1(n_195), .A2(n_235), .B(n_242), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_200), .C(n_201), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_199), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_199), .A2(n_506), .B(n_507), .Y(n_505) );
O2A1O1Ixp33_ASAP7_75t_L g465 ( .A1(n_201), .A2(n_466), .B(n_467), .C(n_468), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_203), .A2(n_451), .B(n_453), .Y(n_450) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g231 ( .A(n_209), .B(n_232), .Y(n_231) );
INVx3_ASAP7_75t_L g249 ( .A(n_209), .Y(n_249) );
AND2x2_ASAP7_75t_L g254 ( .A(n_209), .B(n_234), .Y(n_254) );
AND2x2_ASAP7_75t_L g327 ( .A(n_209), .B(n_306), .Y(n_327) );
AND2x2_ASAP7_75t_L g392 ( .A(n_209), .B(n_382), .Y(n_392) );
OAI311xp33_ASAP7_75t_L g275 ( .A1(n_218), .A2(n_276), .A3(n_280), .B1(n_282), .C1(n_302), .Y(n_275) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g287 ( .A(n_219), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g346 ( .A(n_219), .B(n_254), .Y(n_346) );
AND2x2_ASAP7_75t_L g420 ( .A(n_219), .B(n_301), .Y(n_420) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_220), .B(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g355 ( .A(n_220), .Y(n_355) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx3_ASAP7_75t_L g246 ( .A(n_221), .Y(n_246) );
NOR2x1_ASAP7_75t_L g318 ( .A(n_221), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g375 ( .A(n_221), .B(n_249), .Y(n_375) );
AND2x4_ASAP7_75t_L g221 ( .A(n_222), .B(n_223), .Y(n_221) );
INVx1_ASAP7_75t_L g272 ( .A(n_222), .Y(n_272) );
AO21x1_ASAP7_75t_L g271 ( .A1(n_224), .A2(n_227), .B(n_272), .Y(n_271) );
AO21x2_ASAP7_75t_L g462 ( .A1(n_227), .A2(n_463), .B(n_472), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_227), .B(n_473), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_227), .B(n_485), .Y(n_484) );
AO21x2_ASAP7_75t_L g500 ( .A1(n_227), .A2(n_501), .B(n_508), .Y(n_500) );
INVx3_ASAP7_75t_L g530 ( .A(n_227), .Y(n_530) );
AND2x2_ASAP7_75t_L g250 ( .A(n_230), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g303 ( .A(n_230), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g383 ( .A(n_230), .B(n_384), .Y(n_383) );
AOI221xp5_ASAP7_75t_L g282 ( .A1(n_231), .A2(n_263), .B1(n_283), .B2(n_287), .C(n_289), .Y(n_282) );
INVx1_ASAP7_75t_L g407 ( .A(n_232), .Y(n_407) );
OR2x2_ASAP7_75t_L g373 ( .A(n_233), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g268 ( .A(n_234), .B(n_249), .Y(n_268) );
OR2x2_ASAP7_75t_L g270 ( .A(n_234), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g295 ( .A(n_234), .Y(n_295) );
INVx2_ASAP7_75t_L g306 ( .A(n_234), .Y(n_306) );
AND2x2_ASAP7_75t_L g333 ( .A(n_234), .B(n_271), .Y(n_333) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_234), .Y(n_362) );
AOI221xp5_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_250), .B1(n_253), .B2(n_256), .C(n_259), .Y(n_243) );
INVx1_ASAP7_75t_SL g244 ( .A(n_245), .Y(n_244) );
OR2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
AND2x2_ASAP7_75t_L g344 ( .A(n_246), .B(n_254), .Y(n_344) );
AND2x2_ASAP7_75t_L g394 ( .A(n_246), .B(n_248), .Y(n_394) );
INVx2_ASAP7_75t_SL g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g281 ( .A(n_248), .B(n_252), .Y(n_281) );
AND2x2_ASAP7_75t_L g360 ( .A(n_248), .B(n_333), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_249), .B(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g319 ( .A(n_249), .Y(n_319) );
OAI21xp33_ASAP7_75t_L g329 ( .A1(n_250), .A2(n_330), .B(n_332), .Y(n_329) );
OR2x2_ASAP7_75t_L g273 ( .A(n_251), .B(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g339 ( .A(n_251), .B(n_299), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_251), .B(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g316 ( .A(n_252), .B(n_285), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_252), .B(n_399), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_253), .B(n_279), .Y(n_389) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
AND2x2_ASAP7_75t_L g312 ( .A(n_254), .B(n_267), .Y(n_312) );
INVx1_ASAP7_75t_L g328 ( .A(n_255), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_265), .B1(n_269), .B2(n_273), .Y(n_259) );
INVx2_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
INVx2_ASAP7_75t_L g291 ( .A(n_262), .Y(n_291) );
INVx1_ASAP7_75t_L g304 ( .A(n_262), .Y(n_304) );
INVx1_ASAP7_75t_L g274 ( .A(n_263), .Y(n_274) );
AND2x2_ASAP7_75t_L g345 ( .A(n_263), .B(n_291), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_263), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_268), .Y(n_265) );
OR2x2_ASAP7_75t_L g269 ( .A(n_266), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_266), .B(n_382), .Y(n_381) );
NOR2xp67_ASAP7_75t_L g413 ( .A(n_266), .B(n_414), .Y(n_413) );
INVx3_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g416 ( .A(n_268), .B(n_368), .Y(n_416) );
INVx1_ASAP7_75t_SL g382 ( .A(n_270), .Y(n_382) );
AND2x2_ASAP7_75t_L g322 ( .A(n_271), .B(n_306), .Y(n_322) );
INVx1_ASAP7_75t_L g369 ( .A(n_271), .Y(n_369) );
OAI222xp33_ASAP7_75t_L g410 ( .A1(n_276), .A2(n_366), .B1(n_411), .B2(n_412), .C1(n_415), .C2(n_417), .Y(n_410) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx1_ASAP7_75t_L g331 ( .A(n_278), .Y(n_331) );
AND2x2_ASAP7_75t_L g342 ( .A(n_279), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_279), .B(n_384), .Y(n_411) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_281), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g386 ( .A(n_283), .Y(n_386) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_SL g324 ( .A(n_286), .Y(n_324) );
AND2x2_ASAP7_75t_L g403 ( .A(n_286), .B(n_364), .Y(n_403) );
AND2x2_ASAP7_75t_L g426 ( .A(n_286), .B(n_310), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_288), .B(n_322), .Y(n_321) );
OAI32xp33_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_292), .A3(n_294), .B1(n_296), .B2(n_300), .Y(n_289) );
BUFx2_ASAP7_75t_L g364 ( .A(n_291), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_292), .B(n_310), .Y(n_391) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g330 ( .A(n_293), .B(n_331), .Y(n_330) );
AND2x4_ASAP7_75t_L g398 ( .A(n_293), .B(n_399), .Y(n_398) );
OR2x2_ASAP7_75t_L g387 ( .A(n_294), .B(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AND2x2_ASAP7_75t_L g358 ( .A(n_297), .B(n_331), .Y(n_358) );
INVx2_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
OAI221xp5_ASAP7_75t_SL g320 ( .A1(n_299), .A2(n_321), .B1(n_323), .B2(n_325), .C(n_329), .Y(n_320) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g332 ( .A(n_301), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g338 ( .A(n_301), .B(n_322), .Y(n_338) );
AOI221xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_305), .B1(n_307), .B2(n_312), .C(n_313), .Y(n_302) );
INVx1_ASAP7_75t_L g421 ( .A(n_303), .Y(n_421) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_304), .B(n_398), .Y(n_397) );
NAND2x1p5_ASAP7_75t_L g317 ( .A(n_305), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_310), .B(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g376 ( .A(n_310), .Y(n_376) );
BUFx3_ASAP7_75t_L g399 ( .A(n_311), .Y(n_399) );
INVx1_ASAP7_75t_SL g340 ( .A(n_312), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_312), .B(n_354), .Y(n_353) );
AOI21xp33_ASAP7_75t_SL g313 ( .A1(n_314), .A2(n_315), .B(n_317), .Y(n_313) );
OAI221xp5_ASAP7_75t_L g418 ( .A1(n_314), .A2(n_415), .B1(n_419), .B2(n_421), .C(n_422), .Y(n_418) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g361 ( .A(n_319), .B(n_322), .Y(n_361) );
INVx1_ASAP7_75t_L g425 ( .A(n_319), .Y(n_425) );
INVx2_ASAP7_75t_L g414 ( .A(n_322), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_322), .B(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g367 ( .A(n_327), .B(n_368), .Y(n_367) );
OAI221xp5_ASAP7_75t_SL g334 ( .A1(n_335), .A2(n_337), .B1(n_339), .B2(n_340), .C(n_341), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_344), .B1(n_345), .B2(n_346), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_343), .A2(n_405), .B1(n_406), .B2(n_408), .Y(n_404) );
OAI21xp5_ASAP7_75t_L g422 ( .A1(n_346), .A2(n_423), .B(n_426), .Y(n_422) );
NOR4xp25_ASAP7_75t_SL g347 ( .A(n_348), .B(n_356), .C(n_365), .D(n_385), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_349), .B(n_353), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_359), .B1(n_362), .B2(n_363), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g401 ( .A(n_361), .Y(n_401) );
OAI221xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_370), .B1(n_373), .B2(n_376), .C(n_377), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g388 ( .A(n_368), .Y(n_388) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI21xp5_ASAP7_75t_SL g377 ( .A1(n_378), .A2(n_380), .B(n_383), .Y(n_377) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OAI211xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B(n_389), .C(n_390), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_392), .B1(n_393), .B2(n_394), .Y(n_390) );
CKINVDCx14_ASAP7_75t_R g400 ( .A(n_394), .Y(n_400) );
NOR3xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_410), .C(n_418), .Y(n_395) );
OAI221xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_400), .B1(n_401), .B2(n_402), .C(n_404), .Y(n_396) );
INVxp67_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
CKINVDCx16_ASAP7_75t_R g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g735 ( .A(n_430), .Y(n_735) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g743 ( .A(n_432), .Y(n_743) );
AND2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx2_ASAP7_75t_L g736 ( .A(n_436), .Y(n_736) );
AND3x1_ASAP7_75t_L g436 ( .A(n_437), .B(n_632), .C(n_689), .Y(n_436) );
NOR3xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_577), .C(n_613), .Y(n_437) );
OAI211xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_486), .B(n_532), .C(n_564), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_440), .B(n_459), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AND2x4_ASAP7_75t_L g535 ( .A(n_441), .B(n_536), .Y(n_535) );
INVx5_ASAP7_75t_L g563 ( .A(n_441), .Y(n_563) );
AND2x2_ASAP7_75t_L g636 ( .A(n_441), .B(n_552), .Y(n_636) );
AND2x2_ASAP7_75t_L g674 ( .A(n_441), .B(n_580), .Y(n_674) );
AND2x2_ASAP7_75t_L g694 ( .A(n_441), .B(n_537), .Y(n_694) );
OR2x6_ASAP7_75t_L g441 ( .A(n_442), .B(n_456), .Y(n_441) );
AOI21xp5_ASAP7_75t_SL g442 ( .A1(n_443), .A2(n_447), .B(n_455), .Y(n_442) );
BUFx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx5_ASAP7_75t_L g479 ( .A(n_448), .Y(n_479) );
INVx2_ASAP7_75t_L g454 ( .A(n_452), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_L g480 ( .A1(n_454), .A2(n_481), .B(n_482), .C(n_483), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_L g515 ( .A1(n_454), .A2(n_483), .B(n_516), .C(n_517), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_459), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_474), .Y(n_459) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_460), .Y(n_575) );
AND2x2_ASAP7_75t_L g589 ( .A(n_460), .B(n_536), .Y(n_589) );
INVx1_ASAP7_75t_L g612 ( .A(n_460), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_460), .B(n_563), .Y(n_651) );
OR2x2_ASAP7_75t_L g688 ( .A(n_460), .B(n_534), .Y(n_688) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_461), .Y(n_624) );
AND2x2_ASAP7_75t_L g631 ( .A(n_461), .B(n_537), .Y(n_631) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g552 ( .A(n_462), .B(n_537), .Y(n_552) );
BUFx2_ASAP7_75t_L g580 ( .A(n_462), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_471), .Y(n_463) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_L g524 ( .A1(n_470), .A2(n_479), .B(n_525), .C(n_526), .Y(n_524) );
O2A1O1Ixp33_ASAP7_75t_SL g539 ( .A1(n_470), .A2(n_479), .B(n_540), .C(n_541), .Y(n_539) );
INVx5_ASAP7_75t_L g534 ( .A(n_474), .Y(n_534) );
BUFx2_ASAP7_75t_L g556 ( .A(n_474), .Y(n_556) );
AND2x2_ASAP7_75t_L g713 ( .A(n_474), .B(n_567), .Y(n_713) );
OR2x6_ASAP7_75t_L g474 ( .A(n_475), .B(n_484), .Y(n_474) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND2xp33_ASAP7_75t_L g487 ( .A(n_488), .B(n_519), .Y(n_487) );
OAI221xp5_ASAP7_75t_L g613 ( .A1(n_488), .A2(n_614), .B1(n_621), .B2(n_622), .C(n_625), .Y(n_613) );
OR2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_498), .Y(n_488) );
AND2x2_ASAP7_75t_L g520 ( .A(n_489), .B(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_489), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_SL g489 ( .A(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g548 ( .A(n_490), .B(n_499), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_490), .B(n_500), .Y(n_558) );
OR2x2_ASAP7_75t_L g569 ( .A(n_490), .B(n_521), .Y(n_569) );
AND2x2_ASAP7_75t_L g572 ( .A(n_490), .B(n_560), .Y(n_572) );
AND2x2_ASAP7_75t_L g588 ( .A(n_490), .B(n_510), .Y(n_588) );
OR2x2_ASAP7_75t_L g604 ( .A(n_490), .B(n_500), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_490), .B(n_521), .Y(n_666) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_491), .B(n_510), .Y(n_658) );
AND2x2_ASAP7_75t_L g661 ( .A(n_491), .B(n_500), .Y(n_661) );
OR2x2_ASAP7_75t_L g582 ( .A(n_498), .B(n_569), .Y(n_582) );
INVx2_ASAP7_75t_L g608 ( .A(n_498), .Y(n_608) );
OR2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_510), .Y(n_498) );
AND2x2_ASAP7_75t_L g531 ( .A(n_499), .B(n_511), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_499), .B(n_521), .Y(n_587) );
OR2x2_ASAP7_75t_L g598 ( .A(n_499), .B(n_511), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_499), .B(n_560), .Y(n_657) );
OAI221xp5_ASAP7_75t_L g690 ( .A1(n_499), .A2(n_691), .B1(n_693), .B2(n_695), .C(n_698), .Y(n_690) );
INVx5_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_500), .B(n_521), .Y(n_629) );
OAI21xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_503), .B(n_504), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_510), .B(n_560), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_510), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g576 ( .A(n_510), .B(n_548), .Y(n_576) );
OR2x2_ASAP7_75t_L g620 ( .A(n_510), .B(n_521), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_510), .B(n_572), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_510), .B(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g685 ( .A(n_510), .B(n_686), .Y(n_685) );
INVx5_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_SL g549 ( .A(n_511), .B(n_520), .Y(n_549) );
O2A1O1Ixp33_ASAP7_75t_SL g553 ( .A1(n_511), .A2(n_554), .B(n_557), .C(n_561), .Y(n_553) );
OR2x2_ASAP7_75t_L g591 ( .A(n_511), .B(n_587), .Y(n_591) );
OR2x2_ASAP7_75t_L g627 ( .A(n_511), .B(n_569), .Y(n_627) );
OAI311xp33_ASAP7_75t_L g633 ( .A1(n_511), .A2(n_572), .A3(n_634), .B1(n_637), .C1(n_644), .Y(n_633) );
AND2x2_ASAP7_75t_L g684 ( .A(n_511), .B(n_521), .Y(n_684) );
AND2x2_ASAP7_75t_L g692 ( .A(n_511), .B(n_547), .Y(n_692) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_511), .Y(n_710) );
AND2x2_ASAP7_75t_L g727 ( .A(n_511), .B(n_548), .Y(n_727) );
OR2x6_ASAP7_75t_L g511 ( .A(n_512), .B(n_518), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_531), .Y(n_519) );
AND2x2_ASAP7_75t_L g555 ( .A(n_520), .B(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g711 ( .A(n_520), .Y(n_711) );
AND2x2_ASAP7_75t_L g547 ( .A(n_521), .B(n_548), .Y(n_547) );
INVx3_ASAP7_75t_L g560 ( .A(n_521), .Y(n_560) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_521), .Y(n_603) );
INVxp67_ASAP7_75t_L g642 ( .A(n_521), .Y(n_642) );
OA21x2_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B(n_529), .Y(n_521) );
OA21x2_ASAP7_75t_L g537 ( .A1(n_530), .A2(n_538), .B(n_546), .Y(n_537) );
AND2x2_ASAP7_75t_L g720 ( .A(n_531), .B(n_568), .Y(n_720) );
AOI221xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_547), .B1(n_549), .B2(n_550), .C(n_553), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_534), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g573 ( .A(n_534), .B(n_563), .Y(n_573) );
AND2x2_ASAP7_75t_L g581 ( .A(n_534), .B(n_536), .Y(n_581) );
OR2x2_ASAP7_75t_L g593 ( .A(n_534), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g611 ( .A(n_534), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g635 ( .A(n_534), .B(n_636), .Y(n_635) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_534), .Y(n_655) );
AND2x2_ASAP7_75t_L g707 ( .A(n_534), .B(n_631), .Y(n_707) );
OAI31xp33_ASAP7_75t_L g715 ( .A1(n_534), .A2(n_584), .A3(n_683), .B(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_535), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_SL g679 ( .A(n_535), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_535), .B(n_688), .Y(n_687) );
AND2x4_ASAP7_75t_L g567 ( .A(n_536), .B(n_563), .Y(n_567) );
INVx1_ASAP7_75t_L g654 ( .A(n_536), .Y(n_654) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g704 ( .A(n_537), .B(n_563), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
INVx1_ASAP7_75t_SL g714 ( .A(n_547), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_548), .B(n_619), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_549), .A2(n_661), .B1(n_699), .B2(n_702), .Y(n_698) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g562 ( .A(n_552), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g621 ( .A(n_552), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_552), .B(n_573), .Y(n_726) );
INVx1_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g696 ( .A(n_555), .B(n_697), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_556), .A2(n_615), .B(n_617), .Y(n_614) );
OR2x2_ASAP7_75t_L g622 ( .A(n_556), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g643 ( .A(n_556), .B(n_631), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_556), .B(n_654), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_556), .B(n_694), .Y(n_693) );
OAI221xp5_ASAP7_75t_SL g670 ( .A1(n_557), .A2(n_671), .B1(n_676), .B2(n_679), .C(n_680), .Y(n_670) );
OR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
OR2x2_ASAP7_75t_L g647 ( .A(n_558), .B(n_620), .Y(n_647) );
INVx1_ASAP7_75t_L g686 ( .A(n_558), .Y(n_686) );
INVx2_ASAP7_75t_L g662 ( .A(n_559), .Y(n_662) );
INVx1_ASAP7_75t_L g596 ( .A(n_560), .Y(n_596) );
INVx1_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g601 ( .A(n_563), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_563), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g630 ( .A(n_563), .B(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g718 ( .A(n_563), .B(n_688), .Y(n_718) );
AOI222xp33_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_568), .B1(n_570), .B2(n_573), .C1(n_574), .C2(n_576), .Y(n_564) );
INVxp67_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g574 ( .A(n_567), .B(n_575), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_567), .A2(n_617), .B1(n_645), .B2(n_646), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_567), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
OAI21xp33_ASAP7_75t_SL g605 ( .A1(n_576), .A2(n_606), .B(n_609), .Y(n_605) );
OAI211xp5_ASAP7_75t_SL g577 ( .A1(n_578), .A2(n_582), .B(n_583), .C(n_605), .Y(n_577) );
INVxp67_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
AOI221xp5_ASAP7_75t_L g583 ( .A1(n_581), .A2(n_584), .B1(n_589), .B2(n_590), .C(n_592), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_581), .B(n_669), .Y(n_668) );
INVxp67_ASAP7_75t_L g675 ( .A(n_581), .Y(n_675) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
AND2x2_ASAP7_75t_L g677 ( .A(n_586), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g594 ( .A(n_589), .Y(n_594) );
AND2x2_ASAP7_75t_L g600 ( .A(n_589), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_595), .B1(n_599), .B2(n_602), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_596), .B(n_608), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_597), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g697 ( .A(n_601), .Y(n_697) );
AND2x2_ASAP7_75t_L g716 ( .A(n_601), .B(n_631), .Y(n_716) );
OR2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_608), .B(n_665), .Y(n_724) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_611), .B(n_679), .Y(n_722) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g645 ( .A(n_623), .Y(n_645) );
BUFx2_ASAP7_75t_L g669 ( .A(n_624), .Y(n_669) );
OAI21xp5_ASAP7_75t_SL g625 ( .A1(n_626), .A2(n_628), .B(n_630), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NOR3xp33_ASAP7_75t_L g632 ( .A(n_633), .B(n_648), .C(n_670), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OAI21xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_640), .B(n_643), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
A2O1A1Ixp33_ASAP7_75t_SL g648 ( .A1(n_649), .A2(n_652), .B(n_656), .C(n_659), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g681 ( .A(n_649), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NOR2xp67_ASAP7_75t_SL g653 ( .A(n_654), .B(n_655), .Y(n_653) );
OR2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
INVx1_ASAP7_75t_SL g678 ( .A(n_658), .Y(n_678) );
OAI21xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_663), .B(n_667), .Y(n_659) );
AND2x4_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
AND2x2_ASAP7_75t_L g683 ( .A(n_661), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_675), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_683), .B1(n_685), .B2(n_687), .Y(n_680) );
INVx2_ASAP7_75t_SL g701 ( .A(n_688), .Y(n_701) );
NOR3xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_705), .C(n_717), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVxp67_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVxp67_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_701), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
OAI221xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_708), .B1(n_712), .B2(n_714), .C(n_715), .Y(n_705) );
A2O1A1Ixp33_ASAP7_75t_L g717 ( .A1(n_706), .A2(n_718), .B(n_719), .C(n_721), .Y(n_717) );
INVx1_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
INVxp67_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B1(n_725), .B2(n_727), .Y(n_721) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g737 ( .A(n_729), .Y(n_737) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
OAI22xp5_ASAP7_75t_SL g733 ( .A1(n_734), .A2(n_735), .B1(n_736), .B2(n_737), .Y(n_733) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
BUFx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_SL g757 ( .A(n_745), .Y(n_757) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_750), .Y(n_747) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g761 ( .A(n_749), .Y(n_761) );
INVx1_ASAP7_75t_L g754 ( .A(n_751), .Y(n_754) );
BUFx3_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
endmodule