module fake_jpeg_30835_n_442 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_442);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_442;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_10),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_15),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_47),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_48),
.B(n_53),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_49),
.Y(n_125)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_51),
.Y(n_145)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_55),
.B(n_56),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_18),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_22),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_57),
.Y(n_110)
);

INVx2_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_58),
.B(n_64),
.Y(n_109)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_18),
.B(n_15),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_13),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_65),
.B(n_68),
.Y(n_137)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_67),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_30),
.B(n_13),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_17),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_70),
.B(n_74),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_22),
.B(n_0),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_83),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_30),
.B(n_12),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_38),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_84),
.B(n_85),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_19),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_19),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_86),
.B(n_90),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_34),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_92),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_37),
.B(n_0),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_19),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_36),
.B1(n_41),
.B2(n_20),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_102),
.A2(n_103),
.B1(n_121),
.B2(n_149),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_58),
.A2(n_37),
.B1(n_26),
.B2(n_41),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

INVx3_ASAP7_75t_SL g193 ( 
.A(n_114),
.Y(n_193)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_75),
.A2(n_43),
.B(n_40),
.C(n_16),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_116),
.B(n_57),
.Y(n_157)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_119),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_56),
.A2(n_20),
.B1(n_36),
.B2(n_35),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_120),
.A2(n_128),
.B1(n_142),
.B2(n_57),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_87),
.A2(n_20),
.B1(n_44),
.B2(n_32),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_64),
.A2(n_35),
.B1(n_21),
.B2(n_16),
.Y(n_128)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_77),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_138),
.Y(n_177)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_54),
.Y(n_141)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_59),
.A2(n_21),
.B1(n_43),
.B2(n_32),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_144),
.B(n_1),
.Y(n_191)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_52),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_148),
.B(n_93),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_88),
.A2(n_26),
.B1(n_2),
.B2(n_3),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_104),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_150),
.B(n_152),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_130),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_96),
.A2(n_73),
.B1(n_81),
.B2(n_94),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_153),
.Y(n_218)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_154),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_95),
.B(n_75),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_155),
.B(n_160),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_98),
.Y(n_156)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_156),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_157),
.A2(n_158),
.B1(n_181),
.B2(n_149),
.Y(n_198)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_97),
.B(n_62),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_161),
.Y(n_212)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_107),
.Y(n_163)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_163),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_118),
.B(n_69),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_164),
.B(n_167),
.Y(n_206)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_165),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_166),
.B(n_180),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_105),
.B(n_66),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_168),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_108),
.B(n_80),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_169),
.B(n_171),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_111),
.B(n_76),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_109),
.B(n_78),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_172),
.B(n_183),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_115),
.B(n_123),
.C(n_117),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_185),
.C(n_186),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_103),
.A2(n_61),
.B1(n_72),
.B2(n_49),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_174),
.A2(n_135),
.B1(n_132),
.B2(n_143),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_137),
.B(n_47),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_175),
.B(n_195),
.Y(n_222)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_98),
.Y(n_178)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_178),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_74),
.B(n_2),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g232 ( 
.A1(n_179),
.A2(n_5),
.B(n_7),
.C(n_8),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_113),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_106),
.A2(n_67),
.B1(n_63),
.B2(n_71),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_99),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_182),
.B(n_191),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_116),
.B(n_122),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_100),
.Y(n_184)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_184),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_122),
.B(n_74),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_112),
.B(n_53),
.C(n_51),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_136),
.B(n_19),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_197),
.Y(n_214)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_124),
.Y(n_188)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_188),
.Y(n_234)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_124),
.Y(n_189)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_131),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_190),
.Y(n_236)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_100),
.Y(n_192)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_106),
.Y(n_194)
);

BUFx4f_ASAP7_75t_L g201 ( 
.A(n_194),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_145),
.B(n_51),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_110),
.B(n_53),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_196),
.Y(n_199)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_132),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_198),
.A2(n_202),
.B1(n_204),
.B2(n_216),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_200),
.A2(n_209),
.B1(n_185),
.B2(n_193),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_158),
.A2(n_102),
.B1(n_121),
.B2(n_143),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_L g204 ( 
.A1(n_170),
.A2(n_140),
.B1(n_127),
.B2(n_135),
.Y(n_204)
);

AO22x1_ASAP7_75t_L g207 ( 
.A1(n_183),
.A2(n_114),
.B1(n_140),
.B2(n_127),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_207),
.A2(n_179),
.B(n_169),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_183),
.A2(n_139),
.B1(n_131),
.B2(n_133),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_177),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_233),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_161),
.A2(n_139),
.B1(n_133),
.B2(n_114),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_213),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_160),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_155),
.B(n_1),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_229),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_164),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_227),
.A2(n_163),
.B1(n_188),
.B2(n_159),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_167),
.B(n_11),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_232),
.A2(n_187),
.B(n_185),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_156),
.Y(n_233)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_238),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_173),
.C(n_172),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_240),
.B(n_247),
.C(n_254),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_176),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_241),
.B(n_246),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_242),
.Y(n_285)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_244),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_245),
.B(n_257),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_201),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_203),
.B(n_172),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_248),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_201),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_249),
.Y(n_283)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_215),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_250),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_251),
.A2(n_253),
.B1(n_255),
.B2(n_207),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_206),
.A2(n_208),
.B1(n_218),
.B2(n_204),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_171),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_206),
.A2(n_154),
.B1(n_165),
.B2(n_168),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_189),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_264),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_223),
.B(n_162),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_219),
.Y(n_258)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_187),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_210),
.C(n_220),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_SL g295 ( 
.A(n_260),
.B(n_207),
.C(n_232),
.Y(n_295)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_261),
.Y(n_294)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_226),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_268),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_209),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_214),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_269),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_218),
.A2(n_186),
.B(n_197),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_266),
.Y(n_298)
);

BUFx5_ASAP7_75t_L g267 ( 
.A(n_236),
.Y(n_267)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_267),
.Y(n_275)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_230),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_234),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_230),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_270),
.B(n_272),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_201),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_271),
.Y(n_287)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_234),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_280),
.B(n_281),
.C(n_296),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_247),
.B(n_210),
.Y(n_281)
);

INVxp33_ASAP7_75t_L g282 ( 
.A(n_239),
.Y(n_282)
);

OAI21xp33_ASAP7_75t_SL g307 ( 
.A1(n_282),
.A2(n_295),
.B(n_260),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_222),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_284),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_243),
.A2(n_208),
.B1(n_253),
.B2(n_240),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_286),
.A2(n_269),
.B1(n_244),
.B2(n_250),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_292),
.A2(n_243),
.B1(n_245),
.B2(n_242),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_254),
.B(n_214),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_267),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_297),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_251),
.A2(n_202),
.B1(n_216),
.B2(n_227),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_300),
.A2(n_252),
.B1(n_200),
.B2(n_262),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_239),
.B(n_199),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_301),
.B(n_151),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_259),
.B(n_229),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_252),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_266),
.B(n_225),
.C(n_228),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_281),
.C(n_276),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_275),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_306),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_307),
.A2(n_327),
.B1(n_287),
.B2(n_283),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_290),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_308),
.B(n_312),
.Y(n_333)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_290),
.Y(n_309)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_309),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_310),
.A2(n_313),
.B1(n_285),
.B2(n_298),
.Y(n_334)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_275),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_311),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_291),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_298),
.A2(n_255),
.B1(n_242),
.B2(n_238),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_314),
.Y(n_344)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_315),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_316),
.B(n_292),
.Y(n_341)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_299),
.Y(n_317)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_317),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_318),
.B(n_319),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_274),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_320),
.B(n_321),
.C(n_329),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_276),
.B(n_296),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_282),
.B(n_224),
.Y(n_323)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_323),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_277),
.B(n_248),
.Y(n_324)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_324),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_286),
.B(n_263),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_325),
.A2(n_328),
.B1(n_330),
.B2(n_331),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_279),
.B(n_224),
.Y(n_326)
);

INVxp33_ASAP7_75t_L g351 ( 
.A(n_326),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_300),
.A2(n_261),
.B1(n_268),
.B2(n_270),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_294),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_280),
.B(n_272),
.C(n_236),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_294),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_334),
.A2(n_346),
.B1(n_271),
.B2(n_249),
.Y(n_373)
);

AO22x1_ASAP7_75t_L g335 ( 
.A1(n_308),
.A2(n_295),
.B1(n_285),
.B2(n_277),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_335),
.B(n_304),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_321),
.B(n_302),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_338),
.B(n_339),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_305),
.B(n_303),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_324),
.Y(n_340)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_340),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_341),
.B(n_355),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_320),
.B(n_273),
.C(n_288),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_345),
.B(n_348),
.C(n_353),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_305),
.B(n_329),
.C(n_316),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_318),
.B(n_293),
.C(n_289),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_314),
.B(n_289),
.C(n_258),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_354),
.B(n_304),
.C(n_328),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_309),
.B(n_278),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_344),
.A2(n_313),
.B1(n_317),
.B2(n_315),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_359),
.B(n_360),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_333),
.B(n_322),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_332),
.Y(n_361)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_361),
.Y(n_379)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_347),
.Y(n_362)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_362),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_345),
.B(n_319),
.Y(n_363)
);

OAI21x1_ASAP7_75t_L g389 ( 
.A1(n_363),
.A2(n_351),
.B(n_337),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_352),
.B(n_312),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_364),
.B(n_370),
.Y(n_388)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_349),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_366),
.A2(n_368),
.B(n_237),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_367),
.B(n_335),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g368 ( 
.A(n_350),
.B(n_311),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_369),
.B(n_372),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_336),
.B(n_331),
.C(n_306),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_338),
.B(n_336),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_373),
.A2(n_355),
.B1(n_337),
.B2(n_353),
.Y(n_387)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_356),
.Y(n_374)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_374),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_348),
.B(n_278),
.C(n_219),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_375),
.B(n_376),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_339),
.B(n_190),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_343),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_377),
.Y(n_393)
);

BUFx12_ASAP7_75t_L g380 ( 
.A(n_368),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_380),
.B(n_366),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_386),
.Y(n_398)
);

OAI22xp33_ASAP7_75t_L g385 ( 
.A1(n_367),
.A2(n_344),
.B1(n_354),
.B2(n_334),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_385),
.A2(n_387),
.B1(n_390),
.B2(n_376),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_371),
.B(n_341),
.Y(n_386)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_389),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_358),
.A2(n_342),
.B1(n_351),
.B2(n_246),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_391),
.B(n_237),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_394),
.B(n_396),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_385),
.A2(n_369),
.B1(n_359),
.B2(n_357),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_395),
.B(n_386),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_384),
.B(n_370),
.C(n_365),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_397),
.B(n_404),
.C(n_205),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_382),
.A2(n_365),
.B(n_375),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_399),
.B(n_403),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_383),
.B(n_357),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_400),
.B(n_402),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_401),
.B(n_381),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_383),
.B(n_371),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_378),
.B(n_372),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_384),
.B(n_205),
.C(n_151),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_388),
.B(n_162),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_406),
.B(n_380),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_409),
.B(n_416),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_410),
.B(n_415),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_405),
.B(n_393),
.Y(n_411)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_411),
.Y(n_426)
);

OAI321xp33_ASAP7_75t_L g412 ( 
.A1(n_395),
.A2(n_380),
.A3(n_393),
.B1(n_378),
.B2(n_379),
.C(n_392),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_412),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_413),
.A2(n_193),
.B1(n_178),
.B2(n_184),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_397),
.A2(n_404),
.B(n_398),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_402),
.A2(n_398),
.B(n_400),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_417),
.B(n_221),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_418),
.A2(n_410),
.B(n_413),
.Y(n_427)
);

AO21x1_ASAP7_75t_L g431 ( 
.A1(n_419),
.A2(n_421),
.B(n_426),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_414),
.A2(n_192),
.B(n_194),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_407),
.A2(n_221),
.B(n_7),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_422),
.B(n_424),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_423),
.B(n_9),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_408),
.B(n_9),
.C(n_11),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_427),
.Y(n_436)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_428),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_420),
.B(n_415),
.Y(n_430)
);

OR2x2_ASAP7_75t_L g434 ( 
.A(n_430),
.B(n_431),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_425),
.B(n_11),
.C(n_424),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_432),
.B(n_429),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_435),
.B(n_418),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_437),
.Y(n_439)
);

AOI21x1_ASAP7_75t_L g438 ( 
.A1(n_434),
.A2(n_422),
.B(n_436),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_439),
.B(n_433),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_440),
.B(n_438),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_441),
.Y(n_442)
);


endmodule