module fake_jpeg_7206_n_96 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_96);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_96;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_62;
wire n_43;
wire n_82;

INVx2_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_54),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_44),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_4),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_22),
.Y(n_74)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_6),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_54),
.A2(n_47),
.B1(n_45),
.B2(n_43),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_59),
.A2(n_61),
.B1(n_68),
.B2(n_72),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_56),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_27),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_41),
.B1(n_42),
.B2(n_46),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_64),
.B(n_66),
.Y(n_78)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_65),
.Y(n_77)
);

CKINVDCx12_ASAP7_75t_R g66 ( 
.A(n_52),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_50),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_68)
);

NAND3xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_13),
.C(n_14),
.Y(n_69)
);

OR2x2_ASAP7_75t_SL g81 ( 
.A(n_69),
.B(n_73),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_15),
.Y(n_70)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_70),
.B(n_74),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g73 ( 
.A1(n_50),
.A2(n_19),
.B(n_20),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_63),
.B(n_28),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_29),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_84),
.B(n_78),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_85),
.A2(n_71),
.B(n_82),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_81),
.B(n_79),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_80),
.C(n_83),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_L g89 ( 
.A1(n_88),
.A2(n_76),
.B(n_77),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_75),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_61),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_92),
.B(n_30),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_31),
.B(n_32),
.Y(n_94)
);

BUFx24_ASAP7_75t_SL g95 ( 
.A(n_94),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_35),
.Y(n_96)
);


endmodule