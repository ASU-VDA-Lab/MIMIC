module fake_jpeg_5406_n_340 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_10),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_16),
.B(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_36),
.B(n_44),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_0),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_41),
.Y(n_57)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_42),
.B1(n_19),
.B2(n_31),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_23),
.B(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_30),
.Y(n_72)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_47),
.Y(n_90)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_50),
.Y(n_93)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_53),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_19),
.B1(n_31),
.B2(n_24),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_54),
.A2(n_58),
.B1(n_17),
.B2(n_38),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_42),
.B1(n_23),
.B2(n_24),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_56),
.A2(n_73),
.B1(n_74),
.B2(n_40),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_45),
.B1(n_36),
.B2(n_35),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_62),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_71),
.Y(n_98)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_38),
.B(n_26),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_38),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_83),
.B(n_84),
.Y(n_113)
);

AOI32xp33_ASAP7_75t_L g84 ( 
.A1(n_64),
.A2(n_37),
.A3(n_25),
.B1(n_40),
.B2(n_42),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_38),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_86),
.A2(n_88),
.B(n_97),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_49),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_66),
.A2(n_40),
.B1(n_27),
.B2(n_17),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_91),
.A2(n_52),
.B1(n_50),
.B2(n_60),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_94),
.A2(n_68),
.B1(n_70),
.B2(n_59),
.Y(n_103)
);

AND2x4_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_28),
.Y(n_97)
);

AND2x4_ASAP7_75t_SL g107 ( 
.A(n_97),
.B(n_83),
.Y(n_107)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_99),
.B(n_102),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_61),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_109),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_75),
.B1(n_97),
.B2(n_88),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_101),
.A2(n_105),
.B1(n_55),
.B2(n_57),
.Y(n_146)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_103),
.A2(n_84),
.B1(n_80),
.B2(n_85),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_63),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_104),
.B(n_121),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_75),
.B1(n_97),
.B2(n_88),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_77),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_106),
.B(n_108),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_118),
.B(n_125),
.Y(n_126)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_77),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_110),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_45),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_112),
.Y(n_142)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_86),
.A2(n_70),
.B1(n_68),
.B2(n_73),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_114),
.A2(n_115),
.B1(n_92),
.B2(n_96),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_98),
.A2(n_67),
.B1(n_36),
.B2(n_37),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_81),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_116),
.Y(n_144)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_28),
.Y(n_150)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_48),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_97),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_124),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_113),
.C(n_124),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_113),
.C(n_151),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_131),
.A2(n_139),
.B1(n_146),
.B2(n_95),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_92),
.B1(n_96),
.B2(n_95),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_132),
.A2(n_133),
.B1(n_141),
.B2(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_134),
.B(n_135),
.Y(n_181)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_136),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_101),
.A2(n_83),
.B1(n_69),
.B2(n_82),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_82),
.B1(n_78),
.B2(n_37),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_148),
.Y(n_156)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_152),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_SL g173 ( 
.A(n_150),
.B(n_28),
.C(n_20),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_122),
.A2(n_107),
.B1(n_119),
.B2(n_113),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_107),
.A2(n_26),
.B(n_79),
.C(n_95),
.Y(n_153)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_145),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_155),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_177),
.C(n_150),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_129),
.A2(n_107),
.B1(n_105),
.B2(n_102),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_158),
.Y(n_209)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_154),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_165),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_129),
.A2(n_108),
.B1(n_118),
.B2(n_116),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_160),
.A2(n_183),
.B1(n_147),
.B2(n_33),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_145),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_161),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_126),
.A2(n_112),
.B(n_109),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_162),
.A2(n_33),
.B(n_149),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_144),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_168),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_136),
.A2(n_65),
.B1(n_47),
.B2(n_46),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_170),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_127),
.B(n_110),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_153),
.A2(n_106),
.B1(n_87),
.B2(n_79),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_171),
.A2(n_134),
.B1(n_128),
.B2(n_143),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_130),
.B(n_87),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_179),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_173),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_126),
.B(n_28),
.Y(n_174)
);

A2O1A1O1Ixp25_ASAP7_75t_L g206 ( 
.A1(n_174),
.A2(n_33),
.B(n_18),
.C(n_29),
.D(n_3),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_178),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_78),
.C(n_51),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_127),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_20),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_144),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_18),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_131),
.A2(n_120),
.B1(n_117),
.B2(n_99),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_186),
.C(n_158),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_152),
.C(n_138),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_135),
.Y(n_187)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_138),
.Y(n_190)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_200),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_163),
.A2(n_133),
.B1(n_153),
.B2(n_141),
.Y(n_192)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_192),
.Y(n_222)
);

OAI32xp33_ASAP7_75t_L g195 ( 
.A1(n_166),
.A2(n_128),
.A3(n_140),
.B1(n_32),
.B2(n_30),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_181),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_166),
.A2(n_137),
.B1(n_147),
.B2(n_148),
.Y(n_198)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_198),
.Y(n_227)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_204),
.Y(n_233)
);

NAND3xp33_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_20),
.C(n_33),
.Y(n_200)
);

OAI22x1_ASAP7_75t_SL g201 ( 
.A1(n_174),
.A2(n_32),
.B1(n_28),
.B2(n_20),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_201),
.A2(n_207),
.B1(n_175),
.B2(n_159),
.Y(n_213)
);

OA21x2_ASAP7_75t_L g203 ( 
.A1(n_162),
.A2(n_137),
.B(n_32),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_203),
.A2(n_206),
.B(n_1),
.Y(n_237)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_205),
.A2(n_164),
.B(n_180),
.Y(n_224)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_161),
.B(n_18),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_211),
.B(n_0),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_SL g255 ( 
.A(n_212),
.B(n_213),
.C(n_224),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_218),
.C(n_225),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_164),
.Y(n_215)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_215),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_184),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_216),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_172),
.C(n_176),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_179),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_221),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_177),
.Y(n_221)
);

INVxp33_ASAP7_75t_L g223 ( 
.A(n_211),
.Y(n_223)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_223),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_160),
.C(n_183),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_209),
.A2(n_165),
.B1(n_173),
.B2(n_182),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_231),
.Y(n_245)
);

XNOR2x1_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_182),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_232),
.Y(n_247)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_15),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_201),
.Y(n_234)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_15),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_191),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_236),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_237),
.A2(n_202),
.B(n_189),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_233),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_238),
.B(n_256),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_204),
.Y(n_239)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

INVxp33_ASAP7_75t_SL g240 ( 
.A(n_230),
.Y(n_240)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_240),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_199),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_260),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_257),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_222),
.A2(n_197),
.B1(n_202),
.B2(n_207),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_251),
.A2(n_254),
.B1(n_234),
.B2(n_220),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_228),
.B(n_188),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_252),
.B(n_188),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_227),
.A2(n_224),
.B1(n_234),
.B2(n_212),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_213),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_226),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_258),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_221),
.B(n_187),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_259),
.B(n_219),
.Y(n_261)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_232),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_261),
.B(n_276),
.Y(n_290)
);

AOI21x1_ASAP7_75t_L g262 ( 
.A1(n_243),
.A2(n_203),
.B(n_195),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_262),
.A2(n_265),
.B(n_267),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_218),
.C(n_214),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_263),
.A2(n_275),
.B(n_276),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_253),
.A2(n_243),
.B1(n_260),
.B2(n_244),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_255),
.Y(n_268)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

INVxp67_ASAP7_75t_SL g269 ( 
.A(n_253),
.Y(n_269)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_269),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_242),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_196),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_272),
.A2(n_248),
.B(n_250),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_245),
.A2(n_225),
.B1(n_196),
.B2(n_229),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_273),
.A2(n_279),
.B1(n_247),
.B2(n_235),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_241),
.B(n_193),
.C(n_192),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_246),
.C(n_257),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_242),
.A2(n_193),
.B1(n_203),
.B2(n_237),
.Y(n_279)
);

OR2x2_ASAP7_75t_SL g281 ( 
.A(n_274),
.B(n_255),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_272),
.Y(n_300)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_282),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_223),
.Y(n_284)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_284),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_262),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_285),
.B(n_1),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_273),
.B(n_249),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_294),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_289),
.A2(n_283),
.B(n_270),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_291),
.C(n_292),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_246),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_268),
.A2(n_254),
.B(n_251),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_293),
.A2(n_295),
.B1(n_14),
.B2(n_13),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_265),
.B(n_247),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_278),
.A2(n_206),
.B1(n_2),
.B2(n_3),
.Y(n_295)
);

AOI211xp5_ASAP7_75t_L g299 ( 
.A1(n_288),
.A2(n_266),
.B(n_264),
.C(n_279),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_306),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_300),
.A2(n_13),
.B(n_12),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_277),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_301),
.A2(n_304),
.B(n_288),
.Y(n_310)
);

NOR3xp33_ASAP7_75t_SL g303 ( 
.A(n_292),
.B(n_275),
.C(n_270),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_11),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_280),
.B(n_263),
.C(n_2),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_307),
.C(n_6),
.Y(n_320)
);

NOR2x1_ASAP7_75t_R g306 ( 
.A(n_281),
.B(n_14),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_1),
.C(n_3),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_309),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_310),
.A2(n_311),
.B(n_313),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_300),
.B(n_293),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_302),
.A2(n_290),
.B(n_295),
.Y(n_313)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_314),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_316),
.C(n_317),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_302),
.A2(n_4),
.B(n_5),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_298),
.A2(n_11),
.B1(n_6),
.B2(n_7),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_5),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_297),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_320),
.B(n_307),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_315),
.Y(n_321)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_321),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_325),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_306),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_326),
.A2(n_328),
.B(n_6),
.Y(n_332)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_327),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_303),
.Y(n_328)
);

OAI21xp33_ASAP7_75t_SL g331 ( 
.A1(n_324),
.A2(n_299),
.B(n_305),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_331),
.Y(n_336)
);

AOI321xp33_ASAP7_75t_L g335 ( 
.A1(n_332),
.A2(n_333),
.A3(n_322),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_335)
);

AOI31xp33_ASAP7_75t_L g333 ( 
.A1(n_321),
.A2(n_6),
.A3(n_7),
.B(n_8),
.Y(n_333)
);

NAND3xp33_ASAP7_75t_L g337 ( 
.A(n_335),
.B(n_334),
.C(n_329),
.Y(n_337)
);

OAI321xp33_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_336),
.A3(n_330),
.B1(n_323),
.B2(n_10),
.C(n_9),
.Y(n_338)
);

NAND4xp25_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_10),
.Y(n_340)
);


endmodule