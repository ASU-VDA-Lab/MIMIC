module real_jpeg_2028_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_1),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_54),
.Y(n_102)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_3),
.B(n_43),
.Y(n_42)
);

O2A1O1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_3),
.A2(n_5),
.B(n_34),
.C(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_3),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_3),
.B(n_86),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_3),
.B(n_23),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_3),
.A2(n_30),
.B1(n_34),
.B2(n_76),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_3),
.B(n_52),
.C(n_63),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_76),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_3),
.B(n_57),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_3),
.B(n_71),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_4),
.A2(n_51),
.B1(n_52),
.B2(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_4),
.Y(n_113)
);

AO22x2_ASAP7_75t_L g23 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_23)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

O2A1O1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_5),
.A2(n_23),
.B(n_34),
.C(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_5),
.B(n_34),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_6),
.A2(n_51),
.B1(n_52),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_6),
.Y(n_59)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_7),
.Y(n_88)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_10),
.A2(n_30),
.B1(n_34),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_37),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_10),
.A2(n_37),
.B1(n_51),
.B2(n_52),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_10),
.A2(n_37),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_68),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_11),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_11),
.A2(n_30),
.B1(n_34),
.B2(n_68),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_11),
.A2(n_51),
.B1(n_52),
.B2(n_68),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_13),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_13),
.A2(n_24),
.B1(n_25),
.B2(n_33),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_13),
.A2(n_33),
.B1(n_51),
.B2(n_52),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_116),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_115),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_81),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_19),
.B(n_81),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_60),
.C(n_73),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_20),
.B(n_172),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_40),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_21),
.B(n_41),
.C(n_49),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_28),
.B(n_35),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_23),
.A2(n_29),
.B1(n_38),
.B2(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_23),
.B(n_36),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_24),
.A2(n_25),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_L g75 ( 
.A1(n_24),
.A2(n_27),
.B(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_25),
.B(n_143),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_30),
.A2(n_34),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

NAND2xp33_ASAP7_75t_SL g108 ( 
.A(n_30),
.B(n_46),
.Y(n_108)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI32xp33_ASAP7_75t_L g107 ( 
.A1(n_34),
.A2(n_45),
.A3(n_87),
.B1(n_91),
.B2(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_38),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_48),
.B2(n_49),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_44),
.B(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_45),
.A2(n_46),
.B1(n_86),
.B2(n_87),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_50),
.A2(n_56),
.B(n_78),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_52),
.B1(n_63),
.B2(n_64),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_52),
.B(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_55),
.A2(n_126),
.B(n_127),
.Y(n_125)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_55),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_55),
.A2(n_56),
.B1(n_126),
.B2(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_56),
.B(n_80),
.Y(n_128)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_57),
.A2(n_79),
.B(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_60),
.B(n_73),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_66),
.B(n_69),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_61),
.B(n_72),
.Y(n_103)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_65),
.A2(n_101),
.B(n_103),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_65),
.A2(n_103),
.B(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_65),
.A2(n_67),
.B1(n_122),
.B2(n_136),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_70),
.A2(n_136),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_74),
.B(n_77),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_87),
.B(n_90),
.C(n_92),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_76),
.A2(n_128),
.B(n_156),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_104),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_95),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_89),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_99),
.B2(n_100),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_114),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_170),
.B(n_174),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_138),
.B(n_169),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_129),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_119),
.B(n_129),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.C(n_124),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_121),
.B1(n_123),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_124),
.A2(n_125),
.B1(n_147),
.B2(n_149),
.Y(n_146)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_137),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_135),
.C(n_137),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_133),
.B(n_134),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_150),
.B(n_168),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_146),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_146),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_141),
.A2(n_142),
.B1(n_144),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_147),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_162),
.B(n_167),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_157),
.B(n_161),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_160),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_165),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_173),
.Y(n_174)
);


endmodule