module fake_jpeg_25065_n_257 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_257);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx3_ASAP7_75t_SL g25 ( 
.A(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_14),
.B(n_12),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_31),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_26),
.B1(n_17),
.B2(n_23),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_37),
.A2(n_24),
.B1(n_33),
.B2(n_32),
.Y(n_65)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_23),
.B1(n_17),
.B2(n_26),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_48),
.B1(n_25),
.B2(n_17),
.Y(n_54)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_32),
.A2(n_17),
.B1(n_23),
.B2(n_25),
.Y(n_48)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

OAI21xp33_ASAP7_75t_L g82 ( 
.A1(n_51),
.A2(n_57),
.B(n_59),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_54),
.A2(n_60),
.B1(n_50),
.B2(n_71),
.Y(n_91)
);

NAND2xp33_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_25),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_49),
.B(n_28),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_56),
.B(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_32),
.B1(n_25),
.B2(n_28),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_60),
.A2(n_44),
.B1(n_29),
.B2(n_24),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_16),
.B1(n_27),
.B2(n_21),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_62),
.A2(n_68),
.B1(n_47),
.B2(n_24),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_63),
.B(n_64),
.Y(n_74)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_48),
.B1(n_49),
.B2(n_39),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_30),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_29),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_42),
.A2(n_27),
.B1(n_21),
.B2(n_16),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_39),
.B(n_33),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_33),
.B(n_36),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_47),
.Y(n_72)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_75),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_78),
.A2(n_92),
.B1(n_53),
.B2(n_55),
.Y(n_104)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_84),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_66),
.Y(n_105)
);

INVxp33_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_88),
.Y(n_115)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_89),
.B(n_51),
.Y(n_100)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_96),
.B1(n_57),
.B2(n_71),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_50),
.B1(n_44),
.B2(n_36),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_93),
.Y(n_111)
);

BUFx8_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

CKINVDCx12_ASAP7_75t_R g95 ( 
.A(n_63),
.Y(n_95)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_92),
.B1(n_91),
.B2(n_54),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_97),
.A2(n_104),
.B1(n_117),
.B2(n_118),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_59),
.B1(n_64),
.B2(n_71),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_101),
.B1(n_112),
.B2(n_76),
.Y(n_126)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_105),
.A2(n_113),
.B(n_116),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_77),
.B(n_56),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_110),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_77),
.B(n_35),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_90),
.A2(n_35),
.B1(n_58),
.B2(n_61),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_87),
.A2(n_22),
.B(n_61),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_86),
.B(n_15),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_119),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_29),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_81),
.A2(n_58),
.B1(n_15),
.B2(n_20),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_74),
.A2(n_83),
.B1(n_82),
.B2(n_89),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_20),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_120),
.A2(n_22),
.B(n_94),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_20),
.Y(n_121)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_101),
.A2(n_79),
.B1(n_76),
.B2(n_73),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_126),
.B1(n_131),
.B2(n_120),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_111),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_124),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_79),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_127),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_22),
.B(n_94),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_128),
.B(n_135),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_103),
.A2(n_73),
.B1(n_15),
.B2(n_20),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_94),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_144),
.Y(n_173)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_136),
.Y(n_158)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_143),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_15),
.B1(n_18),
.B2(n_13),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_138),
.A2(n_142),
.B1(n_114),
.B2(n_99),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_18),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_140),
.B(n_99),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_147),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_104),
.A2(n_22),
.B1(n_18),
.B2(n_13),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_115),
.B(n_10),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_148),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_102),
.A2(n_22),
.B(n_1),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_113),
.A2(n_18),
.B(n_13),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_0),
.Y(n_170)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_145),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_152),
.Y(n_178)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_170),
.B1(n_175),
.B2(n_142),
.Y(n_179)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_161),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_157),
.A2(n_168),
.B1(n_150),
.B2(n_130),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_149),
.A2(n_97),
.B1(n_102),
.B2(n_116),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_159),
.A2(n_132),
.B1(n_127),
.B2(n_147),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_116),
.C(n_119),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_165),
.C(n_176),
.Y(n_189)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_113),
.C(n_120),
.Y(n_165)
);

OAI32xp33_ASAP7_75t_L g166 ( 
.A1(n_130),
.A2(n_110),
.A3(n_117),
.B1(n_111),
.B2(n_122),
.Y(n_166)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_149),
.A2(n_107),
.B1(n_13),
.B2(n_2),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_129),
.B(n_10),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_169),
.Y(n_187)
);

XOR2x1_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_0),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_1),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_129),
.B(n_0),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_133),
.B(n_1),
.C(n_2),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_177),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_179),
.B(n_185),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_163),
.Y(n_181)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_154),
.A2(n_132),
.B1(n_131),
.B2(n_148),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_184),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_174),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_137),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_190),
.A2(n_160),
.B(n_164),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_156),
.B(n_144),
.C(n_2),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_195),
.C(n_176),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_194),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_193),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_1),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_173),
.C(n_159),
.Y(n_195)
);

BUFx12_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

INVxp33_ASAP7_75t_SL g220 ( 
.A(n_196),
.Y(n_220)
);

AO221x1_ASAP7_75t_L g197 ( 
.A1(n_180),
.A2(n_172),
.B1(n_171),
.B2(n_162),
.C(n_158),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_198),
.A2(n_207),
.B1(n_186),
.B2(n_183),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_199),
.A2(n_190),
.B1(n_4),
.B2(n_5),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_210),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_172),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_204),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_169),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_192),
.Y(n_219)
);

NAND3xp33_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_174),
.C(n_166),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_209),
.A2(n_190),
.B(n_177),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_168),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_199),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_212),
.A2(n_204),
.B(n_202),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_206),
.A2(n_184),
.B1(n_191),
.B2(n_189),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_189),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_216),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_188),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_208),
.B(n_194),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_217),
.B(n_219),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_222),
.A2(n_220),
.B1(n_196),
.B2(n_200),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_214),
.A2(n_203),
.B1(n_222),
.B2(n_197),
.Y(n_223)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

XNOR2x1_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_218),
.Y(n_224)
);

OAI21x1_ASAP7_75t_L g234 ( 
.A1(n_224),
.A2(n_205),
.B(n_196),
.Y(n_234)
);

OAI21x1_ASAP7_75t_L g226 ( 
.A1(n_221),
.A2(n_202),
.B(n_201),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_196),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_228),
.B(n_3),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_231),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_215),
.B(n_201),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_232),
.A2(n_220),
.B1(n_218),
.B2(n_205),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_233),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_234),
.A2(n_240),
.B(n_4),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_227),
.B(n_225),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_238),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_3),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_239),
.B(n_3),
.Y(n_242)
);

OAI221xp5_ASAP7_75t_L g241 ( 
.A1(n_233),
.A2(n_224),
.B1(n_230),
.B2(n_225),
.C(n_6),
.Y(n_241)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_241),
.Y(n_247)
);

AOI21xp33_ASAP7_75t_L g250 ( 
.A1(n_242),
.A2(n_244),
.B(n_246),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_237),
.C(n_6),
.Y(n_249)
);

INVxp33_ASAP7_75t_L g246 ( 
.A(n_236),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_238),
.Y(n_248)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_248),
.Y(n_252)
);

AOI322xp5_ASAP7_75t_L g253 ( 
.A1(n_249),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_220),
.C1(n_243),
.C2(n_223),
.Y(n_253)
);

OAI21x1_ASAP7_75t_L g251 ( 
.A1(n_247),
.A2(n_4),
.B(n_7),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_251),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_250),
.C(n_249),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_254),
.B(n_255),
.Y(n_256)
);

OAI21x1_ASAP7_75t_L g257 ( 
.A1(n_256),
.A2(n_252),
.B(n_8),
.Y(n_257)
);


endmodule