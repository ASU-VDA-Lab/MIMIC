module fake_netlist_5_1660_n_1038 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_226, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_225, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_223, n_188, n_190, n_8, n_201, n_158, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_222, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_1038);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_222;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_1038;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_380;
wire n_419;
wire n_318;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_316;
wire n_785;
wire n_389;
wire n_855;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_605;
wire n_776;
wire n_928;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_916;
wire n_452;
wire n_885;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_998;
wire n_841;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_719;
wire n_372;
wire n_443;
wire n_293;
wire n_244;
wire n_677;
wire n_864;
wire n_859;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_946;
wire n_612;
wire n_1001;
wire n_498;
wire n_385;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_509;
wire n_568;
wire n_947;
wire n_373;
wire n_820;
wire n_757;
wire n_936;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1032;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_394;
wire n_250;
wire n_579;
wire n_992;
wire n_938;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_406;
wire n_519;
wire n_470;
wire n_919;
wire n_782;
wire n_908;
wire n_325;
wire n_449;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_654;
wire n_370;
wire n_976;
wire n_234;
wire n_343;
wire n_379;
wire n_308;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_795;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_347;
wire n_763;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_622;
wire n_723;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_344;
wire n_287;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_922;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_816;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_680;
wire n_974;
wire n_432;
wire n_395;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_236;
wire n_388;
wire n_761;
wire n_1012;
wire n_1019;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1015;
wire n_1000;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_963;
wire n_954;
wire n_627;
wire n_767;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_707;
wire n_710;
wire n_832;
wire n_695;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_561;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_403;
wire n_453;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1025;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_952;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_809;
wire n_811;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_960;
wire n_759;
wire n_1018;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_904;
wire n_985;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_38),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_181),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_6),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_189),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_88),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_18),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_152),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_34),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_23),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_176),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_215),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_115),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_36),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_103),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_134),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_207),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_21),
.Y(n_243)
);

BUFx8_ASAP7_75t_SL g244 ( 
.A(n_142),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_182),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_128),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_145),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_18),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_90),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_165),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_13),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_120),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_117),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_50),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_204),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_66),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_129),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_143),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_114),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_163),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_31),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_150),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_62),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_74),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_208),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_110),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_201),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_70),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_109),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_79),
.Y(n_271)
);

BUFx10_ASAP7_75t_L g272 ( 
.A(n_147),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_200),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_27),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_54),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_95),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_151),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_211),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_26),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_212),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_12),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_131),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_48),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_53),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_210),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_20),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_31),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_5),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_44),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_154),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_184),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_46),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_223),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_0),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_4),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_20),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_155),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_93),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_205),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_17),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_12),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_87),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_193),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_17),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_162),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_25),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_60),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_35),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_57),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_203),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_11),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_61),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_179),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_106),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_170),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_100),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_123),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_171),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_213),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_73),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_125),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_164),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_144),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_243),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_229),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_252),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_229),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_236),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_274),
.B(n_0),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_231),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_261),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_281),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_281),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_279),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_227),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_231),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_296),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_311),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_240),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_227),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_249),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_249),
.Y(n_342)
);

NAND2xp33_ASAP7_75t_R g343 ( 
.A(n_228),
.B(n_1),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_320),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_241),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_278),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_278),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_242),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_285),
.B(n_1),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_245),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_246),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_230),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_251),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_230),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_237),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_253),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_255),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_272),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_285),
.B(n_2),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_247),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_257),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_237),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_263),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_254),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_258),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_265),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_263),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_244),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_256),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_244),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_259),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_260),
.Y(n_372)
);

BUFx6f_ASAP7_75t_SL g373 ( 
.A(n_272),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_266),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_235),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_267),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_286),
.B(n_2),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_264),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_235),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_348),
.Y(n_380)
);

OA21x2_ASAP7_75t_L g381 ( 
.A1(n_351),
.A2(n_250),
.B(n_239),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_360),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_334),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_346),
.B(n_291),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_337),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_364),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_338),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_369),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_378),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_325),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_358),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_372),
.B(n_341),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_327),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_332),
.Y(n_394)
);

OA21x2_ASAP7_75t_L g395 ( 
.A1(n_349),
.A2(n_250),
.B(n_239),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_342),
.B(n_238),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_347),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_330),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_330),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_336),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_359),
.B(n_315),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_333),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_336),
.B(n_300),
.Y(n_403)
);

INVx4_ASAP7_75t_L g404 ( 
.A(n_328),
.Y(n_404)
);

AND2x6_ASAP7_75t_L g405 ( 
.A(n_358),
.B(n_234),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_371),
.B(n_300),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_329),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_377),
.Y(n_408)
);

OR2x2_ASAP7_75t_SL g409 ( 
.A(n_343),
.B(n_310),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_339),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_345),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_350),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_331),
.B(n_310),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_353),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_344),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_326),
.B(n_272),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_368),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_356),
.B(n_233),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_357),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_361),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_375),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_365),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_366),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_373),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_374),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_376),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_373),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_375),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_379),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_379),
.Y(n_430)
);

INVx4_ASAP7_75t_L g431 ( 
.A(n_324),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_324),
.B(n_271),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_368),
.B(n_233),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_370),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_370),
.B(n_297),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_335),
.B(n_323),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_399),
.B(n_280),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_408),
.Y(n_438)
);

OAI22xp33_ASAP7_75t_SL g439 ( 
.A1(n_401),
.A2(n_289),
.B1(n_292),
.B2(n_284),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_399),
.B(n_298),
.Y(n_440)
);

INVxp67_ASAP7_75t_SL g441 ( 
.A(n_399),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_398),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_398),
.Y(n_443)
);

BUFx10_ASAP7_75t_L g444 ( 
.A(n_432),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_408),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_399),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_398),
.Y(n_447)
);

AND2x6_ASAP7_75t_L g448 ( 
.A(n_410),
.B(n_234),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_395),
.B(n_305),
.Y(n_449)
);

INVx4_ASAP7_75t_L g450 ( 
.A(n_414),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_388),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_388),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_397),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_418),
.B(n_340),
.Y(n_454)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_414),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_395),
.B(n_308),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_414),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_395),
.B(n_313),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_397),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_395),
.B(n_322),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_397),
.Y(n_461)
);

BUFx8_ASAP7_75t_SL g462 ( 
.A(n_434),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_390),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_400),
.B(n_295),
.Y(n_464)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_414),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_436),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_408),
.B(n_352),
.Y(n_467)
);

OR2x6_ASAP7_75t_L g468 ( 
.A(n_431),
.B(n_234),
.Y(n_468)
);

BUFx10_ASAP7_75t_L g469 ( 
.A(n_432),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_400),
.B(n_268),
.Y(n_470)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_414),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_380),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_400),
.B(n_269),
.Y(n_473)
);

AND2x6_ASAP7_75t_L g474 ( 
.A(n_410),
.B(n_234),
.Y(n_474)
);

BUFx10_ASAP7_75t_L g475 ( 
.A(n_432),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_400),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_380),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_381),
.Y(n_478)
);

OAI22xp33_ASAP7_75t_L g479 ( 
.A1(n_401),
.A2(n_232),
.B1(n_248),
.B2(n_262),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_L g480 ( 
.A1(n_413),
.A2(n_304),
.B1(n_287),
.B2(n_288),
.Y(n_480)
);

BUFx10_ASAP7_75t_L g481 ( 
.A(n_432),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_386),
.Y(n_482)
);

AND3x4_ASAP7_75t_L g483 ( 
.A(n_429),
.B(n_367),
.C(n_355),
.Y(n_483)
);

AND2x4_ASAP7_75t_SL g484 ( 
.A(n_414),
.B(n_354),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_380),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_396),
.B(n_294),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_381),
.B(n_270),
.Y(n_487)
);

AND2x6_ASAP7_75t_L g488 ( 
.A(n_410),
.B(n_32),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_381),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_391),
.B(n_323),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_381),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_384),
.B(n_273),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_386),
.B(n_275),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_384),
.B(n_362),
.Y(n_494)
);

INVx4_ASAP7_75t_L g495 ( 
.A(n_420),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_418),
.B(n_363),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_386),
.B(n_276),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_390),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_393),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_382),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_393),
.Y(n_501)
);

INVxp67_ASAP7_75t_SL g502 ( 
.A(n_392),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_394),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_419),
.B(n_422),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_386),
.B(n_277),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_382),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_404),
.B(n_282),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_413),
.B(n_283),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_L g509 ( 
.A1(n_413),
.A2(n_301),
.B1(n_306),
.B2(n_319),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_394),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_396),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_502),
.B(n_420),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_463),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_511),
.B(n_504),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_438),
.B(n_415),
.Y(n_515)
);

AO22x2_ASAP7_75t_L g516 ( 
.A1(n_483),
.A2(n_429),
.B1(n_416),
.B2(n_430),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_498),
.Y(n_517)
);

AO22x2_ASAP7_75t_L g518 ( 
.A1(n_467),
.A2(n_429),
.B1(n_430),
.B2(n_407),
.Y(n_518)
);

NOR2xp67_ASAP7_75t_L g519 ( 
.A(n_457),
.B(n_404),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_499),
.B(n_403),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_511),
.A2(n_411),
.B1(n_412),
.B2(n_426),
.Y(n_521)
);

AO22x2_ASAP7_75t_L g522 ( 
.A1(n_486),
.A2(n_407),
.B1(n_436),
.B2(n_415),
.Y(n_522)
);

AO22x2_ASAP7_75t_L g523 ( 
.A1(n_494),
.A2(n_407),
.B1(n_435),
.B2(n_431),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_501),
.Y(n_524)
);

CKINVDCx14_ASAP7_75t_R g525 ( 
.A(n_466),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_503),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_438),
.B(n_406),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_454),
.A2(n_412),
.B1(n_411),
.B2(n_419),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_510),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_495),
.B(n_420),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_451),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_452),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_461),
.Y(n_533)
);

AO22x2_ASAP7_75t_L g534 ( 
.A1(n_445),
.A2(n_435),
.B1(n_431),
.B2(n_433),
.Y(n_534)
);

AO22x2_ASAP7_75t_L g535 ( 
.A1(n_464),
.A2(n_431),
.B1(n_433),
.B2(n_417),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_447),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_495),
.B(n_420),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_461),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_441),
.B(n_423),
.Y(n_539)
);

BUFx8_ASAP7_75t_L g540 ( 
.A(n_464),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_442),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_443),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_468),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_496),
.A2(n_411),
.B1(n_412),
.B2(n_422),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_468),
.Y(n_545)
);

NAND2x1p5_ASAP7_75t_L g546 ( 
.A(n_450),
.B(n_423),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_444),
.B(n_406),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_482),
.Y(n_548)
);

NAND2x1p5_ASAP7_75t_L g549 ( 
.A(n_450),
.B(n_423),
.Y(n_549)
);

AO22x2_ASAP7_75t_L g550 ( 
.A1(n_439),
.A2(n_417),
.B1(n_409),
.B2(n_413),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_479),
.A2(n_426),
.B1(n_425),
.B2(n_423),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_490),
.B(n_425),
.Y(n_552)
);

AO22x2_ASAP7_75t_L g553 ( 
.A1(n_439),
.A2(n_409),
.B1(n_427),
.B2(n_425),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_453),
.Y(n_554)
);

NAND2x1p5_ASAP7_75t_L g555 ( 
.A(n_455),
.B(n_465),
.Y(n_555)
);

AO22x2_ASAP7_75t_L g556 ( 
.A1(n_508),
.A2(n_427),
.B1(n_425),
.B2(n_404),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_480),
.B(n_421),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_470),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_482),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_470),
.A2(n_404),
.B1(n_392),
.B2(n_405),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_446),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_476),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_459),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_472),
.Y(n_564)
);

AO22x2_ASAP7_75t_L g565 ( 
.A1(n_508),
.A2(n_403),
.B1(n_424),
.B2(n_367),
.Y(n_565)
);

AO22x2_ASAP7_75t_L g566 ( 
.A1(n_492),
.A2(n_402),
.B1(n_428),
.B2(n_387),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_477),
.Y(n_567)
);

NAND2x1p5_ASAP7_75t_L g568 ( 
.A(n_455),
.B(n_402),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_484),
.B(n_383),
.Y(n_569)
);

OAI221xp5_ASAP7_75t_L g570 ( 
.A1(n_509),
.A2(n_383),
.B1(n_385),
.B2(n_387),
.C(n_382),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_485),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_473),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_500),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_506),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_444),
.B(n_428),
.Y(n_575)
);

AO22x2_ASAP7_75t_L g576 ( 
.A1(n_437),
.A2(n_428),
.B1(n_385),
.B2(n_5),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_478),
.B(n_405),
.Y(n_577)
);

AO22x2_ASAP7_75t_L g578 ( 
.A1(n_437),
.A2(n_428),
.B1(n_4),
.B2(n_6),
.Y(n_578)
);

AO22x2_ASAP7_75t_L g579 ( 
.A1(n_440),
.A2(n_428),
.B1(n_7),
.B2(n_8),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_488),
.A2(n_421),
.B1(n_428),
.B2(n_434),
.Y(n_580)
);

OAI221xp5_ASAP7_75t_L g581 ( 
.A1(n_449),
.A2(n_456),
.B1(n_458),
.B2(n_460),
.C(n_389),
.Y(n_581)
);

BUFx8_ASAP7_75t_L g582 ( 
.A(n_462),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_478),
.Y(n_583)
);

AO22x2_ASAP7_75t_L g584 ( 
.A1(n_440),
.A2(n_507),
.B1(n_449),
.B2(n_456),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_473),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_469),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_478),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_SL g588 ( 
.A1(n_488),
.A2(n_434),
.B1(n_405),
.B2(n_312),
.Y(n_588)
);

OR2x6_ASAP7_75t_L g589 ( 
.A(n_468),
.B(n_434),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_465),
.B(n_434),
.Y(n_590)
);

NAND2x1p5_ASAP7_75t_L g591 ( 
.A(n_471),
.B(n_389),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_471),
.B(n_469),
.Y(n_592)
);

OAI221xp5_ASAP7_75t_L g593 ( 
.A1(n_458),
.A2(n_389),
.B1(n_290),
.B2(n_314),
.C(n_321),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_475),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_489),
.B(n_405),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_489),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_514),
.B(n_475),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_SL g598 ( 
.A(n_575),
.B(n_434),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_528),
.B(n_481),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_544),
.B(n_481),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_527),
.B(n_493),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_519),
.B(n_493),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_521),
.B(n_497),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_551),
.B(n_547),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_512),
.B(n_497),
.Y(n_605)
);

AND2x2_ASAP7_75t_SL g606 ( 
.A(n_590),
.B(n_460),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_515),
.B(n_489),
.Y(n_607)
);

NAND2xp33_ASAP7_75t_SL g608 ( 
.A(n_545),
.B(n_505),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_552),
.B(n_505),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_558),
.B(n_488),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_572),
.B(n_491),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_585),
.B(n_488),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_569),
.B(n_491),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_580),
.B(n_491),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_560),
.B(n_487),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_520),
.B(n_487),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_513),
.B(n_517),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_524),
.B(n_293),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_539),
.B(n_448),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_SL g620 ( 
.A(n_543),
.B(n_299),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_526),
.B(n_302),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_529),
.B(n_303),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_531),
.B(n_307),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_583),
.B(n_448),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_532),
.B(n_448),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_594),
.B(n_309),
.Y(n_626)
);

NAND2xp33_ASAP7_75t_SL g627 ( 
.A(n_557),
.B(n_316),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_561),
.B(n_317),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_587),
.B(n_474),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_SL g630 ( 
.A(n_592),
.B(n_318),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_562),
.B(n_33),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_586),
.B(n_448),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_522),
.B(n_405),
.Y(n_633)
);

NAND2xp33_ASAP7_75t_SL g634 ( 
.A(n_530),
.B(n_474),
.Y(n_634)
);

NAND2xp33_ASAP7_75t_SL g635 ( 
.A(n_537),
.B(n_474),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_588),
.B(n_474),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_540),
.B(n_546),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_549),
.B(n_405),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_596),
.B(n_405),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_555),
.B(n_405),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_522),
.B(n_3),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_548),
.B(n_37),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_589),
.B(n_39),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_559),
.B(n_40),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_568),
.B(n_533),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_538),
.B(n_41),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_536),
.B(n_42),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_563),
.B(n_43),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_564),
.B(n_45),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_567),
.B(n_47),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_571),
.B(n_49),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_523),
.B(n_3),
.Y(n_652)
);

NAND2xp33_ASAP7_75t_SL g653 ( 
.A(n_577),
.B(n_7),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_574),
.B(n_51),
.Y(n_654)
);

NAND2xp33_ASAP7_75t_SL g655 ( 
.A(n_595),
.B(n_8),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_554),
.B(n_52),
.Y(n_656)
);

NAND2xp33_ASAP7_75t_SL g657 ( 
.A(n_589),
.B(n_9),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_573),
.B(n_55),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_541),
.B(n_56),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_581),
.B(n_9),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_542),
.B(n_58),
.Y(n_661)
);

AO21x2_ASAP7_75t_L g662 ( 
.A1(n_615),
.A2(n_593),
.B(n_570),
.Y(n_662)
);

NOR2xp67_ASAP7_75t_L g663 ( 
.A(n_626),
.B(n_59),
.Y(n_663)
);

AOI21x1_ASAP7_75t_SL g664 ( 
.A1(n_660),
.A2(n_556),
.B(n_553),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_601),
.B(n_553),
.Y(n_665)
);

OAI21x1_ASAP7_75t_L g666 ( 
.A1(n_624),
.A2(n_629),
.B(n_645),
.Y(n_666)
);

O2A1O1Ixp5_ASAP7_75t_L g667 ( 
.A1(n_609),
.A2(n_556),
.B(n_566),
.C(n_584),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_617),
.Y(n_668)
);

AND2x2_ASAP7_75t_SL g669 ( 
.A(n_643),
.B(n_582),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_607),
.A2(n_550),
.B1(n_579),
.B2(n_578),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_597),
.B(n_523),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_616),
.B(n_550),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_613),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_606),
.B(n_566),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_606),
.B(n_518),
.Y(n_675)
);

NOR2x1_ASAP7_75t_L g676 ( 
.A(n_604),
.B(n_525),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_603),
.B(n_584),
.Y(n_677)
);

AO31x2_ASAP7_75t_L g678 ( 
.A1(n_619),
.A2(n_576),
.A3(n_518),
.B(n_534),
.Y(n_678)
);

NAND3xp33_ASAP7_75t_SL g679 ( 
.A(n_627),
.B(n_535),
.C(n_534),
.Y(n_679)
);

AOI221x1_ASAP7_75t_L g680 ( 
.A1(n_653),
.A2(n_565),
.B1(n_576),
.B2(n_516),
.C(n_535),
.Y(n_680)
);

AOI221x1_ASAP7_75t_L g681 ( 
.A1(n_655),
.A2(n_565),
.B1(n_516),
.B2(n_578),
.C(n_579),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_602),
.A2(n_591),
.B(n_127),
.Y(n_682)
);

NAND2xp33_ASAP7_75t_L g683 ( 
.A(n_608),
.B(n_63),
.Y(n_683)
);

OAI21x1_ASAP7_75t_L g684 ( 
.A1(n_605),
.A2(n_126),
.B(n_225),
.Y(n_684)
);

OAI21x1_ASAP7_75t_L g685 ( 
.A1(n_611),
.A2(n_124),
.B(n_224),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_643),
.B(n_64),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_652),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_614),
.A2(n_610),
.B1(n_612),
.B2(n_600),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_631),
.Y(n_689)
);

AND2x2_ASAP7_75t_SL g690 ( 
.A(n_641),
.B(n_10),
.Y(n_690)
);

O2A1O1Ixp33_ASAP7_75t_SL g691 ( 
.A1(n_647),
.A2(n_130),
.B(n_222),
.C(n_221),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_599),
.B(n_10),
.Y(n_692)
);

OAI21x1_ASAP7_75t_L g693 ( 
.A1(n_636),
.A2(n_122),
.B(n_220),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_631),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_634),
.A2(n_121),
.B(n_219),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_612),
.B(n_65),
.Y(n_696)
);

OAI22xp5_ASAP7_75t_L g697 ( 
.A1(n_610),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_697)
);

OAI22xp5_ASAP7_75t_L g698 ( 
.A1(n_633),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_625),
.Y(n_699)
);

OAI21xp5_ASAP7_75t_L g700 ( 
.A1(n_639),
.A2(n_133),
.B(n_218),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_618),
.B(n_15),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_635),
.A2(n_132),
.B(n_217),
.Y(n_702)
);

OAI21x1_ASAP7_75t_L g703 ( 
.A1(n_638),
.A2(n_119),
.B(n_216),
.Y(n_703)
);

AO32x2_ASAP7_75t_L g704 ( 
.A1(n_657),
.A2(n_16),
.A3(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_704)
);

BUFx2_ASAP7_75t_L g705 ( 
.A(n_620),
.Y(n_705)
);

OAI21x1_ASAP7_75t_L g706 ( 
.A1(n_640),
.A2(n_135),
.B(n_214),
.Y(n_706)
);

INVx3_ASAP7_75t_SL g707 ( 
.A(n_637),
.Y(n_707)
);

AO31x2_ASAP7_75t_L g708 ( 
.A1(n_598),
.A2(n_19),
.A3(n_22),
.B(n_23),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_621),
.A2(n_137),
.B(n_209),
.Y(n_709)
);

OAI21x1_ASAP7_75t_SL g710 ( 
.A1(n_642),
.A2(n_644),
.B(n_659),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_632),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_622),
.B(n_67),
.Y(n_712)
);

AO31x2_ASAP7_75t_L g713 ( 
.A1(n_648),
.A2(n_24),
.A3(n_25),
.B(n_26),
.Y(n_713)
);

AOI22x1_ASAP7_75t_L g714 ( 
.A1(n_649),
.A2(n_138),
.B1(n_206),
.B2(n_202),
.Y(n_714)
);

O2A1O1Ixp5_ASAP7_75t_L g715 ( 
.A1(n_623),
.A2(n_136),
.B(n_198),
.C(n_197),
.Y(n_715)
);

OAI21xp5_ASAP7_75t_L g716 ( 
.A1(n_650),
.A2(n_226),
.B(n_116),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_646),
.Y(n_717)
);

AO21x2_ASAP7_75t_L g718 ( 
.A1(n_677),
.A2(n_661),
.B(n_654),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_668),
.Y(n_719)
);

OR2x6_ASAP7_75t_L g720 ( 
.A(n_689),
.B(n_651),
.Y(n_720)
);

OAI21x1_ASAP7_75t_L g721 ( 
.A1(n_666),
.A2(n_658),
.B(n_656),
.Y(n_721)
);

BUFx2_ASAP7_75t_L g722 ( 
.A(n_687),
.Y(n_722)
);

AO21x2_ASAP7_75t_L g723 ( 
.A1(n_677),
.A2(n_628),
.B(n_630),
.Y(n_723)
);

OAI21x1_ASAP7_75t_L g724 ( 
.A1(n_693),
.A2(n_113),
.B(n_195),
.Y(n_724)
);

AO21x2_ASAP7_75t_L g725 ( 
.A1(n_679),
.A2(n_112),
.B(n_194),
.Y(n_725)
);

OAI21xp5_ASAP7_75t_L g726 ( 
.A1(n_667),
.A2(n_196),
.B(n_111),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_676),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_727)
);

AOI221xp5_ASAP7_75t_L g728 ( 
.A1(n_692),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.C(n_68),
.Y(n_728)
);

INVx8_ASAP7_75t_L g729 ( 
.A(n_671),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_690),
.A2(n_29),
.B1(n_30),
.B2(n_69),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_699),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_672),
.A2(n_71),
.B1(n_72),
.B2(n_75),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_673),
.Y(n_733)
);

BUFx4f_ASAP7_75t_SL g734 ( 
.A(n_707),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_665),
.B(n_694),
.Y(n_735)
);

OAI21x1_ASAP7_75t_L g736 ( 
.A1(n_684),
.A2(n_76),
.B(n_77),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_711),
.Y(n_737)
);

OAI21x1_ASAP7_75t_L g738 ( 
.A1(n_685),
.A2(n_78),
.B(n_80),
.Y(n_738)
);

OAI211xp5_ASAP7_75t_L g739 ( 
.A1(n_680),
.A2(n_81),
.B(n_82),
.C(n_83),
.Y(n_739)
);

AO21x2_ASAP7_75t_L g740 ( 
.A1(n_674),
.A2(n_84),
.B(n_85),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_SL g741 ( 
.A(n_669),
.B(n_698),
.Y(n_741)
);

OR2x6_ASAP7_75t_L g742 ( 
.A(n_688),
.B(n_86),
.Y(n_742)
);

BUFx4f_ASAP7_75t_L g743 ( 
.A(n_705),
.Y(n_743)
);

OAI21x1_ASAP7_75t_L g744 ( 
.A1(n_706),
.A2(n_89),
.B(n_91),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_675),
.Y(n_745)
);

INVx4_ASAP7_75t_L g746 ( 
.A(n_717),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_696),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_670),
.B(n_92),
.Y(n_748)
);

O2A1O1Ixp5_ASAP7_75t_L g749 ( 
.A1(n_670),
.A2(n_94),
.B(n_96),
.C(n_97),
.Y(n_749)
);

OAI21x1_ASAP7_75t_L g750 ( 
.A1(n_682),
.A2(n_98),
.B(n_99),
.Y(n_750)
);

OR2x6_ASAP7_75t_L g751 ( 
.A(n_688),
.B(n_686),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_696),
.B(n_192),
.Y(n_752)
);

INVx1_ASAP7_75t_SL g753 ( 
.A(n_701),
.Y(n_753)
);

O2A1O1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_698),
.A2(n_101),
.B(n_102),
.C(n_104),
.Y(n_754)
);

OR2x2_ASAP7_75t_L g755 ( 
.A(n_678),
.B(n_105),
.Y(n_755)
);

OAI21x1_ASAP7_75t_L g756 ( 
.A1(n_703),
.A2(n_107),
.B(n_108),
.Y(n_756)
);

OR2x2_ASAP7_75t_L g757 ( 
.A(n_678),
.B(n_118),
.Y(n_757)
);

O2A1O1Ixp33_ASAP7_75t_SL g758 ( 
.A1(n_712),
.A2(n_139),
.B(n_140),
.C(n_141),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_662),
.A2(n_146),
.B(n_148),
.Y(n_759)
);

OAI21x1_ASAP7_75t_L g760 ( 
.A1(n_664),
.A2(n_710),
.B(n_695),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_683),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_678),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_713),
.Y(n_763)
);

NAND3xp33_ASAP7_75t_L g764 ( 
.A(n_681),
.B(n_149),
.C(n_153),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_697),
.B(n_156),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_704),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_704),
.Y(n_767)
);

OAI21x1_ASAP7_75t_L g768 ( 
.A1(n_702),
.A2(n_715),
.B(n_716),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_SL g769 ( 
.A(n_697),
.B(n_157),
.Y(n_769)
);

OA21x2_ASAP7_75t_L g770 ( 
.A1(n_716),
.A2(n_158),
.B(n_159),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_662),
.B(n_160),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_743),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_762),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_745),
.B(n_747),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_763),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_743),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_760),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_771),
.Y(n_778)
);

INVx1_ASAP7_75t_SL g779 ( 
.A(n_722),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_771),
.Y(n_780)
);

OA21x2_ASAP7_75t_L g781 ( 
.A1(n_749),
.A2(n_700),
.B(n_709),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_SL g782 ( 
.A1(n_741),
.A2(n_714),
.B1(n_700),
.B2(n_704),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_741),
.B(n_663),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_766),
.Y(n_784)
);

CKINVDCx16_ASAP7_75t_R g785 ( 
.A(n_769),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_753),
.B(n_691),
.Y(n_786)
);

INVx3_ASAP7_75t_L g787 ( 
.A(n_736),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_744),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_737),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_753),
.B(n_161),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_765),
.B(n_731),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_767),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_735),
.B(n_166),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_729),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_756),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_719),
.Y(n_796)
);

BUFx2_ASAP7_75t_L g797 ( 
.A(n_742),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_729),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_721),
.Y(n_799)
);

INVxp33_ASAP7_75t_L g800 ( 
.A(n_733),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_755),
.Y(n_801)
);

INVx3_ASAP7_75t_L g802 ( 
.A(n_724),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_751),
.B(n_713),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_757),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_740),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_770),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_751),
.B(n_713),
.Y(n_807)
);

A2O1A1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_726),
.A2(n_754),
.B(n_769),
.C(n_761),
.Y(n_808)
);

AOI21x1_ASAP7_75t_L g809 ( 
.A1(n_759),
.A2(n_708),
.B(n_168),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_729),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_770),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_734),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_740),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_725),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_718),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_738),
.Y(n_816)
);

OA21x2_ASAP7_75t_L g817 ( 
.A1(n_749),
.A2(n_726),
.B(n_768),
.Y(n_817)
);

INVx1_ASAP7_75t_SL g818 ( 
.A(n_734),
.Y(n_818)
);

AOI221xp5_ASAP7_75t_L g819 ( 
.A1(n_728),
.A2(n_708),
.B1(n_169),
.B2(n_172),
.C(n_173),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_725),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_748),
.B(n_708),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_718),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_748),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_751),
.Y(n_824)
);

INVx4_ASAP7_75t_R g825 ( 
.A(n_761),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_742),
.Y(n_826)
);

OAI21x1_ASAP7_75t_L g827 ( 
.A1(n_750),
.A2(n_167),
.B(n_174),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_746),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_746),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_796),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_774),
.B(n_730),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_796),
.Y(n_832)
);

XOR2xp5_ASAP7_75t_L g833 ( 
.A(n_810),
.B(n_727),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_R g834 ( 
.A(n_829),
.B(n_752),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_796),
.Y(n_835)
);

XNOR2xp5_ASAP7_75t_L g836 ( 
.A(n_818),
.B(n_728),
.Y(n_836)
);

XNOR2xp5_ASAP7_75t_L g837 ( 
.A(n_818),
.B(n_752),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_794),
.B(n_742),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_774),
.B(n_791),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_779),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_773),
.Y(n_841)
);

NAND2xp33_ASAP7_75t_R g842 ( 
.A(n_783),
.B(n_720),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_791),
.B(n_723),
.Y(n_843)
);

BUFx10_ASAP7_75t_L g844 ( 
.A(n_812),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_R g845 ( 
.A(n_772),
.B(n_732),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_789),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_823),
.B(n_723),
.Y(n_847)
);

OR2x4_ASAP7_75t_L g848 ( 
.A(n_790),
.B(n_720),
.Y(n_848)
);

OR2x6_ASAP7_75t_L g849 ( 
.A(n_772),
.B(n_776),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_794),
.B(n_720),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_798),
.B(n_764),
.Y(n_851)
);

BUFx2_ASAP7_75t_L g852 ( 
.A(n_776),
.Y(n_852)
);

NAND2xp33_ASAP7_75t_R g853 ( 
.A(n_797),
.B(n_793),
.Y(n_853)
);

NAND2xp33_ASAP7_75t_R g854 ( 
.A(n_797),
.B(n_759),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_773),
.Y(n_855)
);

NAND2xp33_ASAP7_75t_R g856 ( 
.A(n_826),
.B(n_175),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_800),
.B(n_754),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_773),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_R g859 ( 
.A(n_812),
.B(n_177),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_823),
.B(n_739),
.Y(n_860)
);

NAND2xp33_ASAP7_75t_R g861 ( 
.A(n_826),
.B(n_807),
.Y(n_861)
);

BUFx10_ASAP7_75t_L g862 ( 
.A(n_828),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_798),
.B(n_178),
.Y(n_863)
);

NAND2xp33_ASAP7_75t_SL g864 ( 
.A(n_785),
.B(n_739),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_785),
.B(n_180),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_779),
.B(n_789),
.Y(n_866)
);

NAND2xp33_ASAP7_75t_R g867 ( 
.A(n_826),
.B(n_183),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_789),
.B(n_758),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_R g869 ( 
.A(n_801),
.B(n_185),
.Y(n_869)
);

NAND2xp33_ASAP7_75t_R g870 ( 
.A(n_803),
.B(n_807),
.Y(n_870)
);

NAND2xp33_ASAP7_75t_SL g871 ( 
.A(n_825),
.B(n_186),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_824),
.B(n_187),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_784),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_801),
.B(n_188),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_804),
.B(n_190),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_848),
.B(n_824),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_873),
.B(n_803),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_841),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_855),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_858),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_832),
.B(n_784),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_866),
.B(n_804),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_840),
.B(n_780),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_835),
.B(n_792),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_839),
.B(n_780),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_830),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_843),
.B(n_792),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_SL g888 ( 
.A1(n_869),
.A2(n_824),
.B1(n_781),
.B2(n_821),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_846),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_847),
.B(n_780),
.Y(n_890)
);

INVxp67_ASAP7_75t_L g891 ( 
.A(n_852),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_857),
.B(n_778),
.Y(n_892)
);

OAI22xp5_ASAP7_75t_L g893 ( 
.A1(n_836),
.A2(n_808),
.B1(n_782),
.B2(n_819),
.Y(n_893)
);

AND2x4_ASAP7_75t_SL g894 ( 
.A(n_862),
.B(n_775),
.Y(n_894)
);

INVxp67_ASAP7_75t_SL g895 ( 
.A(n_860),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_838),
.B(n_777),
.Y(n_896)
);

BUFx2_ASAP7_75t_L g897 ( 
.A(n_838),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_874),
.B(n_778),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_850),
.B(n_777),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_868),
.Y(n_900)
);

OR2x2_ASAP7_75t_L g901 ( 
.A(n_831),
.B(n_778),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_850),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_851),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_875),
.Y(n_904)
);

OR2x2_ASAP7_75t_L g905 ( 
.A(n_849),
.B(n_815),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_872),
.B(n_777),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_853),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_872),
.B(n_775),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_864),
.A2(n_786),
.B1(n_821),
.B2(n_781),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_865),
.B(n_775),
.Y(n_910)
);

NOR2x1p5_ASAP7_75t_L g911 ( 
.A(n_851),
.B(n_820),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_877),
.B(n_822),
.Y(n_912)
);

OR2x2_ASAP7_75t_L g913 ( 
.A(n_892),
.B(n_813),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_895),
.B(n_822),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_878),
.Y(n_915)
);

AOI221xp5_ASAP7_75t_L g916 ( 
.A1(n_893),
.A2(n_833),
.B1(n_871),
.B2(n_859),
.C(n_834),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_877),
.B(n_815),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_894),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_880),
.Y(n_919)
);

AND2x4_ASAP7_75t_SL g920 ( 
.A(n_907),
.B(n_862),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_880),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_883),
.B(n_822),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_878),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_887),
.B(n_815),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_887),
.B(n_820),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_879),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_911),
.B(n_799),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_890),
.B(n_814),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_879),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_900),
.B(n_814),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_876),
.B(n_844),
.Y(n_931)
);

OAI211xp5_ASAP7_75t_SL g932 ( 
.A1(n_891),
.A2(n_813),
.B(n_805),
.C(n_842),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_919),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_927),
.B(n_911),
.Y(n_934)
);

OR2x2_ASAP7_75t_L g935 ( 
.A(n_913),
.B(n_890),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_919),
.Y(n_936)
);

INVxp67_ASAP7_75t_SL g937 ( 
.A(n_930),
.Y(n_937)
);

INVx1_ASAP7_75t_SL g938 ( 
.A(n_920),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_928),
.B(n_897),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_915),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_921),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_928),
.B(n_897),
.Y(n_942)
);

OR2x2_ASAP7_75t_L g943 ( 
.A(n_913),
.B(n_905),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_921),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_915),
.Y(n_945)
);

INVx2_ASAP7_75t_SL g946 ( 
.A(n_918),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_925),
.B(n_900),
.Y(n_947)
);

OAI22xp33_ASAP7_75t_L g948 ( 
.A1(n_938),
.A2(n_856),
.B1(n_867),
.B2(n_870),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_937),
.B(n_947),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_935),
.B(n_931),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_943),
.B(n_925),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_943),
.B(n_935),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_934),
.A2(n_916),
.B1(n_854),
.B2(n_932),
.Y(n_953)
);

NOR2x1_ASAP7_75t_L g954 ( 
.A(n_940),
.B(n_918),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_939),
.B(n_920),
.Y(n_955)
);

BUFx2_ASAP7_75t_L g956 ( 
.A(n_954),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_950),
.B(n_934),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_952),
.B(n_934),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_951),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_949),
.Y(n_960)
);

AND2x4_ASAP7_75t_SL g961 ( 
.A(n_953),
.B(n_844),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_948),
.A2(n_888),
.B1(n_909),
.B2(n_903),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_955),
.B(n_941),
.Y(n_963)
);

OA211x2_ASAP7_75t_L g964 ( 
.A1(n_963),
.A2(n_914),
.B(n_910),
.C(n_922),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_963),
.Y(n_965)
);

AOI211xp5_ASAP7_75t_L g966 ( 
.A1(n_962),
.A2(n_837),
.B(n_946),
.C(n_845),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_960),
.B(n_942),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_959),
.B(n_942),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_965),
.B(n_957),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_966),
.B(n_958),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_967),
.B(n_961),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_968),
.B(n_956),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_969),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_972),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_971),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_970),
.Y(n_976)
);

BUFx2_ASAP7_75t_L g977 ( 
.A(n_969),
.Y(n_977)
);

AOI211xp5_ASAP7_75t_L g978 ( 
.A1(n_976),
.A2(n_962),
.B(n_863),
.C(n_946),
.Y(n_978)
);

NAND4xp75_ASAP7_75t_L g979 ( 
.A(n_974),
.B(n_964),
.C(n_825),
.D(n_939),
.Y(n_979)
);

NAND4xp75_ASAP7_75t_L g980 ( 
.A(n_975),
.B(n_781),
.C(n_944),
.D(n_936),
.Y(n_980)
);

NAND4xp25_ASAP7_75t_L g981 ( 
.A(n_975),
.B(n_863),
.C(n_861),
.D(n_904),
.Y(n_981)
);

NOR3xp33_ASAP7_75t_L g982 ( 
.A(n_973),
.B(n_904),
.C(n_903),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_977),
.B(n_933),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_977),
.B(n_945),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_L g985 ( 
.A1(n_976),
.A2(n_902),
.B1(n_901),
.B2(n_908),
.Y(n_985)
);

XNOR2x1_ASAP7_75t_L g986 ( 
.A(n_979),
.B(n_980),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_983),
.Y(n_987)
);

AOI221xp5_ASAP7_75t_L g988 ( 
.A1(n_978),
.A2(n_945),
.B1(n_940),
.B2(n_902),
.C(n_923),
.Y(n_988)
);

NOR3xp33_ASAP7_75t_SL g989 ( 
.A(n_984),
.B(n_981),
.C(n_985),
.Y(n_989)
);

NOR3xp33_ASAP7_75t_L g990 ( 
.A(n_982),
.B(n_901),
.C(n_827),
.Y(n_990)
);

AOI221xp5_ASAP7_75t_L g991 ( 
.A1(n_983),
.A2(n_923),
.B1(n_894),
.B2(n_882),
.C(n_926),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_978),
.A2(n_927),
.B1(n_849),
.B2(n_926),
.Y(n_992)
);

OAI221xp5_ASAP7_75t_L g993 ( 
.A1(n_978),
.A2(n_885),
.B1(n_929),
.B2(n_905),
.C(n_781),
.Y(n_993)
);

NOR2x1_ASAP7_75t_L g994 ( 
.A(n_987),
.B(n_929),
.Y(n_994)
);

XNOR2x1_ASAP7_75t_L g995 ( 
.A(n_986),
.B(n_191),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_992),
.B(n_927),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_989),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_990),
.B(n_991),
.Y(n_998)
);

NAND4xp75_ASAP7_75t_L g999 ( 
.A(n_988),
.B(n_805),
.C(n_817),
.D(n_924),
.Y(n_999)
);

AOI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_993),
.A2(n_924),
.B1(n_899),
.B2(n_896),
.Y(n_1000)
);

AOI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_986),
.A2(n_899),
.B1(n_896),
.B2(n_898),
.Y(n_1001)
);

NOR2x1_ASAP7_75t_L g1002 ( 
.A(n_987),
.B(n_886),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_997),
.B(n_917),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_1002),
.B(n_899),
.Y(n_1004)
);

XOR2x2_ASAP7_75t_L g1005 ( 
.A(n_995),
.B(n_809),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_R g1006 ( 
.A(n_998),
.B(n_809),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_R g1007 ( 
.A(n_996),
.B(n_908),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_994),
.B(n_917),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_R g1009 ( 
.A(n_999),
.B(n_898),
.Y(n_1009)
);

NAND2xp33_ASAP7_75t_SL g1010 ( 
.A(n_1001),
.B(n_1000),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_997),
.B(n_899),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_1003),
.Y(n_1012)
);

OA22x2_ASAP7_75t_L g1013 ( 
.A1(n_1011),
.A2(n_896),
.B1(n_886),
.B2(n_889),
.Y(n_1013)
);

INVxp67_ASAP7_75t_L g1014 ( 
.A(n_1010),
.Y(n_1014)
);

INVxp67_ASAP7_75t_L g1015 ( 
.A(n_1005),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_1008),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_1004),
.Y(n_1017)
);

XNOR2xp5_ASAP7_75t_L g1018 ( 
.A(n_1007),
.B(n_827),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_1009),
.A2(n_896),
.B1(n_889),
.B2(n_906),
.Y(n_1019)
);

AO21x2_ASAP7_75t_L g1020 ( 
.A1(n_1014),
.A2(n_1006),
.B(n_811),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_1017),
.A2(n_906),
.B1(n_817),
.B2(n_912),
.Y(n_1021)
);

OA21x2_ASAP7_75t_L g1022 ( 
.A1(n_1015),
.A2(n_811),
.B(n_806),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_1013),
.Y(n_1023)
);

INVxp67_ASAP7_75t_L g1024 ( 
.A(n_1023),
.Y(n_1024)
);

OAI22xp33_ASAP7_75t_SL g1025 ( 
.A1(n_1020),
.A2(n_1016),
.B1(n_1012),
.B2(n_1019),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_SL g1026 ( 
.A1(n_1020),
.A2(n_1018),
.B(n_817),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_1021),
.B(n_884),
.Y(n_1027)
);

AOI22xp33_ASAP7_75t_L g1028 ( 
.A1(n_1024),
.A2(n_1022),
.B1(n_906),
.B2(n_817),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_L g1029 ( 
.A1(n_1027),
.A2(n_1022),
.B1(n_906),
.B2(n_912),
.Y(n_1029)
);

OAI322xp33_ASAP7_75t_L g1030 ( 
.A1(n_1028),
.A2(n_1026),
.A3(n_1025),
.B1(n_811),
.B2(n_806),
.C1(n_802),
.C2(n_816),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_1029),
.B(n_787),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1030),
.Y(n_1032)
);

OA22x2_ASAP7_75t_L g1033 ( 
.A1(n_1031),
.A2(n_884),
.B1(n_881),
.B2(n_806),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1032),
.Y(n_1034)
);

BUFx4_ASAP7_75t_R g1035 ( 
.A(n_1033),
.Y(n_1035)
);

AOI221xp5_ASAP7_75t_L g1036 ( 
.A1(n_1034),
.A2(n_787),
.B1(n_788),
.B2(n_795),
.C(n_802),
.Y(n_1036)
);

OAI221xp5_ASAP7_75t_R g1037 ( 
.A1(n_1035),
.A2(n_881),
.B1(n_788),
.B2(n_795),
.C(n_802),
.Y(n_1037)
);

AOI211xp5_ASAP7_75t_L g1038 ( 
.A1(n_1036),
.A2(n_1037),
.B(n_799),
.C(n_795),
.Y(n_1038)
);


endmodule