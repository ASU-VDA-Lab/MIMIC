module fake_jpeg_19848_n_176 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_176);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_8),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_48),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_35),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_12),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_4),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_0),
.Y(n_74)
);

BUFx16f_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_7),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_73),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_84),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

BUFx12f_ASAP7_75t_SL g85 ( 
.A(n_61),
.Y(n_85)
);

BUFx4f_ASAP7_75t_SL g97 ( 
.A(n_85),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_85),
.A2(n_50),
.B1(n_77),
.B2(n_67),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_87),
.A2(n_98),
.B1(n_61),
.B2(n_72),
.Y(n_109)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_77),
.B1(n_66),
.B2(n_62),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_96),
.A2(n_70),
.B1(n_58),
.B2(n_64),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_101),
.A2(n_107),
.B1(n_72),
.B2(n_69),
.Y(n_120)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_108),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_L g103 ( 
.A1(n_96),
.A2(n_54),
.B(n_56),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_75),
.C(n_55),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_76),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_0),
.Y(n_127)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_95),
.A2(n_65),
.B1(n_69),
.B2(n_31),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_91),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_111),
.B(n_60),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_75),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_120),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_121),
.B(n_127),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

AO21x1_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_128),
.B(n_2),
.Y(n_142)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_110),
.A2(n_60),
.B1(n_52),
.B2(n_59),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_125),
.A2(n_112),
.B(n_100),
.C(n_74),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_101),
.A2(n_52),
.B1(n_71),
.B2(n_68),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_126),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_1),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_119),
.A2(n_114),
.B(n_113),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_130),
.A2(n_141),
.B(n_133),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_118),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_136),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_133),
.A2(n_119),
.B1(n_5),
.B2(n_6),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_134),
.Y(n_148)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_142),
.Y(n_144)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_139),
.B(n_129),
.Y(n_143)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_146),
.A2(n_153),
.B1(n_140),
.B2(n_14),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_135),
.B(n_3),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_150),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_141),
.A2(n_23),
.B(n_47),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_21),
.Y(n_151)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_148),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_158),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_148),
.A2(n_13),
.B1(n_15),
.B2(n_17),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_153),
.C(n_144),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_154),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_161),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_162),
.A2(n_157),
.B1(n_156),
.B2(n_145),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_160),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_165),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_163),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_149),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_159),
.Y(n_169)
);

NOR2x1_ASAP7_75t_SL g170 ( 
.A(n_169),
.B(n_18),
.Y(n_170)
);

OAI211xp5_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_19),
.B(n_20),
.C(n_24),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_25),
.C(n_26),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_33),
.B(n_34),
.Y(n_173)
);

BUFx24_ASAP7_75t_SL g174 ( 
.A(n_173),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_174),
.A2(n_38),
.B(n_39),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_41),
.C(n_46),
.Y(n_176)
);


endmodule