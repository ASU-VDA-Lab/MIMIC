module real_jpeg_5903_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_0),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_0),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_0),
.B(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_SL g233 ( 
.A(n_0),
.B(n_234),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_0),
.B(n_249),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_0),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_0),
.B(n_266),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_0),
.B(n_442),
.Y(n_441)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_1),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_1),
.Y(n_275)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_1),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_1),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_1),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_2),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_2),
.Y(n_104)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_2),
.Y(n_125)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_2),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_2),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_3),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_3),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_3),
.B(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_3),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_3),
.B(n_58),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_3),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_3),
.B(n_51),
.Y(n_363)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_4),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_4),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_4),
.B(n_211),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g236 ( 
.A(n_4),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_4),
.B(n_413),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_5),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_5),
.B(n_223),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_5),
.B(n_246),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_5),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_5),
.B(n_323),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_5),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_5),
.B(n_303),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_5),
.B(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_6),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_6),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_6),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_6),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_6),
.B(n_211),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_6),
.B(n_404),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_6),
.B(n_329),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_7),
.Y(n_101)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_7),
.Y(n_116)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_7),
.Y(n_140)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_8),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_9),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_9),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_9),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_9),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_9),
.B(n_171),
.Y(n_170)
);

AND2x2_ASAP7_75t_SL g400 ( 
.A(n_9),
.B(n_401),
.Y(n_400)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_10),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g329 ( 
.A(n_10),
.Y(n_329)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_12),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_12),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_12),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_13),
.B(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_13),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_13),
.B(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_13),
.B(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_13),
.B(n_130),
.Y(n_129)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_15),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_49),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_16),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_16),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_16),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_16),
.B(n_181),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_16),
.B(n_273),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_16),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_16),
.B(n_329),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_17),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_17),
.B(n_190),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_17),
.B(n_252),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_17),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_17),
.B(n_301),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_17),
.B(n_311),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_17),
.B(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_17),
.B(n_257),
.Y(n_424)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_19),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_19),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_19),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_19),
.B(n_321),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_19),
.B(n_329),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_19),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_19),
.B(n_231),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_491),
.B(n_494),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_192),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_191),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_153),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_25),
.B(n_153),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_110),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_78),
.C(n_91),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_27),
.B(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_47),
.C(n_60),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_28),
.B(n_47),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_33),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_29),
.B(n_39),
.C(n_46),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_30),
.B(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_30),
.B(n_269),
.Y(n_268)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_32),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_39),
.B1(n_40),
.B2(n_46),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx8_ASAP7_75t_L g266 ( 
.A(n_36),
.Y(n_266)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_38),
.Y(n_131)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_38),
.Y(n_187)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_38),
.Y(n_247)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_44),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_44),
.Y(n_361)
);

INVx6_ASAP7_75t_L g415 ( 
.A(n_44),
.Y(n_415)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_45),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g235 ( 
.A(n_45),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_45),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_47),
.B(n_162),
.C(n_165),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_47),
.B(n_165),
.Y(n_464)
);

FAx1_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_52),
.CI(n_55),
.CON(n_47),
.SN(n_47)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_59),
.Y(n_250)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_59),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_60),
.B(n_483),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_66),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_61),
.B(n_67),
.C(n_77),
.Y(n_151)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_63),
.Y(n_215)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_65),
.Y(n_225)
);

INVx6_ASAP7_75t_L g445 ( 
.A(n_65),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_71),
.B2(n_77),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_114),
.C(n_117),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_67),
.A2(n_68),
.B1(n_117),
.B2(n_118),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_94),
.C(n_98),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_71),
.A2(n_77),
.B1(n_94),
.B2(n_95),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_76),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_76),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_78),
.A2(n_91),
.B1(n_92),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_78),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_79),
.B(n_83),
.C(n_86),
.Y(n_136)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_102),
.C(n_105),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_93),
.B(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_94),
.B(n_166),
.C(n_170),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_94),
.A2(n_95),
.B1(n_170),
.B2(n_455),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_97),
.Y(n_213)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_97),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_98),
.B(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_101),
.Y(n_218)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_101),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_102),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.Y(n_174)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_105),
.A2(n_106),
.B1(n_188),
.B2(n_189),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_106),
.B(n_176),
.C(n_188),
.Y(n_175)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_109),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_148),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_135),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_121),
.B1(n_133),
.B2(n_134),
.Y(n_112)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_118),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx5_ASAP7_75t_L g333 ( 
.A(n_120),
.Y(n_333)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_126),
.B1(n_127),
.B2(n_132),
.Y(n_121)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_125),
.Y(n_231)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_141),
.B1(n_142),
.B2(n_147),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_138),
.Y(n_147)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.C(n_152),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_152),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.C(n_159),
.Y(n_153)
);

FAx1_ASAP7_75t_SL g487 ( 
.A(n_154),
.B(n_157),
.CI(n_159),
.CON(n_487),
.SN(n_487)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_173),
.C(n_175),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_160),
.A2(n_161),
.B1(n_480),
.B2(n_481),
.Y(n_479)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_162),
.A2(n_163),
.B1(n_464),
.B2(n_465),
.Y(n_463)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_166),
.A2(n_167),
.B1(n_453),
.B2(n_454),
.Y(n_452)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_170),
.Y(n_455)
);

BUFx5_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_172),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_173),
.B(n_175),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_177),
.B(n_472),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.C(n_184),
.Y(n_177)
);

FAx1_ASAP7_75t_SL g449 ( 
.A(n_178),
.B(n_180),
.CI(n_184),
.CON(n_449),
.SN(n_449)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_183),
.Y(n_252)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

AO21x1_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_486),
.B(n_489),
.Y(n_192)
);

OAI21x1_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_476),
.B(n_485),
.Y(n_193)
);

AOI21x1_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_459),
.B(n_475),
.Y(n_194)
);

OAI21x1_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_428),
.B(n_458),
.Y(n_195)
);

AOI21x1_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_390),
.B(n_427),
.Y(n_196)
);

AO21x1_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_314),
.B(n_389),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_294),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_199),
.B(n_294),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_242),
.B2(n_293),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_200),
.B(n_243),
.C(n_276),
.Y(n_426)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_219),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_202),
.B(n_220),
.C(n_241),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_214),
.C(n_216),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_203),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_209),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_204),
.A2(n_205),
.B1(n_209),
.B2(n_210),
.Y(n_299)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_214),
.B(n_216),
.Y(n_313)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_227),
.B1(n_240),
.B2(n_241),
.Y(n_219)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_220),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B(n_226),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_222),
.Y(n_226)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g405 ( 
.A(n_226),
.B(n_406),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_226),
.B(n_395),
.C(n_406),
.Y(n_435)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_232),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_228),
.B(n_233),
.C(n_236),
.Y(n_425)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx5_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_242),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_276),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_253),
.C(n_267),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_244),
.B(n_296),
.Y(n_295)
);

BUFx24_ASAP7_75t_SL g498 ( 
.A(n_244),
.Y(n_498)
);

FAx1_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_248),
.CI(n_251),
.CON(n_244),
.SN(n_244)
);

MAJx2_ASAP7_75t_L g292 ( 
.A(n_245),
.B(n_248),
.C(n_251),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_247),
.Y(n_279)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_253),
.A2(n_254),
.B1(n_267),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

MAJx2_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_259),
.C(n_264),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_255),
.A2(n_256),
.B1(n_264),
.B2(n_265),
.Y(n_382)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_259),
.B(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_267),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_272),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_272),
.Y(n_291)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx8_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

BUFx5_ASAP7_75t_L g311 ( 
.A(n_271),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_271),
.Y(n_404)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_275),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_290),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_277),
.B(n_291),
.C(n_292),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

MAJx2_ASAP7_75t_L g406 ( 
.A(n_278),
.B(n_285),
.C(n_288),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_285),
.B1(n_288),
.B2(n_289),
.Y(n_280)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_281),
.Y(n_288)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx8_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_285),
.Y(n_289)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_298),
.C(n_312),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_295),
.B(n_387),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_298),
.B(n_312),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.C(n_305),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_299),
.B(n_300),
.Y(n_375)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_305),
.B(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_310),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_306),
.B(n_310),
.Y(n_355)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

OAI21x1_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_384),
.B(n_388),
.Y(n_314)
);

OA21x2_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_369),
.B(n_383),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_352),
.B(n_368),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_318),
.A2(n_342),
.B(n_351),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_325),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_319),
.B(n_325),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_322),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_320),
.B(n_322),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_320),
.B(n_347),
.Y(n_346)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_327),
.B1(n_334),
.B2(n_335),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_330),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_328),
.B(n_330),
.C(n_334),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_340),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_336),
.B(n_340),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_343),
.A2(n_346),
.B(n_350),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_344),
.B(n_345),
.Y(n_350)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_353),
.B(n_367),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_353),
.B(n_367),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_357),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_355),
.B(n_356),
.C(n_371),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_357),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_358),
.B(n_362),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_358),
.B(n_364),
.C(n_366),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

INVx11_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_363),
.A2(n_364),
.B1(n_365),
.B2(n_366),
.Y(n_362)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_363),
.Y(n_366)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_372),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_370),
.B(n_372),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_373),
.A2(n_374),
.B1(n_376),
.B2(n_377),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_373),
.B(n_379),
.C(n_380),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_379),
.B1(n_380),
.B2(n_381),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_381),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_386),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_385),
.B(n_386),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_391),
.B(n_426),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_391),
.B(n_426),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_408),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_394),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_393),
.B(n_394),
.C(n_408),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_395),
.A2(n_396),
.B1(n_405),
.B2(n_407),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_397),
.B(n_398),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_397),
.B(n_400),
.C(n_402),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_399),
.A2(n_400),
.B1(n_402),
.B2(n_403),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_405),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_409),
.B(n_411),
.C(n_421),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_421),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_416),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_412),
.B(n_417),
.C(n_418),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_425),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_423),
.B(n_424),
.C(n_425),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_429),
.B(n_430),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_432),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_431),
.B(n_448),
.C(n_456),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_433),
.A2(n_448),
.B1(n_456),
.B2(n_457),
.Y(n_432)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_433),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_434),
.A2(n_435),
.B1(n_436),
.B2(n_447),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_434),
.B(n_437),
.C(n_438),
.Y(n_461)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_436),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_437),
.B(n_438),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_446),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_441),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_440),
.B(n_441),
.C(n_446),
.Y(n_470)
);

INVx6_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx5_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_448),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_450),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_449),
.B(n_451),
.C(n_452),
.Y(n_468)
);

BUFx24_ASAP7_75t_SL g500 ( 
.A(n_449),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_452),
.Y(n_450)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_460),
.B(n_474),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_460),
.B(n_474),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_462),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_461),
.B(n_463),
.C(n_466),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_466),
.Y(n_462)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_464),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_467),
.A2(n_468),
.B1(n_469),
.B2(n_473),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_467),
.B(n_470),
.C(n_471),
.Y(n_478)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_469),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_SL g469 ( 
.A(n_470),
.B(n_471),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_477),
.B(n_484),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_477),
.B(n_484),
.Y(n_485)
);

BUFx24_ASAP7_75t_SL g499 ( 
.A(n_477),
.Y(n_499)
);

FAx1_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_479),
.CI(n_482),
.CON(n_477),
.SN(n_477)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_478),
.B(n_479),
.C(n_482),
.Y(n_488)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_488),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_487),
.B(n_488),
.Y(n_490)
);

BUFx24_ASAP7_75t_SL g497 ( 
.A(n_487),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx13_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx6_ASAP7_75t_L g495 ( 
.A(n_493),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_496),
.Y(n_494)
);


endmodule