module fake_jpeg_1151_n_607 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_607);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_607;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_419;
wire n_132;
wire n_133;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_19),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_57),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_58),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_20),
.B(n_9),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_60),
.B(n_68),
.Y(n_125)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_62),
.Y(n_146)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_64),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_65),
.Y(n_155)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_20),
.B(n_9),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_69),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_70),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_71),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_72),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_37),
.A2(n_9),
.B1(n_1),
.B2(n_2),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_73),
.A2(n_48),
.B1(n_24),
.B2(n_52),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_74),
.Y(n_161)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_76),
.Y(n_171)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_78),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_83),
.Y(n_173)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

BUFx24_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_86),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_10),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_87),
.B(n_109),
.Y(n_139)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_21),
.B(n_10),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_90),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_47),
.B(n_8),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_91),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_21),
.B(n_8),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_108),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_94),
.Y(n_165)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_97),
.Y(n_158)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_98),
.Y(n_162)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_37),
.Y(n_100)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_40),
.Y(n_102)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

BUFx10_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_44),
.Y(n_107)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_37),
.B(n_8),
.Y(n_108)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_44),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_46),
.Y(n_110)
);

BUFx12f_ASAP7_75t_SL g113 ( 
.A(n_110),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_23),
.B(n_11),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_26),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_75),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_116),
.B(n_76),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_64),
.A2(n_44),
.B1(n_54),
.B2(n_51),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g187 ( 
.A1(n_121),
.A2(n_170),
.B1(n_86),
.B2(n_69),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_91),
.C(n_108),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_123),
.B(n_42),
.C(n_27),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_56),
.B(n_23),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_127),
.B(n_138),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_59),
.B(n_55),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_55),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_141),
.B(n_152),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_63),
.B(n_26),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_153),
.B(n_43),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_174),
.B1(n_48),
.B2(n_41),
.Y(n_182)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_82),
.Y(n_164)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_66),
.B(n_50),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_83),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_57),
.A2(n_46),
.B1(n_49),
.B2(n_51),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_168),
.A2(n_48),
.B1(n_49),
.B2(n_54),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_72),
.A2(n_54),
.B1(n_49),
.B2(n_51),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_73),
.A2(n_54),
.B1(n_51),
.B2(n_49),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_86),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_175),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_122),
.A2(n_80),
.B1(n_105),
.B2(n_103),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_177),
.A2(n_180),
.B1(n_186),
.B2(n_201),
.Y(n_275)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_179),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_124),
.A2(n_65),
.B1(n_62),
.B2(n_102),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_168),
.A2(n_70),
.B1(n_58),
.B2(n_101),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_181),
.A2(n_182),
.B1(n_209),
.B2(n_221),
.Y(n_272)
);

AO22x1_ASAP7_75t_SL g183 ( 
.A1(n_139),
.A2(n_110),
.B1(n_92),
.B2(n_71),
.Y(n_183)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_183),
.Y(n_246)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_132),
.Y(n_184)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_184),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_187),
.B(n_211),
.Y(n_285)
);

BUFx12f_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_189),
.Y(n_269)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_114),
.Y(n_190)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_190),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_191),
.Y(n_241)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_128),
.Y(n_193)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_193),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_194),
.B(n_212),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_137),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_195),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_149),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_196),
.B(n_204),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_153),
.B(n_29),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_197),
.B(n_200),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_149),
.A2(n_104),
.B1(n_110),
.B2(n_52),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_198),
.Y(n_248)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_118),
.Y(n_199)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_199),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_125),
.B(n_50),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_139),
.A2(n_170),
.B1(n_121),
.B2(n_130),
.Y(n_201)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_137),
.Y(n_202)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_202),
.Y(n_271)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_147),
.Y(n_203)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_203),
.Y(n_293)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_205),
.Y(n_267)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_206),
.Y(n_270)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_115),
.Y(n_207)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_207),
.Y(n_251)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_151),
.Y(n_208)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_208),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_119),
.A2(n_94),
.B1(n_74),
.B2(n_29),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_134),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_210),
.Y(n_265)
);

OA22x2_ASAP7_75t_L g211 ( 
.A1(n_129),
.A2(n_24),
.B1(n_27),
.B2(n_32),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_145),
.B(n_43),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_156),
.Y(n_213)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_213),
.Y(n_279)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_140),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_214),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_126),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_215),
.Y(n_292)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_140),
.Y(n_216)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_216),
.Y(n_280)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_136),
.Y(n_217)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_217),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_158),
.B(n_33),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_220),
.Y(n_249)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_157),
.Y(n_219)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_219),
.Y(n_294)
);

INVx3_ASAP7_75t_SL g220 ( 
.A(n_126),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_113),
.A2(n_24),
.B1(n_52),
.B2(n_45),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_157),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_223),
.Y(n_254)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_150),
.Y(n_223)
);

AND2x2_ASAP7_75t_SL g224 ( 
.A(n_173),
.B(n_45),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_0),
.Y(n_250)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_166),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_227),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_154),
.A2(n_33),
.B1(n_53),
.B2(n_30),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_226),
.A2(n_235),
.B1(n_237),
.B2(n_238),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_133),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_146),
.Y(n_228)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

AOI32xp33_ASAP7_75t_L g229 ( 
.A1(n_144),
.A2(n_30),
.A3(n_53),
.B1(n_45),
.B2(n_32),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_230),
.Y(n_258)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_112),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_232),
.Y(n_259)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_120),
.Y(n_232)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_135),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_233),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_146),
.Y(n_234)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_L g235 ( 
.A1(n_154),
.A2(n_42),
.B1(n_27),
.B2(n_32),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_133),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_236),
.B(n_239),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_161),
.A2(n_41),
.B1(n_42),
.B2(n_88),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_L g238 ( 
.A1(n_161),
.A2(n_41),
.B1(n_99),
.B2(n_78),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_117),
.B(n_67),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_144),
.A2(n_109),
.B1(n_25),
.B2(n_2),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_240),
.A2(n_135),
.B1(n_148),
.B2(n_165),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_181),
.A2(n_171),
.B1(n_155),
.B2(n_176),
.Y(n_242)
);

AO22x1_ASAP7_75t_L g326 ( 
.A1(n_242),
.A2(n_234),
.B1(n_228),
.B2(n_131),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_238),
.A2(n_176),
.B1(n_155),
.B2(n_163),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_245),
.A2(n_286),
.B1(n_165),
.B2(n_131),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_250),
.B(n_211),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_224),
.B(n_171),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_260),
.B(n_261),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_224),
.B(n_163),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_188),
.A2(n_148),
.B(n_160),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_264),
.A2(n_25),
.B(n_143),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_215),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_287),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_192),
.B(n_172),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_277),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_230),
.B(n_142),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_278),
.B(n_290),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_282),
.A2(n_248),
.B1(n_286),
.B2(n_242),
.Y(n_341)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_195),
.Y(n_284)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_284),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_183),
.A2(n_160),
.B1(n_120),
.B2(n_131),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_233),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_183),
.B(n_165),
.Y(n_290)
);

AND2x6_ASAP7_75t_L g291 ( 
.A(n_204),
.B(n_143),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_264),
.Y(n_297)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_263),
.Y(n_296)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_296),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_297),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_246),
.A2(n_187),
.B1(n_221),
.B2(n_198),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_298),
.A2(n_311),
.B1(n_326),
.B2(n_248),
.Y(n_351)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_263),
.Y(n_299)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_299),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_300),
.B(n_303),
.Y(n_364)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_255),
.Y(n_301)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_301),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_278),
.B(n_185),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_246),
.A2(n_211),
.B1(n_235),
.B2(n_219),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_304),
.A2(n_341),
.B1(n_273),
.B2(n_269),
.Y(n_370)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_280),
.Y(n_305)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_305),
.Y(n_360)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_280),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_306),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_241),
.B(n_178),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_307),
.B(n_313),
.Y(n_377)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_279),
.Y(n_308)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_308),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_243),
.B(n_178),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_310),
.B(n_316),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_275),
.A2(n_187),
.B1(n_240),
.B2(n_202),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_249),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_312),
.B(n_327),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_276),
.B(n_203),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_244),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_314),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_276),
.B(n_222),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_315),
.B(n_320),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_258),
.B(n_231),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_279),
.Y(n_317)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_317),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_285),
.A2(n_207),
.B1(n_208),
.B2(n_220),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_319),
.A2(n_325),
.B(n_342),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_274),
.B(n_268),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_268),
.Y(n_321)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_321),
.Y(n_355)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_244),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_322),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_260),
.B(n_179),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_323),
.B(n_333),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_261),
.B(n_189),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_324),
.B(n_334),
.Y(n_361)
);

NAND2xp33_ASAP7_75t_SL g325 ( 
.A(n_285),
.B(n_189),
.Y(n_325)
);

NAND3xp33_ASAP7_75t_L g327 ( 
.A(n_262),
.B(n_216),
.C(n_214),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_253),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_328),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_SL g380 ( 
.A1(n_329),
.A2(n_343),
.B1(n_324),
.B2(n_300),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_250),
.B(n_205),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_330),
.B(n_294),
.C(n_287),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_270),
.B(n_205),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_331),
.A2(n_307),
.B(n_295),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_254),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_332),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_290),
.B(n_0),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_285),
.B(n_0),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_259),
.B(n_0),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_335),
.B(n_336),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_247),
.B(n_1),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_270),
.Y(n_337)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_337),
.Y(n_372)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_288),
.Y(n_339)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_339),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_294),
.B(n_3),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_340),
.B(n_265),
.Y(n_387)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_288),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_318),
.A2(n_333),
.B1(n_303),
.B2(n_275),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_345),
.A2(n_369),
.B1(n_326),
.B2(n_336),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_351),
.A2(n_370),
.B1(n_374),
.B2(n_379),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_352),
.B(n_339),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_318),
.B(n_291),
.C(n_252),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_357),
.B(n_324),
.C(n_334),
.Y(n_389)
);

O2A1O1Ixp33_ASAP7_75t_SL g362 ( 
.A1(n_298),
.A2(n_283),
.B(n_272),
.C(n_282),
.Y(n_362)
);

OA21x2_ASAP7_75t_L g407 ( 
.A1(n_362),
.A2(n_351),
.B(n_368),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_295),
.Y(n_366)
);

CKINVDCx14_ASAP7_75t_R g391 ( 
.A(n_366),
.Y(n_391)
);

FAx1_ASAP7_75t_SL g368 ( 
.A(n_316),
.B(n_247),
.CI(n_283),
.CON(n_368),
.SN(n_368)
);

FAx1_ASAP7_75t_SL g394 ( 
.A(n_368),
.B(n_376),
.CI(n_342),
.CON(n_394),
.SN(n_394)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_302),
.A2(n_271),
.B1(n_284),
.B2(n_253),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_325),
.A2(n_269),
.B(n_251),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_371),
.A2(n_385),
.B(n_337),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_373),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_309),
.A2(n_271),
.B1(n_281),
.B2(n_251),
.Y(n_374)
);

MAJx2_ASAP7_75t_L g376 ( 
.A(n_330),
.B(n_252),
.C(n_257),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_311),
.A2(n_266),
.B1(n_281),
.B2(n_289),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_380),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_300),
.A2(n_266),
.B1(n_289),
.B2(n_293),
.Y(n_381)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_381),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_331),
.Y(n_383)
);

NAND3xp33_ASAP7_75t_L g419 ( 
.A(n_383),
.B(n_256),
.C(n_338),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_320),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_384),
.B(n_5),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_334),
.A2(n_257),
.B(n_267),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_387),
.B(n_343),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_364),
.B(n_301),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_388),
.B(n_390),
.C(n_396),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_389),
.B(n_401),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_352),
.B(n_302),
.C(n_315),
.Y(n_390)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_346),
.Y(n_392)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_392),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_394),
.B(n_424),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_376),
.B(n_313),
.C(n_323),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_384),
.B(n_335),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_398),
.B(n_420),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_399),
.A2(n_407),
.B1(n_415),
.B2(n_418),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_359),
.A2(n_319),
.B(n_340),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_400),
.A2(n_406),
.B(n_417),
.Y(n_452)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_346),
.Y(n_403)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_403),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_357),
.B(n_296),
.C(n_299),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_404),
.B(n_405),
.C(n_413),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_364),
.B(n_321),
.C(n_317),
.Y(n_405)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_347),
.Y(n_408)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_408),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_350),
.B(n_308),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_409),
.B(n_416),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_362),
.A2(n_379),
.B1(n_366),
.B2(n_368),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_410),
.A2(n_412),
.B1(n_361),
.B2(n_377),
.Y(n_433)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_347),
.Y(n_411)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_411),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_362),
.A2(n_329),
.B1(n_326),
.B2(n_306),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_349),
.B(n_305),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_414),
.B(n_361),
.C(n_387),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_345),
.A2(n_328),
.B1(n_322),
.B2(n_314),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_350),
.B(n_265),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_359),
.A2(n_267),
.B(n_293),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_369),
.A2(n_338),
.B1(n_256),
.B2(n_292),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_419),
.A2(n_400),
.B1(n_393),
.B2(n_395),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_373),
.Y(n_420)
);

OAI21x1_ASAP7_75t_R g421 ( 
.A1(n_377),
.A2(n_143),
.B(n_292),
.Y(n_421)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_421),
.Y(n_439)
);

BUFx24_ASAP7_75t_SL g422 ( 
.A(n_344),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_422),
.B(n_423),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_365),
.B(n_4),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_353),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_353),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_425),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_426),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_417),
.B(n_385),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_431),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_432),
.B(n_25),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_433),
.A2(n_449),
.B1(n_394),
.B2(n_424),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_391),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_434),
.B(n_443),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_404),
.B(n_349),
.C(n_361),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_435),
.B(n_442),
.Y(n_468)
);

AOI22x1_ASAP7_75t_L g438 ( 
.A1(n_410),
.A2(n_382),
.B1(n_344),
.B2(n_372),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_438),
.B(n_378),
.Y(n_480)
);

OA21x2_ASAP7_75t_L g440 ( 
.A1(n_407),
.A2(n_371),
.B(n_382),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_440),
.A2(n_453),
.B(n_457),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_413),
.B(n_356),
.C(n_365),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_426),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_414),
.B(n_375),
.C(n_354),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_444),
.B(n_450),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_421),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_448),
.B(n_454),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_407),
.A2(n_358),
.B1(n_354),
.B2(n_372),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_389),
.B(n_375),
.C(n_355),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_395),
.A2(n_386),
.B(n_355),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_421),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_456),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_406),
.A2(n_386),
.B(n_348),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_399),
.A2(n_393),
.B1(n_397),
.B2(n_415),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_459),
.A2(n_461),
.B1(n_396),
.B2(n_392),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_394),
.A2(n_348),
.B1(n_360),
.B2(n_363),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_418),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_462),
.B(n_12),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_464),
.A2(n_470),
.B1(n_485),
.B2(n_486),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_441),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_465),
.B(n_467),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_452),
.A2(n_402),
.B(n_388),
.Y(n_467)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_427),
.Y(n_469)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_469),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_433),
.A2(n_412),
.B1(n_408),
.B2(n_403),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_453),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_471),
.B(n_479),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_452),
.A2(n_405),
.B(n_390),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_472),
.A2(n_474),
.B1(n_478),
.B2(n_490),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_455),
.Y(n_473)
);

CKINVDCx14_ASAP7_75t_R g510 ( 
.A(n_473),
.Y(n_510)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_427),
.Y(n_475)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_475),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_438),
.Y(n_476)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_476),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_459),
.A2(n_360),
.B1(n_367),
.B2(n_363),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_451),
.Y(n_479)
);

OA21x2_ASAP7_75t_L g506 ( 
.A1(n_480),
.A2(n_494),
.B(n_431),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_460),
.B(n_378),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_482),
.B(n_436),
.Y(n_513)
);

INVx8_ASAP7_75t_L g484 ( 
.A(n_442),
.Y(n_484)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_484),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_449),
.A2(n_367),
.B1(n_6),
.B2(n_7),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_462),
.A2(n_5),
.B1(n_7),
.B2(n_11),
.Y(n_486)
);

MAJx2_ASAP7_75t_L g517 ( 
.A(n_487),
.B(n_489),
.C(n_458),
.Y(n_517)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_488),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_430),
.B(n_12),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_429),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_437),
.B(n_12),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_491),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_437),
.B(n_12),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_492),
.B(n_429),
.Y(n_497)
);

OA21x2_ASAP7_75t_L g494 ( 
.A1(n_447),
.A2(n_14),
.B(n_15),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_473),
.A2(n_447),
.B1(n_431),
.B2(n_457),
.Y(n_495)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_495),
.Y(n_529)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_497),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_SL g499 ( 
.A(n_472),
.B(n_445),
.Y(n_499)
);

XNOR2x2_ASAP7_75t_L g535 ( 
.A(n_499),
.B(n_501),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_SL g501 ( 
.A(n_464),
.B(n_445),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_468),
.B(n_430),
.C(n_450),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_504),
.B(n_515),
.Y(n_523)
);

O2A1O1Ixp33_ASAP7_75t_L g527 ( 
.A1(n_506),
.A2(n_471),
.B(n_477),
.C(n_493),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_468),
.B(n_435),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_507),
.B(n_517),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_470),
.A2(n_461),
.B1(n_440),
.B2(n_448),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_508),
.A2(n_514),
.B1(n_516),
.B2(n_480),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_474),
.B(n_428),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_511),
.B(n_518),
.Y(n_524)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_513),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_465),
.A2(n_438),
.B1(n_440),
.B2(n_454),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_483),
.B(n_428),
.C(n_444),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_466),
.A2(n_439),
.B1(n_436),
.B2(n_432),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_487),
.B(n_446),
.C(n_439),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_467),
.B(n_446),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_520),
.B(n_478),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_519),
.A2(n_493),
.B(n_466),
.Y(n_522)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_522),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_497),
.B(n_481),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_526),
.A2(n_528),
.B1(n_531),
.B2(n_532),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_527),
.B(n_506),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_505),
.A2(n_508),
.B1(n_502),
.B2(n_509),
.Y(n_528)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_502),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_498),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_520),
.A2(n_463),
.B(n_480),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_533),
.A2(n_534),
.B1(n_536),
.B2(n_537),
.Y(n_553)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_503),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_512),
.B(n_492),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_496),
.B(n_491),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_539),
.B(n_540),
.Y(n_545)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_521),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_541),
.B(n_542),
.Y(n_544)
);

OA21x2_ASAP7_75t_L g542 ( 
.A1(n_495),
.A2(n_477),
.B(n_463),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_543),
.A2(n_556),
.B1(n_539),
.B2(n_527),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_538),
.A2(n_510),
.B1(n_505),
.B2(n_479),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_547),
.B(n_548),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_531),
.A2(n_516),
.B1(n_488),
.B2(n_484),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_524),
.B(n_500),
.Y(n_549)
);

NOR2xp67_ASAP7_75t_SL g565 ( 
.A(n_549),
.B(n_550),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_523),
.B(n_507),
.C(n_504),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_530),
.B(n_499),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_551),
.B(n_557),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_529),
.A2(n_490),
.B1(n_475),
.B2(n_469),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_554),
.B(n_555),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_524),
.B(n_515),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_529),
.A2(n_506),
.B1(n_458),
.B2(n_494),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g557 ( 
.A(n_530),
.B(n_511),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_541),
.B(n_518),
.C(n_501),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_558),
.B(n_559),
.C(n_560),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_533),
.B(n_517),
.C(n_489),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_522),
.B(n_494),
.C(n_485),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_528),
.B(n_486),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_SL g564 ( 
.A(n_561),
.B(n_544),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_SL g563 ( 
.A1(n_552),
.A2(n_542),
.B(n_526),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_563),
.B(n_564),
.Y(n_583)
);

CKINVDCx14_ASAP7_75t_R g566 ( 
.A(n_546),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_566),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_550),
.B(n_542),
.C(n_525),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_567),
.B(n_569),
.Y(n_585)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_568),
.B(n_573),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_549),
.B(n_535),
.C(n_537),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_557),
.B(n_535),
.C(n_534),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_570),
.B(n_574),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_553),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_SL g578 ( 
.A(n_571),
.B(n_545),
.Y(n_578)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_543),
.A2(n_532),
.B(n_15),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_561),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_560),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_575),
.B(n_574),
.Y(n_581)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_578),
.Y(n_591)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_581),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_567),
.B(n_544),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_SL g595 ( 
.A(n_584),
.B(n_586),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_SL g586 ( 
.A(n_577),
.B(n_558),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_SL g587 ( 
.A1(n_569),
.A2(n_559),
.B1(n_551),
.B2(n_18),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_SL g593 ( 
.A1(n_587),
.A2(n_575),
.B(n_573),
.Y(n_593)
);

BUFx24_ASAP7_75t_SL g588 ( 
.A(n_576),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_588),
.B(n_562),
.Y(n_589)
);

NOR2x1_ASAP7_75t_L g596 ( 
.A(n_589),
.B(n_580),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_585),
.B(n_562),
.Y(n_590)
);

NOR2xp67_ASAP7_75t_L g598 ( 
.A(n_590),
.B(n_592),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_582),
.B(n_565),
.Y(n_592)
);

INVxp67_ASAP7_75t_L g599 ( 
.A(n_593),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_596),
.B(n_594),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_SL g597 ( 
.A1(n_591),
.A2(n_583),
.B(n_570),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_SL g601 ( 
.A1(n_597),
.A2(n_594),
.B(n_587),
.Y(n_601)
);

OAI21xp5_ASAP7_75t_L g602 ( 
.A1(n_600),
.A2(n_601),
.B(n_598),
.Y(n_602)
);

AOI322xp5_ASAP7_75t_L g603 ( 
.A1(n_602),
.A2(n_599),
.A3(n_593),
.B1(n_595),
.B2(n_579),
.C1(n_568),
.C2(n_564),
.Y(n_603)
);

OAI211xp5_ASAP7_75t_L g604 ( 
.A1(n_603),
.A2(n_579),
.B(n_572),
.C(n_18),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_604),
.B(n_572),
.C(n_17),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_L g606 ( 
.A1(n_605),
.A2(n_16),
.B(n_19),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_L g607 ( 
.A1(n_606),
.A2(n_19),
.B(n_434),
.Y(n_607)
);


endmodule