module fake_jpeg_8605_n_78 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx3_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_5),
.B(n_0),
.Y(n_12)
);

BUFx12_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_18),
.Y(n_25)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_21),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_21),
.A2(n_12),
.B1(n_11),
.B2(n_14),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_23),
.A2(n_11),
.B1(n_15),
.B2(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_12),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_25),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_31),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_35),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_36),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_26),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_10),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_42),
.B(n_43),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_15),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_40),
.B1(n_36),
.B2(n_35),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_27),
.B1(n_33),
.B2(n_9),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_32),
.C(n_31),
.Y(n_48)
);

NOR3xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_49),
.C(n_27),
.Y(n_55)
);

AO21x1_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_20),
.B(n_17),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_24),
.C(n_17),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_9),
.C(n_24),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_7),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_55),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_46),
.C(n_13),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_49),
.A2(n_13),
.B(n_1),
.Y(n_56)
);

XNOR2x1_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_13),
.Y(n_63)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_4),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_57),
.B(n_48),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_61),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_53),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_55),
.C(n_13),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_64),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_60),
.C(n_1),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_59),
.Y(n_68)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_70),
.C(n_0),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_65),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_71),
.B(n_66),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_73),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_69),
.C(n_1),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_74),
.B(n_0),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_2),
.Y(n_78)
);


endmodule