module real_aes_6868_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_374;
wire n_379;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
A2O1A1Ixp33_ASAP7_75t_SL g236 ( .A1(n_0), .A2(n_237), .B(n_240), .C(n_244), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_1), .B(n_228), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_2), .A2(n_80), .B1(n_81), .B2(n_161), .Y(n_79) );
INVx1_ASAP7_75t_L g161 ( .A(n_2), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_3), .B(n_238), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_4), .A2(n_197), .B(n_293), .Y(n_292) );
AO21x2_ASAP7_75t_L g301 ( .A1(n_5), .A2(n_230), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g183 ( .A(n_6), .Y(n_183) );
AND2x6_ASAP7_75t_L g202 ( .A(n_6), .B(n_181), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_6), .B(n_517), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g318 ( .A1(n_7), .A2(n_202), .B(n_204), .C(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g84 ( .A(n_8), .B(n_85), .Y(n_84) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_9), .A2(n_21), .B1(n_89), .B2(n_94), .Y(n_93) );
INVx1_ASAP7_75t_L g222 ( .A(n_10), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g141 ( .A1(n_11), .A2(n_76), .B1(n_142), .B2(n_145), .Y(n_141) );
AOI22xp5_ASAP7_75t_L g163 ( .A1(n_12), .A2(n_164), .B1(n_165), .B2(n_166), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_12), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g308 ( .A(n_12), .B(n_238), .Y(n_308) );
AO22x2_ASAP7_75t_L g88 ( .A1(n_13), .A2(n_23), .B1(n_89), .B2(n_90), .Y(n_88) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_14), .A2(n_204), .B(n_207), .C(n_215), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g304 ( .A1(n_15), .A2(n_204), .B(n_215), .C(n_305), .Y(n_304) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_16), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g156 ( .A1(n_17), .A2(n_18), .B1(n_157), .B2(n_159), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_19), .A2(n_197), .B(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g200 ( .A(n_20), .Y(n_200) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_22), .A2(n_254), .B(n_255), .C(n_259), .Y(n_253) );
OAI221xp5_ASAP7_75t_L g174 ( .A1(n_23), .A2(n_39), .B1(n_51), .B2(n_175), .C(n_176), .Y(n_174) );
INVxp67_ASAP7_75t_L g177 ( .A(n_23), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_24), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_25), .B(n_196), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g323 ( .A(n_26), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_27), .A2(n_58), .B1(n_106), .B2(n_112), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g99 ( .A(n_28), .B(n_100), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_29), .B(n_238), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_29), .A2(n_80), .B1(n_81), .B2(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_29), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g133 ( .A1(n_30), .A2(n_46), .B1(n_134), .B2(n_137), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_31), .B(n_197), .Y(n_303) );
INVx1_ASAP7_75t_L g122 ( .A(n_32), .Y(n_122) );
A2O1A1Ixp33_ASAP7_75t_L g283 ( .A1(n_33), .A2(n_254), .B(n_259), .C(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g241 ( .A(n_34), .Y(n_241) );
INVx1_ASAP7_75t_L g285 ( .A(n_35), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g162 ( .A1(n_36), .A2(n_163), .B1(n_169), .B2(n_170), .Y(n_162) );
INVx1_ASAP7_75t_L g169 ( .A(n_36), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_37), .B(n_197), .Y(n_282) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_38), .Y(n_224) );
AO22x2_ASAP7_75t_L g98 ( .A1(n_39), .A2(n_61), .B1(n_89), .B2(n_90), .Y(n_98) );
INVxp67_ASAP7_75t_L g178 ( .A(n_39), .Y(n_178) );
OAI22xp5_ASAP7_75t_SL g166 ( .A1(n_40), .A2(n_63), .B1(n_167), .B2(n_168), .Y(n_166) );
INVx1_ASAP7_75t_L g168 ( .A(n_40), .Y(n_168) );
INVx1_ASAP7_75t_L g181 ( .A(n_41), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_42), .B(n_197), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_43), .B(n_228), .Y(n_298) );
A2O1A1Ixp33_ASAP7_75t_L g295 ( .A1(n_44), .A2(n_214), .B(n_270), .C(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g221 ( .A(n_45), .Y(n_221) );
AOI22xp33_ASAP7_75t_SL g150 ( .A1(n_47), .A2(n_54), .B1(n_151), .B2(n_153), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_48), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_49), .B(n_238), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_50), .B(n_239), .Y(n_320) );
AO22x2_ASAP7_75t_L g96 ( .A1(n_51), .A2(n_67), .B1(n_89), .B2(n_94), .Y(n_96) );
AOI22xp5_ASAP7_75t_L g123 ( .A1(n_52), .A2(n_71), .B1(n_124), .B2(n_127), .Y(n_123) );
CKINVDCx16_ASAP7_75t_R g234 ( .A(n_53), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_55), .B(n_209), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_56), .A2(n_204), .B(n_259), .C(n_268), .Y(n_267) );
CKINVDCx16_ASAP7_75t_R g294 ( .A(n_57), .Y(n_294) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_59), .B(n_212), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g261 ( .A(n_60), .Y(n_261) );
INVx2_ASAP7_75t_L g219 ( .A(n_62), .Y(n_219) );
INVx1_ASAP7_75t_L g167 ( .A(n_63), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g277 ( .A(n_64), .Y(n_277) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_65), .B(n_243), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_66), .B(n_197), .Y(n_252) );
INVx1_ASAP7_75t_L g256 ( .A(n_68), .Y(n_256) );
INVxp67_ASAP7_75t_L g297 ( .A(n_69), .Y(n_297) );
INVx1_ASAP7_75t_L g89 ( .A(n_70), .Y(n_89) );
INVx1_ASAP7_75t_L g91 ( .A(n_70), .Y(n_91) );
INVx1_ASAP7_75t_L g269 ( .A(n_72), .Y(n_269) );
INVx1_ASAP7_75t_L g316 ( .A(n_73), .Y(n_316) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_74), .A2(n_80), .B1(n_81), .B2(n_525), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_74), .Y(n_525) );
AND2x2_ASAP7_75t_L g287 ( .A(n_75), .B(n_218), .Y(n_287) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_171), .B1(n_184), .B2(n_506), .C(n_511), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_162), .Y(n_78) );
INVx1_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
NAND2x1p5_ASAP7_75t_L g81 ( .A(n_82), .B(n_131), .Y(n_81) );
NOR2xp33_ASAP7_75t_L g82 ( .A(n_83), .B(n_116), .Y(n_82) );
NAND3xp33_ASAP7_75t_L g83 ( .A(n_84), .B(n_99), .C(n_105), .Y(n_83) );
BUFx2_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
AND2x6_ASAP7_75t_L g86 ( .A(n_87), .B(n_95), .Y(n_86) );
AND2x4_ASAP7_75t_L g152 ( .A(n_87), .B(n_120), .Y(n_152) );
AND2x2_ASAP7_75t_L g155 ( .A(n_87), .B(n_139), .Y(n_155) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_92), .Y(n_87) );
OR2x2_ASAP7_75t_L g104 ( .A(n_88), .B(n_92), .Y(n_104) );
INVx2_ASAP7_75t_L g110 ( .A(n_88), .Y(n_110) );
INVx1_ASAP7_75t_L g115 ( .A(n_88), .Y(n_115) );
AND2x2_ASAP7_75t_L g119 ( .A(n_88), .B(n_93), .Y(n_119) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g94 ( .A(n_91), .Y(n_94) );
AND2x2_ASAP7_75t_L g140 ( .A(n_92), .B(n_110), .Y(n_140) );
INVx2_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
AND2x2_ASAP7_75t_L g111 ( .A(n_93), .B(n_98), .Y(n_111) );
AND2x4_ASAP7_75t_L g102 ( .A(n_95), .B(n_103), .Y(n_102) );
AND2x4_ASAP7_75t_L g158 ( .A(n_95), .B(n_140), .Y(n_158) );
AND2x2_ASAP7_75t_L g95 ( .A(n_96), .B(n_97), .Y(n_95) );
INVx1_ASAP7_75t_L g109 ( .A(n_96), .Y(n_109) );
INVx1_ASAP7_75t_L g121 ( .A(n_96), .Y(n_121) );
INVx1_ASAP7_75t_L g130 ( .A(n_96), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_96), .B(n_98), .Y(n_148) );
AND2x2_ASAP7_75t_L g120 ( .A(n_97), .B(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x2_ASAP7_75t_L g139 ( .A(n_98), .B(n_130), .Y(n_139) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx4_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x6_ASAP7_75t_L g136 ( .A(n_103), .B(n_120), .Y(n_136) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x4_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g126 ( .A(n_109), .Y(n_126) );
AND2x4_ASAP7_75t_L g113 ( .A(n_111), .B(n_114), .Y(n_113) );
AND2x4_ASAP7_75t_L g125 ( .A(n_111), .B(n_126), .Y(n_125) );
BUFx3_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OR2x6_ASAP7_75t_L g160 ( .A(n_115), .B(n_148), .Y(n_160) );
OAI21xp5_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_122), .B(n_123), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x6_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
AND2x4_ASAP7_75t_L g128 ( .A(n_119), .B(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g144 ( .A(n_120), .B(n_140), .Y(n_144) );
BUFx12f_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NOR2x1_ASAP7_75t_L g131 ( .A(n_132), .B(n_149), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_141), .Y(n_132) );
INVx2_ASAP7_75t_SL g134 ( .A(n_135), .Y(n_134) );
INVx11_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x4_ASAP7_75t_L g146 ( .A(n_140), .B(n_147), .Y(n_146) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_150), .B(n_156), .Y(n_149) );
BUFx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx5_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx8_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_SL g159 ( .A(n_160), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_163), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_166), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g171 ( .A(n_172), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_173), .Y(n_172) );
AND3x1_ASAP7_75t_SL g173 ( .A(n_174), .B(n_179), .C(n_182), .Y(n_173) );
INVxp67_ASAP7_75t_L g517 ( .A(n_174), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
INVx1_ASAP7_75t_SL g518 ( .A(n_179), .Y(n_518) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_179), .A2(n_521), .B(n_523), .Y(n_520) );
INVx1_ASAP7_75t_L g527 ( .A(n_179), .Y(n_527) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_180), .B(n_183), .Y(n_523) );
HB1xp67_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
OR2x2_ASAP7_75t_SL g526 ( .A(n_182), .B(n_527), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_SL g185 ( .A(n_186), .B(n_461), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_187), .B(n_396), .Y(n_186) );
NAND4xp25_ASAP7_75t_SL g187 ( .A(n_188), .B(n_341), .C(n_365), .D(n_388), .Y(n_187) );
AOI221xp5_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_278), .B1(n_312), .B2(n_325), .C(n_328), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_191), .B(n_248), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_191), .A2(n_226), .B1(n_279), .B2(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_191), .B(n_249), .Y(n_399) );
AND2x2_ASAP7_75t_L g418 ( .A(n_191), .B(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_191), .B(n_402), .Y(n_488) );
AND2x4_ASAP7_75t_L g191 ( .A(n_192), .B(n_226), .Y(n_191) );
AND2x2_ASAP7_75t_L g356 ( .A(n_192), .B(n_249), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_192), .B(n_371), .Y(n_370) );
OR2x2_ASAP7_75t_L g379 ( .A(n_192), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g384 ( .A(n_192), .B(n_227), .Y(n_384) );
INVx2_ASAP7_75t_L g416 ( .A(n_192), .Y(n_416) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_192), .Y(n_460) );
AND2x2_ASAP7_75t_L g477 ( .A(n_192), .B(n_354), .Y(n_477) );
INVx5_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
AND2x2_ASAP7_75t_L g395 ( .A(n_193), .B(n_354), .Y(n_395) );
AND2x4_ASAP7_75t_L g409 ( .A(n_193), .B(n_226), .Y(n_409) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_193), .Y(n_413) );
AND2x2_ASAP7_75t_L g433 ( .A(n_193), .B(n_348), .Y(n_433) );
AND2x2_ASAP7_75t_L g483 ( .A(n_193), .B(n_250), .Y(n_483) );
AND2x2_ASAP7_75t_L g493 ( .A(n_193), .B(n_227), .Y(n_493) );
OR2x6_ASAP7_75t_L g193 ( .A(n_194), .B(n_223), .Y(n_193) );
AOI21xp5_ASAP7_75t_SL g194 ( .A1(n_195), .A2(n_203), .B(n_216), .Y(n_194) );
BUFx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x4_ASAP7_75t_L g197 ( .A(n_198), .B(n_202), .Y(n_197) );
NAND2x1p5_ASAP7_75t_L g317 ( .A(n_198), .B(n_202), .Y(n_317) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_201), .Y(n_198) );
INVx1_ASAP7_75t_L g214 ( .A(n_199), .Y(n_214) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g205 ( .A(n_200), .Y(n_205) );
INVx1_ASAP7_75t_L g311 ( .A(n_200), .Y(n_311) );
INVx1_ASAP7_75t_L g206 ( .A(n_201), .Y(n_206) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_201), .Y(n_210) );
INVx3_ASAP7_75t_L g239 ( .A(n_201), .Y(n_239) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_201), .Y(n_243) );
INVx1_ASAP7_75t_L g307 ( .A(n_201), .Y(n_307) );
BUFx3_ASAP7_75t_L g215 ( .A(n_202), .Y(n_215) );
INVx4_ASAP7_75t_SL g246 ( .A(n_202), .Y(n_246) );
INVx5_ASAP7_75t_L g235 ( .A(n_204), .Y(n_235) );
AND2x6_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
BUFx3_ASAP7_75t_L g245 ( .A(n_205), .Y(n_245) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_205), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_211), .B(n_213), .Y(n_207) );
INVx2_ASAP7_75t_L g212 ( .A(n_209), .Y(n_212) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx4_ASAP7_75t_L g271 ( .A(n_210), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_L g255 ( .A1(n_212), .A2(n_256), .B(n_257), .C(n_258), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_L g284 ( .A1(n_212), .A2(n_258), .B(n_285), .C(n_286), .Y(n_284) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_212), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_213), .B(n_246), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_213), .B(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g225 ( .A(n_218), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_218), .A2(n_252), .B(n_253), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_218), .A2(n_282), .B(n_283), .Y(n_281) );
AND2x2_ASAP7_75t_SL g218 ( .A(n_219), .B(n_220), .Y(n_218) );
AND2x2_ASAP7_75t_L g231 ( .A(n_219), .B(n_220), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
AND2x2_ASAP7_75t_L g349 ( .A(n_226), .B(n_249), .Y(n_349) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_226), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_226), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g439 ( .A(n_226), .Y(n_439) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g327 ( .A(n_227), .B(n_264), .Y(n_327) );
AND2x2_ASAP7_75t_L g354 ( .A(n_227), .B(n_265), .Y(n_354) );
OA21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_232), .B(n_247), .Y(n_227) );
INVx3_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_229), .B(n_261), .Y(n_260) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_229), .A2(n_266), .B(n_276), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_229), .B(n_277), .Y(n_276) );
AO21x2_ASAP7_75t_L g314 ( .A1(n_229), .A2(n_315), .B(n_322), .Y(n_314) );
INVx4_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_230), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_230), .A2(n_303), .B(n_304), .Y(n_302) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g324 ( .A(n_231), .Y(n_324) );
O2A1O1Ixp33_ASAP7_75t_SL g233 ( .A1(n_234), .A2(n_235), .B(n_236), .C(n_246), .Y(n_233) );
INVx2_ASAP7_75t_L g254 ( .A(n_235), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_L g293 ( .A1(n_235), .A2(n_246), .B(n_294), .C(n_295), .Y(n_293) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_238), .B(n_297), .Y(n_296) );
INVx5_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
INVx4_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_245), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_246), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_248), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_262), .Y(n_248) );
OR2x2_ASAP7_75t_L g380 ( .A(n_249), .B(n_263), .Y(n_380) );
AND2x2_ASAP7_75t_L g417 ( .A(n_249), .B(n_327), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_249), .B(n_348), .Y(n_428) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_249), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_249), .B(n_384), .Y(n_501) );
INVx5_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
BUFx2_ASAP7_75t_L g326 ( .A(n_250), .Y(n_326) );
AND2x2_ASAP7_75t_L g335 ( .A(n_250), .B(n_263), .Y(n_335) );
AND2x2_ASAP7_75t_L g451 ( .A(n_250), .B(n_346), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_250), .B(n_384), .Y(n_473) );
OR2x6_ASAP7_75t_L g250 ( .A(n_251), .B(n_260), .Y(n_250) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_263), .Y(n_419) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_264), .Y(n_371) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
BUFx2_ASAP7_75t_L g348 ( .A(n_265), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_275), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_270), .B(n_272), .C(n_273), .Y(n_268) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_279), .B(n_288), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_279), .B(n_361), .Y(n_480) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_280), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g332 ( .A(n_280), .B(n_333), .Y(n_332) );
INVx5_ASAP7_75t_SL g340 ( .A(n_280), .Y(n_340) );
OR2x2_ASAP7_75t_L g363 ( .A(n_280), .B(n_333), .Y(n_363) );
OR2x2_ASAP7_75t_L g373 ( .A(n_280), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g436 ( .A(n_280), .B(n_290), .Y(n_436) );
AND2x2_ASAP7_75t_SL g474 ( .A(n_280), .B(n_289), .Y(n_474) );
NOR4xp25_ASAP7_75t_L g495 ( .A(n_280), .B(n_416), .C(n_496), .D(n_497), .Y(n_495) );
AND2x2_ASAP7_75t_L g505 ( .A(n_280), .B(n_337), .Y(n_505) );
OR2x6_ASAP7_75t_L g280 ( .A(n_281), .B(n_287), .Y(n_280) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g330 ( .A(n_289), .B(n_326), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_289), .B(n_332), .Y(n_499) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_299), .Y(n_289) );
OR2x2_ASAP7_75t_L g339 ( .A(n_290), .B(n_340), .Y(n_339) );
INVx3_ASAP7_75t_L g346 ( .A(n_290), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_290), .B(n_314), .Y(n_358) );
INVxp67_ASAP7_75t_L g361 ( .A(n_290), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_290), .B(n_333), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_290), .B(n_300), .Y(n_427) );
AND2x2_ASAP7_75t_L g442 ( .A(n_290), .B(n_337), .Y(n_442) );
OR2x2_ASAP7_75t_L g471 ( .A(n_290), .B(n_300), .Y(n_471) );
OA21x2_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_292), .B(n_298), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_299), .B(n_376), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_299), .B(n_340), .Y(n_479) );
OR2x2_ASAP7_75t_L g500 ( .A(n_299), .B(n_377), .Y(n_500) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g313 ( .A(n_300), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g337 ( .A(n_300), .B(n_333), .Y(n_337) );
NAND2xp5_ASAP7_75t_SL g352 ( .A(n_300), .B(n_314), .Y(n_352) );
AND2x2_ASAP7_75t_L g422 ( .A(n_300), .B(n_346), .Y(n_422) );
AND2x2_ASAP7_75t_L g456 ( .A(n_300), .B(n_340), .Y(n_456) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_301), .B(n_340), .Y(n_359) );
AND2x2_ASAP7_75t_L g387 ( .A(n_301), .B(n_314), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_308), .B(n_309), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g319 ( .A1(n_309), .A2(n_320), .B(n_321), .Y(n_319) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx3_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_312), .B(n_395), .Y(n_394) );
AOI221xp5_ASAP7_75t_L g454 ( .A1(n_313), .A2(n_402), .B1(n_438), .B2(n_455), .C(n_457), .Y(n_454) );
INVx5_ASAP7_75t_SL g333 ( .A(n_314), .Y(n_333) );
OAI21xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_317), .B(n_318), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
OAI33xp33_ASAP7_75t_L g353 ( .A1(n_326), .A2(n_354), .A3(n_355), .B1(n_357), .B2(n_360), .B3(n_364), .Y(n_353) );
OR2x2_ASAP7_75t_L g369 ( .A(n_326), .B(n_370), .Y(n_369) );
AOI322xp5_ASAP7_75t_L g478 ( .A1(n_326), .A2(n_395), .A3(n_402), .B1(n_479), .B2(n_480), .C1(n_481), .C2(n_484), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_326), .B(n_354), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_SL g502 ( .A1(n_326), .A2(n_354), .B(n_503), .C(n_505), .Y(n_502) );
AOI221xp5_ASAP7_75t_L g341 ( .A1(n_327), .A2(n_342), .B1(n_347), .B2(n_350), .C(n_353), .Y(n_341) );
INVx1_ASAP7_75t_L g434 ( .A(n_327), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_327), .B(n_483), .Y(n_482) );
OAI22xp33_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_331), .B1(n_334), .B2(n_336), .Y(n_328) );
INVx1_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g411 ( .A(n_332), .B(n_346), .Y(n_411) );
AND2x2_ASAP7_75t_L g469 ( .A(n_332), .B(n_470), .Y(n_469) );
OR2x2_ASAP7_75t_L g377 ( .A(n_333), .B(n_340), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_333), .B(n_346), .Y(n_405) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_335), .B(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_335), .B(n_413), .Y(n_467) );
OAI321xp33_ASAP7_75t_L g486 ( .A1(n_335), .A2(n_408), .A3(n_487), .B1(n_488), .B2(n_489), .C(n_490), .Y(n_486) );
INVx1_ASAP7_75t_L g453 ( .A(n_336), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_337), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g392 ( .A(n_337), .B(n_340), .Y(n_392) );
AOI321xp33_ASAP7_75t_L g450 ( .A1(n_337), .A2(n_354), .A3(n_451), .B1(n_452), .B2(n_453), .C(n_454), .Y(n_450) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g367 ( .A(n_339), .B(n_352), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_340), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_340), .B(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_340), .B(n_426), .Y(n_463) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g386 ( .A(n_344), .B(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g351 ( .A(n_345), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g459 ( .A(n_346), .Y(n_459) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_349), .B(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g382 ( .A(n_354), .Y(n_382) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_356), .B(n_391), .Y(n_440) );
OR2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
OR2x2_ASAP7_75t_L g404 ( .A(n_359), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g449 ( .A(n_359), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_360), .A2(n_407), .B1(n_410), .B2(n_412), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g504 ( .A(n_363), .B(n_427), .Y(n_504) );
AOI221xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_368), .B1(n_372), .B2(n_378), .C(n_381), .Y(n_365) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx2_ASAP7_75t_L g402 ( .A(n_371), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_375), .Y(n_372) );
INVx1_ASAP7_75t_SL g448 ( .A(n_374), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_376), .B(n_426), .Y(n_425) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_376), .A2(n_444), .B(n_446), .Y(n_443) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g489 ( .A(n_377), .B(n_471), .Y(n_489) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_SL g391 ( .A(n_380), .Y(n_391) );
AOI21xp33_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_383), .B(n_385), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g435 ( .A(n_387), .B(n_436), .Y(n_435) );
INVxp67_ASAP7_75t_L g497 ( .A(n_387), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_392), .B(n_393), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_391), .B(n_409), .Y(n_445) );
INVxp67_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g466 ( .A(n_395), .Y(n_466) );
NAND5xp2_ASAP7_75t_L g396 ( .A(n_397), .B(n_414), .C(n_423), .D(n_443), .E(n_450), .Y(n_396) );
O2A1O1Ixp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_400), .B(n_403), .C(n_406), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g438 ( .A(n_402), .Y(n_438) );
CKINVDCx16_ASAP7_75t_R g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_410), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g452 ( .A(n_412), .Y(n_452) );
OAI21xp5_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_418), .B(n_420), .Y(n_414) );
AOI221xp5_ASAP7_75t_L g468 ( .A1(n_415), .A2(n_469), .B1(n_472), .B2(n_474), .C(n_475), .Y(n_468) );
AND2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
AOI321xp33_ASAP7_75t_L g423 ( .A1(n_416), .A2(n_424), .A3(n_428), .B1(n_429), .B2(n_435), .C(n_437), .Y(n_423) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g494 ( .A(n_428), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g429 ( .A(n_430), .B(n_434), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g446 ( .A(n_431), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
NOR2xp67_ASAP7_75t_SL g458 ( .A(n_432), .B(n_439), .Y(n_458) );
AOI321xp33_ASAP7_75t_SL g490 ( .A1(n_435), .A2(n_491), .A3(n_492), .B1(n_493), .B2(n_494), .C(n_495), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_439), .B(n_440), .C(n_441), .Y(n_437) );
INVx1_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_448), .B(n_456), .Y(n_485) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND3xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .C(n_460), .Y(n_457) );
NOR3xp33_ASAP7_75t_L g461 ( .A(n_462), .B(n_486), .C(n_498), .Y(n_461) );
OAI211xp5_ASAP7_75t_SL g462 ( .A1(n_463), .A2(n_464), .B(n_468), .C(n_478), .Y(n_462) );
INVxp67_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_466), .B(n_467), .Y(n_465) );
OAI221xp5_ASAP7_75t_L g498 ( .A1(n_467), .A2(n_499), .B1(n_500), .B2(n_501), .C(n_502), .Y(n_498) );
INVx1_ASAP7_75t_L g487 ( .A(n_469), .Y(n_487) );
INVx1_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_SL g491 ( .A(n_489), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
CKINVDCx14_ASAP7_75t_R g503 ( .A(n_504), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_507), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_510), .Y(n_508) );
INVx1_ASAP7_75t_L g522 ( .A(n_509), .Y(n_522) );
OAI322xp33_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .A3(n_514), .B1(n_518), .B2(n_519), .C1(n_524), .C2(n_526), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_515), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_516), .Y(n_515) );
CKINVDCx16_ASAP7_75t_R g519 ( .A(n_520), .Y(n_519) );
endmodule