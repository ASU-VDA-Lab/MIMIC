module fake_jpeg_9752_n_301 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_41),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_39),
.C(n_40),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_20),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_23),
.B1(n_26),
.B2(n_16),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_47),
.B1(n_55),
.B2(n_25),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_23),
.B1(n_26),
.B2(n_16),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_16),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_33),
.Y(n_74)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_22),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_52),
.B(n_17),
.Y(n_72)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_54),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_42),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g88 ( 
.A(n_58),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_61),
.B(n_31),
.Y(n_90)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx4f_ASAP7_75t_SL g84 ( 
.A(n_62),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_70),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_26),
.B1(n_33),
.B2(n_20),
.Y(n_66)
);

OAI32xp33_ASAP7_75t_L g102 ( 
.A1(n_66),
.A2(n_78),
.A3(n_83),
.B1(n_68),
.B2(n_77),
.Y(n_102)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_67),
.B(n_68),
.Y(n_103)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_63),
.A2(n_48),
.B1(n_49),
.B2(n_57),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_69),
.A2(n_81),
.B1(n_59),
.B2(n_19),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_54),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_28),
.C(n_18),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_73),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_86),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_33),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_82),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_76),
.Y(n_101)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_63),
.A2(n_33),
.B1(n_20),
.B2(n_32),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_28),
.B1(n_25),
.B2(n_18),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_31),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_43),
.B(n_31),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_29),
.Y(n_89)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

NOR2x1_ASAP7_75t_R g91 ( 
.A(n_82),
.B(n_53),
.Y(n_91)
);

XNOR2x1_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_84),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_57),
.B(n_62),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_92),
.A2(n_91),
.B(n_94),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_10),
.C(n_14),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_94),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_75),
.B(n_74),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_95),
.A2(n_78),
.B(n_66),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_71),
.B(n_29),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_96),
.B(n_109),
.Y(n_142)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_98),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_99),
.A2(n_102),
.B1(n_67),
.B2(n_78),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_81),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_106),
.Y(n_122)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_65),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_79),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_73),
.A2(n_24),
.B(n_56),
.C(n_61),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_112),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_69),
.A2(n_59),
.B1(n_60),
.B2(n_19),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_113),
.A2(n_88),
.B1(n_78),
.B2(n_66),
.Y(n_121)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_117),
.B(n_118),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_125),
.B1(n_126),
.B2(n_108),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_123),
.B(n_2),
.Y(n_170)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_97),
.A2(n_88),
.B1(n_66),
.B2(n_85),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_97),
.A2(n_85),
.B1(n_87),
.B2(n_65),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_98),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_130),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_137),
.C(n_138),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_87),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_129),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_105),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_17),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_131),
.Y(n_173)
);

OAI21xp33_ASAP7_75t_L g153 ( 
.A1(n_132),
.A2(n_107),
.B(n_104),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_115),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_141),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_101),
.A2(n_17),
.B(n_1),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_135),
.B(n_96),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_80),
.C(n_17),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_17),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_0),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_139),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_92),
.Y(n_140)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_113),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_0),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_110),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_93),
.B(n_0),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_3),
.B(n_6),
.Y(n_172)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_158),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_122),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_156),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_151),
.A2(n_123),
.B1(n_136),
.B2(n_128),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_153),
.B(n_170),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_115),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_160),
.C(n_132),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_155),
.A2(n_157),
.B(n_166),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_135),
.A2(n_109),
.B(n_102),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_163),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_100),
.C(n_99),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_106),
.Y(n_161)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_143),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_169),
.Y(n_183)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_100),
.Y(n_164)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_123),
.A2(n_1),
.B(n_2),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_125),
.A2(n_112),
.B1(n_111),
.B2(n_1),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_168),
.A2(n_174),
.B1(n_141),
.B2(n_119),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_139),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_118),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_171),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_172),
.B(n_134),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_121),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_177),
.A2(n_171),
.B1(n_145),
.B2(n_163),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_182),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_137),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_191),
.C(n_196),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_147),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_165),
.A2(n_120),
.B1(n_127),
.B2(n_130),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_184),
.A2(n_200),
.B1(n_202),
.B2(n_174),
.Y(n_205)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_147),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_189),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_161),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_148),
.B(n_120),
.Y(n_190)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_190),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_117),
.Y(n_192)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_158),
.B(n_131),
.Y(n_193)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_193),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_194),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_146),
.B(n_144),
.C(n_8),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_156),
.B(n_164),
.Y(n_197)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_146),
.B(n_144),
.C(n_8),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_199),
.C(n_172),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_155),
.B(n_7),
.C(n_8),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_152),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_189),
.Y(n_210)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_204),
.B(n_199),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_205),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_160),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_213),
.Y(n_226)
);

FAx1_ASAP7_75t_SL g209 ( 
.A(n_195),
.B(n_157),
.CI(n_170),
.CON(n_209),
.SN(n_209)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_186),
.Y(n_231)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_152),
.C(n_150),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_217),
.C(n_220),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_167),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_188),
.A2(n_149),
.B(n_165),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_214),
.A2(n_222),
.B(n_186),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_202),
.A2(n_188),
.B1(n_187),
.B2(n_201),
.Y(n_215)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_173),
.C(n_151),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_218),
.A2(n_206),
.B1(n_207),
.B2(n_217),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_182),
.A2(n_168),
.B1(n_166),
.B2(n_169),
.Y(n_219)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_219),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_175),
.C(n_12),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_176),
.A2(n_11),
.B(n_12),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_11),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_200),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_228),
.B(n_232),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_237),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_234),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_218),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_206),
.A2(n_179),
.B1(n_185),
.B2(n_178),
.Y(n_236)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_236),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_179),
.C(n_185),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_211),
.C(n_213),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_210),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_183),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_241),
.B(n_243),
.Y(n_257)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_242),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_214),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_219),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_238),
.Y(n_254)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_237),
.Y(n_247)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_247),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_236),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_250),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_230),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_239),
.C(n_235),
.Y(n_260)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_233),
.A2(n_216),
.B1(n_223),
.B2(n_224),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_253),
.A2(n_244),
.B1(n_238),
.B2(n_233),
.Y(n_263)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_221),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_258),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_261),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_256),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_263),
.A2(n_245),
.B1(n_209),
.B2(n_234),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_257),
.A2(n_227),
.B1(n_240),
.B2(n_229),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_269),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_249),
.A2(n_229),
.B(n_222),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_268),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_253),
.B(n_177),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_256),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_226),
.Y(n_280)
);

OAI221xp5_ASAP7_75t_L g271 ( 
.A1(n_268),
.A2(n_249),
.B1(n_252),
.B2(n_255),
.C(n_235),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_271),
.A2(n_279),
.B(n_280),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_247),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_273),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_246),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_277),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_245),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_259),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_260),
.C(n_261),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_282),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_263),
.C(n_226),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_278),
.A2(n_270),
.B(n_203),
.Y(n_284)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_284),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_220),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_288),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_274),
.A2(n_203),
.B(n_204),
.Y(n_288)
);

NOR2x1_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_225),
.Y(n_291)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_291),
.Y(n_296)
);

NOR2xp67_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_209),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_292),
.B(n_285),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_294),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_293),
.B(n_13),
.C(n_14),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_297),
.B(n_290),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_295),
.C(n_289),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_299),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_296),
.Y(n_301)
);


endmodule