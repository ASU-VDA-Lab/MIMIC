module fake_netlist_1_8791_n_41 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_41);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_40;
wire n_29;
wire n_39;
BUFx2_ASAP7_75t_L g11 ( .A(n_1), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_3), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_3), .B(n_2), .Y(n_13) );
BUFx6f_ASAP7_75t_L g14 ( .A(n_4), .Y(n_14) );
OA21x2_ASAP7_75t_L g15 ( .A1(n_0), .A2(n_9), .B(n_2), .Y(n_15) );
NAND2xp33_ASAP7_75t_R g16 ( .A(n_1), .B(n_7), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_10), .Y(n_17) );
OR2x2_ASAP7_75t_L g18 ( .A(n_11), .B(n_0), .Y(n_18) );
BUFx6f_ASAP7_75t_L g19 ( .A(n_14), .Y(n_19) );
AO22x1_ASAP7_75t_L g20 ( .A1(n_12), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_14), .Y(n_21) );
BUFx6f_ASAP7_75t_L g22 ( .A(n_14), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
BUFx2_ASAP7_75t_L g24 ( .A(n_18), .Y(n_24) );
OAI21xp5_ASAP7_75t_L g25 ( .A1(n_19), .A2(n_17), .B(n_13), .Y(n_25) );
OAI21xp5_ASAP7_75t_SL g26 ( .A1(n_24), .A2(n_14), .B(n_20), .Y(n_26) );
OAI31xp33_ASAP7_75t_L g27 ( .A1(n_24), .A2(n_12), .A3(n_16), .B(n_5), .Y(n_27) );
BUFx2_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
INVxp67_ASAP7_75t_SL g29 ( .A(n_28), .Y(n_29) );
OR2x6_ASAP7_75t_L g30 ( .A(n_26), .B(n_15), .Y(n_30) );
HB1xp67_ASAP7_75t_L g31 ( .A(n_30), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g32 ( .A(n_29), .B(n_27), .Y(n_32) );
OAI211xp5_ASAP7_75t_SL g33 ( .A1(n_32), .A2(n_23), .B(n_30), .C(n_17), .Y(n_33) );
AOI211xp5_ASAP7_75t_L g34 ( .A1(n_31), .A2(n_14), .B(n_28), .C(n_22), .Y(n_34) );
OR2x2_ASAP7_75t_L g35 ( .A(n_32), .B(n_30), .Y(n_35) );
CKINVDCx5p33_ASAP7_75t_R g36 ( .A(n_35), .Y(n_36) );
OR3x2_ASAP7_75t_L g37 ( .A(n_33), .B(n_15), .C(n_23), .Y(n_37) );
NAND4xp25_ASAP7_75t_L g38 ( .A(n_34), .B(n_15), .C(n_22), .D(n_19), .Y(n_38) );
NAND2xp5_ASAP7_75t_L g39 ( .A(n_36), .B(n_22), .Y(n_39) );
INVx1_ASAP7_75t_L g40 ( .A(n_37), .Y(n_40) );
AOI32xp33_ASAP7_75t_L g41 ( .A1(n_40), .A2(n_8), .A3(n_19), .B1(n_38), .B2(n_39), .Y(n_41) );
endmodule