module fake_aes_12564_n_718 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_718);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_718;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_638;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx3_ASAP7_75t_L g104 ( .A(n_9), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_34), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_95), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_63), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_99), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_82), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_46), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_27), .Y(n_111) );
INVx3_ASAP7_75t_L g112 ( .A(n_19), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_78), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_93), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_76), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_15), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_90), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_18), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_67), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_80), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_60), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_56), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_87), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_53), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_7), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_70), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_24), .B(n_64), .Y(n_127) );
CKINVDCx16_ASAP7_75t_R g128 ( .A(n_51), .Y(n_128) );
CKINVDCx14_ASAP7_75t_R g129 ( .A(n_15), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_1), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_22), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_71), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_38), .Y(n_133) );
INVx1_ASAP7_75t_SL g134 ( .A(n_96), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_89), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_69), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_65), .Y(n_137) );
INVxp67_ASAP7_75t_L g138 ( .A(n_43), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_30), .Y(n_139) );
HB1xp67_ASAP7_75t_L g140 ( .A(n_62), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_3), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_14), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_48), .B(n_88), .Y(n_143) );
INVx2_ASAP7_75t_SL g144 ( .A(n_98), .Y(n_144) );
INVx2_ASAP7_75t_SL g145 ( .A(n_25), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_10), .Y(n_146) );
CKINVDCx16_ASAP7_75t_R g147 ( .A(n_57), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_33), .Y(n_148) );
CKINVDCx8_ASAP7_75t_R g149 ( .A(n_128), .Y(n_149) );
CKINVDCx11_ASAP7_75t_R g150 ( .A(n_113), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_112), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_144), .Y(n_152) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_129), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_144), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_145), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_140), .B(n_0), .Y(n_156) );
INVx1_ASAP7_75t_SL g157 ( .A(n_131), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_145), .Y(n_158) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_112), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_112), .Y(n_160) );
NAND2xp33_ASAP7_75t_L g161 ( .A(n_106), .B(n_23), .Y(n_161) );
OAI21x1_ASAP7_75t_L g162 ( .A1(n_105), .A2(n_44), .B(n_102), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_107), .Y(n_163) );
INVxp67_ASAP7_75t_L g164 ( .A(n_104), .Y(n_164) );
OAI22xp5_ASAP7_75t_L g165 ( .A1(n_131), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_108), .Y(n_166) );
AND2x6_ASAP7_75t_L g167 ( .A(n_115), .B(n_26), .Y(n_167) );
INVx2_ASAP7_75t_SL g168 ( .A(n_151), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_163), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_163), .Y(n_170) );
NOR2xp33_ASAP7_75t_SL g171 ( .A(n_167), .B(n_147), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_163), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_163), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_159), .B(n_104), .Y(n_174) );
AND2x4_ASAP7_75t_L g175 ( .A(n_151), .B(n_118), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_151), .B(n_106), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_163), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_149), .Y(n_178) );
INVx2_ASAP7_75t_SL g179 ( .A(n_167), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_164), .B(n_119), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_166), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_166), .Y(n_182) );
INVx3_ASAP7_75t_L g183 ( .A(n_166), .Y(n_183) );
AOI22xp33_ASAP7_75t_L g184 ( .A1(n_167), .A2(n_130), .B1(n_125), .B2(n_142), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_152), .B(n_123), .Y(n_185) );
INVx4_ASAP7_75t_L g186 ( .A(n_167), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_152), .B(n_133), .Y(n_187) );
CKINVDCx6p67_ASAP7_75t_R g188 ( .A(n_167), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_166), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_166), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_153), .B(n_109), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_154), .B(n_135), .Y(n_192) );
INVx3_ASAP7_75t_L g193 ( .A(n_160), .Y(n_193) );
XNOR2xp5_ASAP7_75t_L g194 ( .A(n_178), .B(n_157), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_176), .B(n_156), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_171), .B(n_149), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_176), .B(n_154), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_193), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_186), .B(n_136), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_186), .B(n_137), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g201 ( .A1(n_184), .A2(n_126), .B1(n_121), .B2(n_158), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_171), .B(n_109), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_176), .B(n_174), .Y(n_203) );
OR2x6_ASAP7_75t_L g204 ( .A(n_191), .B(n_165), .Y(n_204) );
AOI221xp5_ASAP7_75t_L g205 ( .A1(n_174), .A2(n_146), .B1(n_141), .B2(n_116), .C(n_160), .Y(n_205) );
INVx2_ASAP7_75t_SL g206 ( .A(n_191), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_174), .B(n_155), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_180), .B(n_155), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_180), .B(n_158), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_175), .B(n_110), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_168), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g212 ( .A1(n_191), .A2(n_161), .B1(n_141), .B2(n_146), .Y(n_212) );
OAI221xp5_ASAP7_75t_L g213 ( .A1(n_185), .A2(n_161), .B1(n_138), .B2(n_148), .C(n_111), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_186), .B(n_110), .Y(n_214) );
AOI22xp33_ASAP7_75t_L g215 ( .A1(n_175), .A2(n_167), .B1(n_162), .B2(n_132), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_186), .B(n_111), .Y(n_216) );
INVx2_ASAP7_75t_SL g217 ( .A(n_175), .Y(n_217) );
BUFx12f_ASAP7_75t_SL g218 ( .A(n_175), .Y(n_218) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_186), .Y(n_219) );
INVxp67_ASAP7_75t_L g220 ( .A(n_175), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_177), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_175), .B(n_114), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_168), .B(n_114), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_178), .B(n_150), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_186), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_168), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_193), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_195), .B(n_184), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_199), .A2(n_179), .B(n_192), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_199), .A2(n_179), .B(n_192), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g231 ( .A1(n_220), .A2(n_188), .B1(n_179), .B2(n_187), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_206), .B(n_150), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_200), .A2(n_185), .B(n_187), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_203), .A2(n_188), .B1(n_193), .B2(n_132), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_203), .B(n_193), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_217), .A2(n_188), .B1(n_124), .B2(n_139), .Y(n_236) );
O2A1O1Ixp5_ASAP7_75t_SL g237 ( .A1(n_196), .A2(n_169), .B(n_170), .C(n_189), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_219), .B(n_124), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_219), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_204), .A2(n_193), .B1(n_139), .B2(n_148), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_207), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_SL g242 ( .A1(n_200), .A2(n_127), .B(n_189), .C(n_170), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_197), .Y(n_243) );
INVx3_ASAP7_75t_SL g244 ( .A(n_224), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g245 ( .A1(n_204), .A2(n_117), .B1(n_120), .B2(n_122), .Y(n_245) );
OAI21xp5_ASAP7_75t_L g246 ( .A1(n_215), .A2(n_162), .B(n_189), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_197), .A2(n_173), .B(n_182), .C(n_169), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_218), .B(n_134), .Y(n_248) );
OR2x6_ASAP7_75t_L g249 ( .A(n_204), .B(n_143), .Y(n_249) );
OA22x2_ASAP7_75t_L g250 ( .A1(n_212), .A2(n_173), .B1(n_182), .B2(n_170), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_215), .A2(n_169), .B1(n_172), .B2(n_182), .Y(n_251) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_194), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_219), .B(n_183), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_208), .B(n_183), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_209), .Y(n_255) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_219), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_214), .A2(n_173), .B(n_172), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_208), .B(n_183), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_255), .Y(n_259) );
INVx5_ASAP7_75t_L g260 ( .A(n_239), .Y(n_260) );
AO22x2_ASAP7_75t_L g261 ( .A1(n_251), .A2(n_201), .B1(n_245), .B2(n_243), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_241), .B(n_205), .Y(n_262) );
AOI221x1_ASAP7_75t_L g263 ( .A1(n_251), .A2(n_222), .B1(n_172), .B2(n_210), .C(n_211), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_232), .B(n_222), .Y(n_264) );
OAI21x1_ASAP7_75t_L g265 ( .A1(n_237), .A2(n_246), .B(n_257), .Y(n_265) );
OAI21xp5_ASAP7_75t_L g266 ( .A1(n_228), .A2(n_202), .B(n_216), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_233), .A2(n_213), .B(n_227), .C(n_198), .Y(n_267) );
AO31x2_ASAP7_75t_L g268 ( .A1(n_247), .A2(n_177), .A3(n_181), .B(n_190), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_229), .A2(n_230), .B(n_231), .Y(n_269) );
NAND3x1_ASAP7_75t_L g270 ( .A(n_248), .B(n_223), .C(n_3), .Y(n_270) );
INVx2_ASAP7_75t_SL g271 ( .A(n_244), .Y(n_271) );
AOI21x1_ASAP7_75t_L g272 ( .A1(n_246), .A2(n_226), .B(n_190), .Y(n_272) );
AO32x2_ASAP7_75t_L g273 ( .A1(n_250), .A2(n_198), .A3(n_4), .B1(n_5), .B2(n_6), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_253), .A2(n_225), .B(n_221), .Y(n_274) );
AOI21xp33_ASAP7_75t_L g275 ( .A1(n_250), .A2(n_225), .B(n_221), .Y(n_275) );
OAI22xp5_ASAP7_75t_L g276 ( .A1(n_249), .A2(n_225), .B1(n_190), .B2(n_181), .Y(n_276) );
O2A1O1Ixp5_ASAP7_75t_L g277 ( .A1(n_238), .A2(n_190), .B(n_181), .C(n_177), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_254), .A2(n_225), .B(n_181), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_240), .B(n_2), .Y(n_279) );
NOR4xp25_ASAP7_75t_L g280 ( .A(n_235), .B(n_177), .C(n_183), .D(n_6), .Y(n_280) );
AOI221xp5_ASAP7_75t_SL g281 ( .A1(n_234), .A2(n_183), .B1(n_5), .B2(n_7), .C(n_8), .Y(n_281) );
CKINVDCx20_ASAP7_75t_R g282 ( .A(n_252), .Y(n_282) );
OA21x2_ASAP7_75t_L g283 ( .A1(n_258), .A2(n_50), .B(n_101), .Y(n_283) );
OAI21x1_ASAP7_75t_L g284 ( .A1(n_272), .A2(n_236), .B(n_242), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_259), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_273), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_273), .Y(n_287) );
OAI21x1_ASAP7_75t_L g288 ( .A1(n_265), .A2(n_256), .B(n_239), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_269), .A2(n_256), .B(n_239), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_267), .A2(n_256), .B(n_249), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_278), .A2(n_249), .B(n_52), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_273), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_262), .B(n_4), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_268), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_268), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_268), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_261), .Y(n_297) );
OR2x2_ASAP7_75t_L g298 ( .A(n_280), .B(n_8), .Y(n_298) );
INVx6_ASAP7_75t_L g299 ( .A(n_260), .Y(n_299) );
OA21x2_ASAP7_75t_L g300 ( .A1(n_263), .A2(n_54), .B(n_100), .Y(n_300) );
AOI22xp5_ASAP7_75t_L g301 ( .A1(n_261), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_260), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_283), .Y(n_303) );
AOI21x1_ASAP7_75t_L g304 ( .A1(n_283), .A2(n_55), .B(n_97), .Y(n_304) );
BUFx3_ASAP7_75t_L g305 ( .A(n_260), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_288), .Y(n_306) );
OR2x6_ASAP7_75t_L g307 ( .A(n_290), .B(n_276), .Y(n_307) );
OA21x2_ASAP7_75t_L g308 ( .A1(n_303), .A2(n_281), .B(n_275), .Y(n_308) );
BUFx2_ASAP7_75t_L g309 ( .A(n_297), .Y(n_309) );
AO21x2_ASAP7_75t_L g310 ( .A1(n_294), .A2(n_280), .B(n_266), .Y(n_310) );
INVxp67_ASAP7_75t_SL g311 ( .A(n_295), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_288), .Y(n_312) );
OAI33xp33_ASAP7_75t_L g313 ( .A1(n_298), .A2(n_279), .A3(n_276), .B1(n_270), .B2(n_281), .B3(n_16), .Y(n_313) );
INVxp67_ASAP7_75t_SL g314 ( .A(n_295), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_297), .B(n_266), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_286), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_286), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_287), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_295), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_287), .B(n_271), .Y(n_320) );
AO21x2_ASAP7_75t_L g321 ( .A1(n_294), .A2(n_274), .B(n_264), .Y(n_321) );
OAI21x1_ASAP7_75t_L g322 ( .A1(n_303), .A2(n_277), .B(n_260), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_296), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_292), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_292), .Y(n_325) );
AO21x2_ASAP7_75t_L g326 ( .A1(n_303), .A2(n_11), .B(n_12), .Y(n_326) );
INVx1_ASAP7_75t_SL g327 ( .A(n_305), .Y(n_327) );
AO21x2_ASAP7_75t_L g328 ( .A1(n_296), .A2(n_12), .B(n_13), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_298), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_300), .Y(n_330) );
BUFx12f_ASAP7_75t_L g331 ( .A(n_299), .Y(n_331) );
OAI21xp5_ASAP7_75t_L g332 ( .A1(n_301), .A2(n_289), .B(n_291), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_306), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_316), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_316), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_311), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_329), .B(n_301), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_316), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_319), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_329), .B(n_285), .Y(n_340) );
NOR2x1_ASAP7_75t_L g341 ( .A(n_328), .B(n_305), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_319), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_319), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_329), .B(n_285), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_319), .B(n_300), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_323), .Y(n_346) );
BUFx2_ASAP7_75t_L g347 ( .A(n_311), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_317), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_323), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_317), .B(n_300), .Y(n_350) );
BUFx2_ASAP7_75t_L g351 ( .A(n_314), .Y(n_351) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_314), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_309), .B(n_293), .Y(n_353) );
INVx2_ASAP7_75t_SL g354 ( .A(n_323), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_323), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_306), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_317), .B(n_324), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_309), .B(n_293), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_324), .B(n_300), .Y(n_359) );
BUFx3_ASAP7_75t_L g360 ( .A(n_331), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_324), .B(n_302), .Y(n_361) );
NOR2x1_ASAP7_75t_SL g362 ( .A(n_331), .B(n_305), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_318), .Y(n_363) );
AND2x4_ASAP7_75t_SL g364 ( .A(n_307), .B(n_302), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_318), .B(n_284), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_306), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_325), .B(n_284), .Y(n_367) );
BUFx6f_ASAP7_75t_L g368 ( .A(n_306), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_312), .Y(n_369) );
AND2x4_ASAP7_75t_L g370 ( .A(n_312), .B(n_304), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_325), .B(n_304), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_310), .B(n_13), .Y(n_372) );
INVxp67_ASAP7_75t_SL g373 ( .A(n_312), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_310), .B(n_14), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_310), .B(n_16), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_312), .Y(n_376) );
NAND4xp25_ASAP7_75t_L g377 ( .A(n_372), .B(n_320), .C(n_309), .D(n_332), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_334), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_334), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_335), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_340), .B(n_320), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_352), .B(n_320), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_335), .Y(n_383) );
BUFx3_ASAP7_75t_L g384 ( .A(n_360), .Y(n_384) );
AOI22xp33_ASAP7_75t_SL g385 ( .A1(n_360), .A2(n_327), .B1(n_331), .B2(n_328), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_342), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_357), .B(n_310), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_338), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_342), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_352), .B(n_310), .Y(n_390) );
CKINVDCx16_ASAP7_75t_R g391 ( .A(n_360), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_336), .B(n_315), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_357), .B(n_321), .Y(n_393) );
INVxp67_ASAP7_75t_L g394 ( .A(n_362), .Y(n_394) );
NOR2x1_ASAP7_75t_L g395 ( .A(n_341), .B(n_328), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_357), .B(n_321), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_336), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_347), .B(n_315), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_338), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_348), .Y(n_400) );
INVx5_ASAP7_75t_L g401 ( .A(n_347), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_342), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_340), .B(n_344), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_340), .B(n_321), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_344), .B(n_327), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_344), .B(n_321), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_343), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_348), .B(n_321), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_363), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_363), .Y(n_410) );
BUFx2_ASAP7_75t_SL g411 ( .A(n_351), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_361), .B(n_328), .Y(n_412) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_351), .B(n_331), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_361), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_361), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_354), .B(n_328), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_362), .B(n_282), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_354), .B(n_330), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_354), .B(n_330), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_353), .B(n_326), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_346), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_355), .B(n_330), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_355), .B(n_330), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_339), .B(n_326), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_339), .B(n_372), .Y(n_425) );
INVx3_ASAP7_75t_L g426 ( .A(n_333), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_346), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_346), .Y(n_428) );
BUFx3_ASAP7_75t_L g429 ( .A(n_339), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_343), .Y(n_430) );
BUFx2_ASAP7_75t_L g431 ( .A(n_339), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_353), .B(n_326), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_372), .B(n_326), .Y(n_433) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_343), .Y(n_434) );
INVxp67_ASAP7_75t_SL g435 ( .A(n_341), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_353), .B(n_326), .Y(n_436) );
BUFx2_ASAP7_75t_SL g437 ( .A(n_349), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_374), .B(n_307), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_349), .Y(n_439) );
NOR2x1_ASAP7_75t_L g440 ( .A(n_374), .B(n_332), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_349), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_374), .B(n_308), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_358), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_403), .B(n_375), .Y(n_444) );
INVxp67_ASAP7_75t_L g445 ( .A(n_411), .Y(n_445) );
AND2x4_ASAP7_75t_L g446 ( .A(n_425), .B(n_364), .Y(n_446) );
BUFx2_ASAP7_75t_L g447 ( .A(n_391), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_409), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_403), .B(n_364), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_404), .B(n_365), .Y(n_450) );
INVxp67_ASAP7_75t_L g451 ( .A(n_411), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_443), .B(n_382), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_404), .B(n_365), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_406), .B(n_365), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_409), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_377), .A2(n_337), .B1(n_375), .B2(n_358), .Y(n_456) );
AND2x4_ASAP7_75t_SL g457 ( .A(n_397), .B(n_375), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_410), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_410), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_406), .B(n_367), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_393), .B(n_367), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_393), .B(n_367), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_396), .B(n_350), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_391), .B(n_394), .Y(n_464) );
AND2x2_ASAP7_75t_SL g465 ( .A(n_431), .B(n_358), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_378), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_378), .Y(n_467) );
NAND2x1_ASAP7_75t_L g468 ( .A(n_431), .B(n_337), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_414), .B(n_337), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_396), .B(n_359), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_379), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_414), .B(n_364), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_379), .Y(n_473) );
OAI21xp5_ASAP7_75t_SL g474 ( .A1(n_417), .A2(n_359), .B(n_350), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_415), .B(n_359), .Y(n_475) );
AOI211xp5_ASAP7_75t_L g476 ( .A1(n_413), .A2(n_313), .B(n_350), .C(n_371), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_425), .B(n_371), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_387), .B(n_371), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_387), .B(n_345), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_380), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_386), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_415), .B(n_345), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_380), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_386), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_383), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_389), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_383), .Y(n_487) );
OAI21xp33_ASAP7_75t_L g488 ( .A1(n_440), .A2(n_307), .B(n_345), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_388), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_438), .B(n_307), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_438), .B(n_376), .Y(n_491) );
INVx1_ASAP7_75t_SL g492 ( .A(n_384), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_389), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_388), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_402), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_412), .B(n_376), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_412), .B(n_376), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_381), .B(n_366), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_399), .B(n_366), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_440), .A2(n_313), .B1(n_307), .B2(n_368), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_402), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_384), .B(n_17), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_399), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_400), .B(n_366), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_400), .Y(n_505) );
NAND3xp33_ASAP7_75t_L g506 ( .A(n_385), .B(n_333), .C(n_368), .Y(n_506) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_434), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_408), .B(n_356), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_382), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_408), .B(n_356), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_407), .Y(n_511) );
INVxp67_ASAP7_75t_L g512 ( .A(n_437), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_424), .B(n_356), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_405), .B(n_369), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_392), .Y(n_515) );
INVx1_ASAP7_75t_SL g516 ( .A(n_437), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_392), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_424), .B(n_369), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_398), .Y(n_519) );
INVxp67_ASAP7_75t_L g520 ( .A(n_398), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_407), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_420), .B(n_369), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_433), .B(n_308), .Y(n_523) );
INVx3_ASAP7_75t_SL g524 ( .A(n_401), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_420), .B(n_373), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_421), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_461), .B(n_401), .Y(n_527) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_507), .Y(n_528) );
AOI21xp33_ASAP7_75t_L g529 ( .A1(n_502), .A2(n_435), .B(n_390), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_515), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_517), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_461), .B(n_401), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_462), .B(n_401), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_478), .B(n_390), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_478), .B(n_432), .Y(n_535) );
NOR3xp33_ASAP7_75t_L g536 ( .A(n_502), .B(n_395), .C(n_442), .Y(n_536) );
NAND2x1_ASAP7_75t_SL g537 ( .A(n_524), .B(n_395), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_519), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_452), .B(n_432), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_509), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_462), .B(n_401), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_506), .A2(n_401), .B(n_373), .Y(n_542) );
OAI21xp5_ASAP7_75t_SL g543 ( .A1(n_456), .A2(n_436), .B(n_416), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_463), .B(n_436), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_507), .Y(n_545) );
INVx1_ASAP7_75t_SL g546 ( .A(n_447), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_481), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_481), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_463), .B(n_421), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_520), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_450), .B(n_429), .Y(n_551) );
NOR2x1_ASAP7_75t_L g552 ( .A(n_492), .B(n_429), .Y(n_552) );
INVx2_ASAP7_75t_SL g553 ( .A(n_449), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_450), .B(n_453), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_484), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_470), .B(n_428), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_453), .B(n_429), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_454), .B(n_416), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_448), .Y(n_559) );
OR2x6_ASAP7_75t_L g560 ( .A(n_468), .B(n_419), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_455), .Y(n_561) );
AND2x4_ASAP7_75t_L g562 ( .A(n_446), .B(n_419), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_454), .B(n_428), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_458), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_470), .B(n_427), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_460), .B(n_427), .Y(n_566) );
INVxp67_ASAP7_75t_L g567 ( .A(n_526), .Y(n_567) );
NAND2x1p5_ASAP7_75t_L g568 ( .A(n_516), .B(n_418), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_484), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_460), .B(n_430), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_491), .B(n_479), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_459), .Y(n_572) );
INVxp67_ASAP7_75t_SL g573 ( .A(n_486), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_466), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_467), .Y(n_575) );
INVxp67_ASAP7_75t_SL g576 ( .A(n_486), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_471), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_473), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_464), .B(n_17), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_444), .B(n_430), .Y(n_580) );
AND2x4_ASAP7_75t_SL g581 ( .A(n_464), .B(n_441), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_469), .B(n_18), .Y(n_582) );
AND2x4_ASAP7_75t_L g583 ( .A(n_446), .B(n_418), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_491), .B(n_423), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_475), .B(n_441), .Y(n_585) );
INVx1_ASAP7_75t_SL g586 ( .A(n_524), .Y(n_586) );
OAI31xp33_ASAP7_75t_L g587 ( .A1(n_457), .A2(n_423), .A3(n_422), .B(n_426), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_479), .B(n_439), .Y(n_588) );
OAI21xp5_ASAP7_75t_L g589 ( .A1(n_465), .A2(n_307), .B(n_426), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_493), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_510), .B(n_439), .Y(n_591) );
AND2x4_ASAP7_75t_SL g592 ( .A(n_446), .B(n_422), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_510), .B(n_426), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_474), .B(n_426), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_480), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_457), .B(n_307), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_493), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_496), .B(n_368), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_445), .B(n_19), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_495), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_495), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_501), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_465), .A2(n_299), .B1(n_368), .B2(n_333), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_534), .B(n_508), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_534), .B(n_482), .Y(n_605) );
OAI21xp5_ASAP7_75t_SL g606 ( .A1(n_587), .A2(n_451), .B(n_500), .Y(n_606) );
OAI322xp33_ASAP7_75t_L g607 ( .A1(n_546), .A2(n_525), .A3(n_498), .B1(n_523), .B2(n_514), .C1(n_472), .C2(n_512), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_567), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_550), .B(n_477), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_560), .A2(n_500), .B1(n_476), .B2(n_477), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_554), .B(n_477), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_567), .Y(n_612) );
AOI221xp5_ASAP7_75t_L g613 ( .A1(n_543), .A2(n_488), .B1(n_487), .B2(n_489), .C(n_494), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_592), .B(n_490), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_528), .Y(n_615) );
OAI221xp5_ASAP7_75t_L g616 ( .A1(n_536), .A2(n_483), .B1(n_485), .B2(n_503), .C(n_505), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_540), .B(n_522), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_530), .B(n_496), .Y(n_618) );
OAI221xp5_ASAP7_75t_L g619 ( .A1(n_536), .A2(n_579), .B1(n_529), .B2(n_560), .C(n_599), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_531), .B(n_497), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_538), .B(n_497), .Y(n_621) );
AOI21xp33_ASAP7_75t_L g622 ( .A1(n_582), .A2(n_504), .B(n_499), .Y(n_622) );
NAND2x1_ASAP7_75t_L g623 ( .A(n_560), .B(n_511), .Y(n_623) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_545), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_549), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_535), .B(n_513), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_571), .B(n_518), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g628 ( .A(n_552), .B(n_521), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_535), .B(n_513), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_544), .B(n_518), .Y(n_630) );
BUFx2_ASAP7_75t_L g631 ( .A(n_568), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_549), .Y(n_632) );
OAI211xp5_ASAP7_75t_L g633 ( .A1(n_529), .A2(n_521), .B(n_511), .C(n_501), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_556), .Y(n_634) );
OAI21xp5_ASAP7_75t_L g635 ( .A1(n_568), .A2(n_370), .B(n_322), .Y(n_635) );
OAI211xp5_ASAP7_75t_SL g636 ( .A1(n_589), .A2(n_20), .B(n_21), .C(n_22), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_594), .A2(n_368), .B1(n_333), .B2(n_370), .C(n_20), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_556), .Y(n_638) );
NOR2xp67_ASAP7_75t_L g639 ( .A(n_542), .B(n_21), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_588), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_565), .Y(n_641) );
CKINVDCx16_ASAP7_75t_R g642 ( .A(n_553), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_547), .Y(n_643) );
INVx2_ASAP7_75t_SL g644 ( .A(n_581), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_586), .A2(n_299), .B1(n_368), .B2(n_333), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_565), .B(n_299), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_562), .B(n_368), .Y(n_647) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_573), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_594), .A2(n_333), .B1(n_370), .B2(n_308), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_562), .A2(n_333), .B1(n_370), .B2(n_308), .Y(n_650) );
OAI21xp5_ASAP7_75t_L g651 ( .A1(n_542), .A2(n_370), .B(n_322), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_527), .A2(n_308), .B1(n_322), .B2(n_31), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_596), .A2(n_308), .B1(n_29), .B2(n_32), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_642), .B(n_603), .Y(n_654) );
OAI21xp5_ASAP7_75t_SL g655 ( .A1(n_619), .A2(n_532), .B(n_533), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_625), .Y(n_656) );
NAND4xp25_ASAP7_75t_L g657 ( .A(n_619), .B(n_541), .C(n_544), .D(n_539), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_632), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_644), .B(n_583), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_634), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_638), .Y(n_661) );
OAI32xp33_ASAP7_75t_L g662 ( .A1(n_648), .A2(n_563), .A3(n_566), .B1(n_570), .B2(n_585), .Y(n_662) );
OAI22xp33_ASAP7_75t_SL g663 ( .A1(n_623), .A2(n_583), .B1(n_566), .B2(n_573), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_641), .Y(n_664) );
NOR3xp33_ASAP7_75t_L g665 ( .A(n_636), .B(n_575), .C(n_559), .Y(n_665) );
OAI21xp5_ASAP7_75t_L g666 ( .A1(n_639), .A2(n_537), .B(n_576), .Y(n_666) );
OAI22xp33_ASAP7_75t_L g667 ( .A1(n_610), .A2(n_570), .B1(n_585), .B2(n_598), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_606), .A2(n_551), .B1(n_557), .B2(n_593), .Y(n_668) );
NOR3x1_ASAP7_75t_L g669 ( .A(n_631), .B(n_593), .C(n_598), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_608), .Y(n_670) );
NOR3xp33_ASAP7_75t_L g671 ( .A(n_636), .B(n_577), .C(n_561), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_612), .Y(n_672) );
O2A1O1Ixp5_ASAP7_75t_L g673 ( .A1(n_628), .A2(n_576), .B(n_564), .C(n_572), .Y(n_673) );
AOI221xp5_ASAP7_75t_L g674 ( .A1(n_607), .A2(n_574), .B1(n_578), .B2(n_595), .C(n_591), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_618), .Y(n_675) );
AOI32xp33_ASAP7_75t_L g676 ( .A1(n_613), .A2(n_558), .A3(n_584), .B1(n_591), .B2(n_580), .Y(n_676) );
A2O1A1Ixp33_ASAP7_75t_L g677 ( .A1(n_613), .A2(n_602), .B(n_601), .C(n_600), .Y(n_677) );
OAI221xp5_ASAP7_75t_L g678 ( .A1(n_616), .A2(n_597), .B1(n_590), .B2(n_569), .C(n_555), .Y(n_678) );
OAI211xp5_ASAP7_75t_L g679 ( .A1(n_637), .A2(n_548), .B(n_35), .C(n_36), .Y(n_679) );
OAI32xp33_ASAP7_75t_L g680 ( .A1(n_616), .A2(n_28), .A3(n_37), .B1(n_39), .B2(n_40), .Y(n_680) );
NAND2xp5_ASAP7_75t_SL g681 ( .A(n_637), .B(n_41), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_646), .A2(n_42), .B1(n_45), .B2(n_47), .Y(n_682) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_622), .A2(n_49), .B1(n_58), .B2(n_59), .C(n_61), .Y(n_683) );
AOI311xp33_ASAP7_75t_L g684 ( .A1(n_609), .A2(n_66), .A3(n_68), .B(n_72), .C(n_73), .Y(n_684) );
NOR2x1_ASAP7_75t_L g685 ( .A(n_633), .B(n_74), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_633), .A2(n_75), .B(n_77), .Y(n_686) );
OAI31xp33_ASAP7_75t_L g687 ( .A1(n_615), .A2(n_79), .A3(n_81), .B(n_83), .Y(n_687) );
NAND3xp33_ASAP7_75t_L g688 ( .A(n_651), .B(n_84), .C(n_85), .Y(n_688) );
AOI211xp5_ASAP7_75t_L g689 ( .A1(n_650), .A2(n_86), .B(n_91), .C(n_92), .Y(n_689) );
OAI21xp33_ASAP7_75t_L g690 ( .A1(n_617), .A2(n_94), .B(n_103), .Y(n_690) );
XNOR2x1_ASAP7_75t_L g691 ( .A(n_614), .B(n_605), .Y(n_691) );
AOI221x1_ASAP7_75t_L g692 ( .A1(n_645), .A2(n_635), .B1(n_611), .B2(n_620), .C(n_621), .Y(n_692) );
OAI221xp5_ASAP7_75t_L g693 ( .A1(n_649), .A2(n_653), .B1(n_604), .B2(n_626), .C(n_630), .Y(n_693) );
AOI222xp33_ASAP7_75t_L g694 ( .A1(n_624), .A2(n_629), .B1(n_640), .B2(n_627), .C1(n_647), .C2(n_643), .Y(n_694) );
NOR2x1_ASAP7_75t_L g695 ( .A(n_685), .B(n_679), .Y(n_695) );
NOR2xp67_ASAP7_75t_L g696 ( .A(n_657), .B(n_655), .Y(n_696) );
NOR3xp33_ASAP7_75t_L g697 ( .A(n_667), .B(n_674), .C(n_679), .Y(n_697) );
AOI211xp5_ASAP7_75t_L g698 ( .A1(n_663), .A2(n_674), .B(n_681), .C(n_654), .Y(n_698) );
NOR2xp67_ASAP7_75t_L g699 ( .A(n_668), .B(n_678), .Y(n_699) );
NOR4xp25_ASAP7_75t_L g700 ( .A(n_676), .B(n_677), .C(n_670), .D(n_672), .Y(n_700) );
O2A1O1Ixp33_ASAP7_75t_L g701 ( .A1(n_673), .A2(n_662), .B(n_665), .C(n_671), .Y(n_701) );
NAND3xp33_ASAP7_75t_L g702 ( .A(n_698), .B(n_692), .C(n_683), .Y(n_702) );
AND2x4_ASAP7_75t_L g703 ( .A(n_696), .B(n_659), .Y(n_703) );
NAND3x1_ASAP7_75t_L g704 ( .A(n_697), .B(n_666), .C(n_686), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_695), .Y(n_705) );
OR2x2_ASAP7_75t_L g706 ( .A(n_705), .B(n_700), .Y(n_706) );
NAND2xp33_ASAP7_75t_SL g707 ( .A(n_703), .B(n_691), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_702), .B(n_699), .Y(n_708) );
AOI211xp5_ASAP7_75t_L g709 ( .A1(n_707), .A2(n_701), .B(n_704), .C(n_680), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_708), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_710), .Y(n_711) );
AO22x1_ASAP7_75t_L g712 ( .A1(n_709), .A2(n_706), .B1(n_669), .B2(n_658), .Y(n_712) );
OAI22x1_ASAP7_75t_L g713 ( .A1(n_711), .A2(n_712), .B1(n_682), .B2(n_688), .Y(n_713) );
AOI22x1_ASAP7_75t_L g714 ( .A1(n_711), .A2(n_694), .B1(n_675), .B2(n_660), .Y(n_714) );
AOI21xp33_ASAP7_75t_L g715 ( .A1(n_713), .A2(n_687), .B(n_693), .Y(n_715) );
AOI21xp5_ASAP7_75t_SL g716 ( .A1(n_715), .A2(n_714), .B(n_656), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_716), .A2(n_661), .B1(n_664), .B2(n_689), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_717), .A2(n_690), .B1(n_652), .B2(n_684), .Y(n_718) );
endmodule