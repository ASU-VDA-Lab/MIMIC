module fake_jpeg_14832_n_244 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_244);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_244;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_22),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_34),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_40),
.Y(n_56)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_39),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_23),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_37),
.A2(n_18),
.B1(n_21),
.B2(n_32),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_44),
.A2(n_46),
.B1(n_52),
.B2(n_1),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_18),
.B1(n_21),
.B2(n_32),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_31),
.B1(n_23),
.B2(n_30),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_57),
.B1(n_39),
.B2(n_38),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_49),
.B(n_34),
.Y(n_71)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_31),
.B1(n_30),
.B2(n_27),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_27),
.B1(n_28),
.B2(n_19),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_65),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_33),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_63),
.A2(n_59),
.B(n_25),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_64),
.A2(n_79),
.B1(n_43),
.B2(n_50),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_48),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_38),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_80),
.C(n_59),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_70),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_34),
.Y(n_70)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_26),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_25),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_46),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_74),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_54),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_52),
.B(n_60),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_75),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_76),
.B(n_2),
.Y(n_105)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_39),
.B1(n_43),
.B2(n_50),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_26),
.C(n_25),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_49),
.B(n_26),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_81),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_82),
.Y(n_95)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_79),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_17),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_90),
.B(n_105),
.Y(n_112)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

AND2x6_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_1),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_92),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_63),
.B(n_80),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_100),
.B(n_96),
.Y(n_118)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_101),
.A2(n_107),
.B1(n_43),
.B2(n_58),
.Y(n_126)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_58),
.B1(n_51),
.B2(n_38),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_45),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_77),
.Y(n_119)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_72),
.C(n_77),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_93),
.C(n_100),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_124),
.B1(n_97),
.B2(n_94),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_96),
.B(n_63),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_115),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_94),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_83),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_117),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_119),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_99),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_126),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_127),
.A2(n_122),
.B1(n_123),
.B2(n_111),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_131),
.B1(n_107),
.B2(n_102),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_98),
.A2(n_76),
.B1(n_64),
.B2(n_45),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_129),
.A2(n_105),
.B1(n_92),
.B2(n_95),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_83),
.Y(n_130)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_51),
.Y(n_132)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_140),
.C(n_145),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_85),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_134),
.A2(n_136),
.B1(n_146),
.B2(n_128),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_85),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_138),
.A2(n_153),
.B1(n_112),
.B2(n_110),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_97),
.C(n_99),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_144),
.A2(n_149),
.B1(n_151),
.B2(n_67),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_95),
.C(n_106),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_123),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_87),
.B1(n_106),
.B2(n_35),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_128),
.A2(n_26),
.B(n_87),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_150),
.A2(n_120),
.B(n_42),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_114),
.A2(n_42),
.B1(n_35),
.B2(n_36),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_129),
.A2(n_42),
.B1(n_35),
.B2(n_82),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_125),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_124),
.Y(n_157)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_156),
.Y(n_160)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_164),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_140),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_175),
.C(n_177),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_120),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_162),
.B(n_166),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_118),
.Y(n_163)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_163),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_142),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_165),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_181)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_120),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_170),
.A2(n_171),
.B(n_136),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_155),
.A2(n_127),
.B1(n_116),
.B2(n_111),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_172),
.A2(n_144),
.B1(n_148),
.B2(n_152),
.Y(n_180)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_173),
.A2(n_174),
.B1(n_135),
.B2(n_155),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_116),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_121),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_176),
.A2(n_170),
.B1(n_134),
.B2(n_135),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_121),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_152),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_24),
.C(n_20),
.Y(n_204)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_189),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_183),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_161),
.B(n_146),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_164),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_170),
.A2(n_136),
.B(n_143),
.Y(n_185)
);

XOR2x1_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_134),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_153),
.B1(n_121),
.B2(n_28),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_159),
.A2(n_19),
.B1(n_67),
.B2(n_82),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_191),
.B(n_172),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_158),
.A2(n_67),
.B1(n_3),
.B2(n_4),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_2),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_196),
.A2(n_201),
.B1(n_179),
.B2(n_188),
.Y(n_214)
);

OAI31xp33_ASAP7_75t_SL g197 ( 
.A1(n_183),
.A2(n_171),
.A3(n_175),
.B(n_158),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_198),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_194),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_203),
.C(n_207),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_202),
.B(n_185),
.Y(n_212)
);

OAI311xp33_ASAP7_75t_L g203 ( 
.A1(n_178),
.A2(n_17),
.A3(n_20),
.B1(n_4),
.C1(n_5),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_3),
.C(n_4),
.Y(n_217)
);

MAJx2_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_187),
.C(n_190),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_205),
.A2(n_180),
.B(n_17),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_24),
.C(n_17),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_192),
.C(n_193),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_213),
.C(n_215),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_206),
.B(n_190),
.Y(n_211)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_211),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_212),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_205),
.C(n_204),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_216),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_2),
.C(n_3),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_201),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_220),
.B(n_221),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_211),
.A2(n_200),
.B1(n_207),
.B2(n_195),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_208),
.A2(n_197),
.B1(n_7),
.B2(n_8),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_222),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_208),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_223),
.B(n_209),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_227),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_6),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_224),
.B(n_7),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_230),
.B(n_231),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_218),
.B(n_10),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_228),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_232),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_228),
.A2(n_10),
.B(n_11),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_235),
.A2(n_236),
.B1(n_12),
.B2(n_13),
.Y(n_238)
);

NOR2xp67_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_11),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_234),
.B(n_232),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_237),
.A2(n_233),
.B(n_14),
.Y(n_240)
);

BUFx24_ASAP7_75t_SL g241 ( 
.A(n_238),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_240),
.Y(n_242)
);

OAI321xp33_ASAP7_75t_L g243 ( 
.A1(n_242),
.A2(n_241),
.A3(n_239),
.B1(n_15),
.B2(n_14),
.C(n_12),
.Y(n_243)
);

XNOR2x2_ASAP7_75t_SL g244 ( 
.A(n_243),
.B(n_15),
.Y(n_244)
);


endmodule