module real_jpeg_26481_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_0),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_0),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_0),
.B(n_85),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_2),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_2),
.B(n_100),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_2),
.B(n_85),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_2),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_2),
.B(n_34),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_2),
.B(n_52),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_2),
.B(n_38),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_3),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_3),
.B(n_85),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_3),
.B(n_96),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_3),
.B(n_60),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_3),
.B(n_49),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_3),
.B(n_34),
.Y(n_227)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_3),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_3),
.B(n_203),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_5),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_5),
.B(n_60),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_5),
.B(n_100),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_5),
.B(n_108),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_5),
.B(n_49),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_5),
.B(n_34),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_5),
.B(n_52),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_5),
.B(n_203),
.Y(n_261)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_6),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_7),
.Y(n_101)
);

INVx8_ASAP7_75t_SL g28 ( 
.A(n_8),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_9),
.B(n_49),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_9),
.B(n_34),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_9),
.B(n_60),
.Y(n_129)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_9),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_9),
.B(n_100),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_9),
.B(n_52),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_10),
.B(n_38),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_10),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_10),
.B(n_100),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_10),
.B(n_85),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_10),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_10),
.B(n_49),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_10),
.B(n_34),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_11),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_11),
.B(n_52),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_11),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_11),
.B(n_100),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_11),
.B(n_85),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_11),
.B(n_60),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_11),
.B(n_49),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_11),
.B(n_34),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_12),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_12),
.B(n_100),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_12),
.B(n_85),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_12),
.B(n_60),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_12),
.B(n_49),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_12),
.B(n_34),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_12),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_12),
.B(n_203),
.Y(n_333)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_15),
.B(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_15),
.B(n_197),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_15),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_15),
.B(n_85),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_15),
.B(n_60),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_15),
.B(n_49),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_15),
.B(n_34),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_15),
.B(n_52),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_16),
.B(n_60),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_16),
.B(n_49),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_16),
.B(n_85),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_16),
.B(n_100),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_16),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_16),
.B(n_34),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_16),
.B(n_52),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_16),
.B(n_203),
.Y(n_243)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_17),
.Y(n_97)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_17),
.Y(n_109)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_17),
.Y(n_145)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_17),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_65),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_41),
.B2(n_42),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_32),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx11_ASAP7_75t_L g203 ( 
.A(n_25),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_26),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_SL g32 ( 
.A(n_26),
.B(n_33),
.C(n_37),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_26),
.A2(n_31),
.B1(n_33),
.B2(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_27),
.B(n_257),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_27),
.B(n_288),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_27),
.B(n_252),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_29),
.B(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_29),
.B(n_266),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_29),
.B(n_239),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_62),
.C(n_63),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_43),
.B(n_391),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_54),
.C(n_55),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_44),
.B(n_389),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_51),
.B2(n_53),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g379 ( 
.A1(n_47),
.A2(n_48),
.B1(n_58),
.B2(n_347),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_56),
.C(n_58),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_50),
.C(n_53),
.Y(n_62)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_49),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_51),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_54),
.B(n_55),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_56),
.A2(n_57),
.B1(n_379),
.B2(n_380),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_58),
.A2(n_319),
.B1(n_320),
.B2(n_347),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_58),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_SL g377 ( 
.A(n_58),
.B(n_320),
.C(n_345),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_59),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_59),
.B(n_252),
.Y(n_251)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_62),
.B(n_63),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_390),
.C(n_392),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_384),
.C(n_385),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_366),
.C(n_367),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_337),
.C(n_338),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_312),
.C(n_313),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_280),
.C(n_281),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_245),
.C(n_246),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_209),
.C(n_210),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_176),
.C(n_177),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_150),
.C(n_151),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_111),
.C(n_122),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_92),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_87),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_78),
.B(n_87),
.C(n_92),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_81),
.C(n_83),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_79),
.A2(n_80),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

BUFx24_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_88),
.B(n_90),
.C(n_91),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_102),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_93),
.B(n_103),
.C(n_104),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_98),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_94),
.A2(n_95),
.B1(n_98),
.B2(n_99),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_97),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_100),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_107),
.B2(n_110),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_105),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_106),
.B(n_110),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_109),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_115),
.C(n_121),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_115),
.A2(n_116),
.B1(n_121),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_119),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_146),
.C(n_147),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_131),
.C(n_136),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_129),
.C(n_130),
.Y(n_146)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.C(n_141),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_139),
.B(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_165),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_166),
.C(n_175),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_161),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_160),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_160),
.C(n_161),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_155),
.Y(n_159)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_156),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_159),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx24_ASAP7_75t_SL g393 ( 
.A(n_161),
.Y(n_393)
);

FAx1_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_163),
.CI(n_164),
.CON(n_161),
.SN(n_161)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_163),
.C(n_164),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_175),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_173),
.B2(n_174),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_169),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_172),
.C(n_174),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_173),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_192),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_181),
.C(n_192),
.Y(n_209)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_187),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_188),
.C(n_191),
.Y(n_213)
);

BUFx24_ASAP7_75t_SL g397 ( 
.A(n_183),
.Y(n_397)
);

FAx1_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_185),
.CI(n_186),
.CON(n_183),
.SN(n_183)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_184),
.B(n_185),
.C(n_186),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_193),
.B(n_200),
.C(n_207),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_200),
.B1(n_207),
.B2(n_208),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_195),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_198),
.B(n_199),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_198),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_234),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_199),
.B(n_234),
.C(n_235),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_200),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_205),
.C(n_206),
.Y(n_229)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_230),
.B2(n_244),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_211),
.B(n_231),
.C(n_232),
.Y(n_245)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_215),
.C(n_223),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_223),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_216),
.B(n_219),
.C(n_222),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_255),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_221),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_229),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_225),
.B(n_228),
.C(n_229),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_227),
.Y(n_228)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_230),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_236),
.B(n_275),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_236),
.B(n_276),
.C(n_277),
.Y(n_301)
);

FAx1_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_240),
.CI(n_243),
.CON(n_236),
.SN(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_278),
.B2(n_279),
.Y(n_246)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_247),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_248),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_270),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_249),
.B(n_270),
.C(n_278),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_258),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_250),
.B(n_259),
.C(n_260),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_251),
.B(n_254),
.C(n_256),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_263),
.B2(n_269),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_261),
.Y(n_269)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_267),
.B2(n_268),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_265),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_264),
.B(n_268),
.C(n_269),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_264),
.B(n_287),
.C(n_290),
.Y(n_335)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_273),
.C(n_274),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_282),
.B(n_284),
.C(n_311),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_298),
.B2(n_311),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_292),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_286),
.B(n_293),
.C(n_294),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_289),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_290),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_290),
.A2(n_291),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_SL g351 ( 
.A(n_290),
.B(n_317),
.C(n_320),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

BUFx24_ASAP7_75t_SL g395 ( 
.A(n_294),
.Y(n_395)
);

FAx1_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_296),
.CI(n_297),
.CON(n_294),
.SN(n_294)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_295),
.B(n_296),
.C(n_297),
.Y(n_322)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_298),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_299),
.B(n_301),
.C(n_302),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_305),
.B2(n_310),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_306),
.C(n_308),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_305),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_306),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_307),
.A2(n_308),
.B1(n_333),
.B2(n_334),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_308),
.B(n_334),
.C(n_335),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_336),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_327),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_315),
.B(n_327),
.C(n_336),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_321),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_316),
.B(n_322),
.C(n_323),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

BUFx24_ASAP7_75t_SL g396 ( 
.A(n_323),
.Y(n_396)
);

FAx1_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_325),
.CI(n_326),
.CON(n_323),
.SN(n_323)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_324),
.B(n_325),
.C(n_326),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_330),
.C(n_331),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_335),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_333),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_339),
.B(n_341),
.C(n_353),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_342),
.B1(n_352),
.B2(n_353),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_343),
.A2(n_344),
.B1(n_348),
.B2(n_349),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_343),
.B(n_350),
.C(n_351),
.Y(n_369)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_354),
.B(n_356),
.C(n_359),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_356),
.A2(n_357),
.B1(n_358),
.B2(n_359),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_359),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_360),
.B(n_362),
.C(n_365),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_363),
.B1(n_364),
.B2(n_365),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_363),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_364),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_368),
.A2(n_381),
.B1(n_382),
.B2(n_383),
.Y(n_367)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_368),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_369),
.B(n_370),
.C(n_383),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_376),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_371),
.B(n_377),
.C(n_378),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_372),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_372),
.B(n_388),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_372),
.B(n_386),
.C(n_388),
.Y(n_392)
);

FAx1_ASAP7_75t_SL g372 ( 
.A(n_373),
.B(n_374),
.CI(n_375),
.CON(n_372),
.SN(n_372)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_378),
.Y(n_376)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_379),
.Y(n_380)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_381),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);


endmodule