module fake_jpeg_3426_n_229 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_229);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_6),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_52),
.Y(n_58)
);

BUFx8_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_10),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_18),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_25),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_21),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_28),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_35),
.Y(n_69)
);

BUFx4f_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_15),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_9),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_30),
.Y(n_74)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_36),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_54),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_77),
.B1(n_72),
.B2(n_78),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_70),
.B1(n_78),
.B2(n_57),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_55),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_100),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_61),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_97),
.B(n_98),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_63),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_71),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_72),
.B(n_57),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_86),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_99),
.A2(n_102),
.B1(n_88),
.B2(n_101),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_112),
.B1(n_113),
.B2(n_56),
.Y(n_125)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_81),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_114),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_70),
.B1(n_56),
.B2(n_80),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_81),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_118),
.Y(n_128)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_121),
.B(n_122),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_97),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_70),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_123),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_125),
.A2(n_105),
.B1(n_62),
.B2(n_67),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_80),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_135),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_104),
.A2(n_79),
.B1(n_73),
.B2(n_58),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_68),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_115),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_139),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_113),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_120),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_109),
.B(n_64),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_140),
.B(n_74),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_76),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_65),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_146),
.A2(n_163),
.B1(n_170),
.B2(n_145),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_119),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_150),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_128),
.A2(n_79),
.B1(n_67),
.B2(n_62),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_149),
.A2(n_160),
.B1(n_162),
.B2(n_168),
.Y(n_182)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_124),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_153),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_159),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_75),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_156),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_69),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_155),
.B(n_157),
.Y(n_171)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_144),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_66),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_131),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_142),
.B(n_0),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_161),
.B(n_164),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_137),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_4),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_129),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_33),
.Y(n_189)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_137),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_7),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_169),
.B(n_49),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_141),
.A2(n_24),
.B1(n_47),
.B2(n_45),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_153),
.C(n_165),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_174),
.C(n_187),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_129),
.C(n_132),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_176),
.A2(n_12),
.B(n_13),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_145),
.Y(n_177)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_148),
.A2(n_132),
.B(n_23),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_SL g202 ( 
.A1(n_178),
.A2(n_181),
.B(n_32),
.C(n_31),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_159),
.A2(n_22),
.B1(n_43),
.B2(n_42),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_147),
.Y(n_184)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_149),
.B(n_37),
.C(n_34),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_168),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_8),
.Y(n_195)
);

AOI221xp5_ASAP7_75t_L g193 ( 
.A1(n_172),
.A2(n_170),
.B1(n_9),
.B2(n_10),
.C(n_11),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_R g207 ( 
.A(n_193),
.B(n_199),
.C(n_187),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_195),
.B(n_200),
.Y(n_204)
);

FAx1_ASAP7_75t_SL g199 ( 
.A(n_174),
.B(n_11),
.CI(n_12),
.CON(n_199),
.SN(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_186),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_201),
.A2(n_181),
.B1(n_182),
.B2(n_175),
.Y(n_205)
);

NOR2xp67_ASAP7_75t_SL g211 ( 
.A(n_202),
.B(n_26),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_192),
.A2(n_173),
.B1(n_178),
.B2(n_182),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_203),
.B(n_205),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_183),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_196),
.C(n_198),
.Y(n_214)
);

NOR3xp33_ASAP7_75t_SL g212 ( 
.A(n_207),
.B(n_210),
.C(n_194),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_197),
.A2(n_177),
.B1(n_180),
.B2(n_179),
.Y(n_208)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_208),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_171),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_209),
.A2(n_211),
.B(n_202),
.Y(n_217)
);

NOR3xp33_ASAP7_75t_SL g210 ( 
.A(n_199),
.B(n_29),
.C(n_27),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_217),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_215),
.C(n_193),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_209),
.B(n_204),
.Y(n_215)
);

OAI21x1_ASAP7_75t_L g223 ( 
.A1(n_218),
.A2(n_219),
.B(n_221),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_213),
.A2(n_210),
.B(n_202),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_216),
.A2(n_13),
.B(n_14),
.Y(n_221)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_220),
.Y(n_222)
);

OAI21xp33_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_216),
.B(n_16),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_14),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_225),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_226),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_227),
.A2(n_223),
.B1(n_18),
.B2(n_19),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_17),
.Y(n_229)
);


endmodule