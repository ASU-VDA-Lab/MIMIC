module fake_jpeg_27669_n_82 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_82);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_82;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_36),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_14),
.B1(n_24),
.B2(n_22),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_0),
.Y(n_47)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_12),
.B1(n_21),
.B2(n_20),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_38),
.A2(n_39),
.B1(n_31),
.B2(n_30),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_10),
.B1(n_19),
.B2(n_18),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_49),
.B1(n_4),
.B2(n_5),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_3),
.Y(n_58)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_1),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_31),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_50),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_34),
.A2(n_30),
.B1(n_8),
.B2(n_13),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_53),
.B(n_55),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_58),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_51),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_57),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_2),
.Y(n_57)
);

INVxp33_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

MAJx2_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_16),
.C(n_6),
.Y(n_61)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_4),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_52),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_73),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_67),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_68),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_52),
.C(n_71),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_66),
.Y(n_77)
);

AOI321xp33_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_76),
.A3(n_65),
.B1(n_72),
.B2(n_59),
.C(n_64),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_78),
.B(n_64),
.Y(n_79)
);

AO21x1_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_70),
.B(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_80),
.B(n_68),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_81),
.Y(n_82)
);


endmodule