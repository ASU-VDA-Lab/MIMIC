module fake_netlist_1_832_n_1279 (n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_292, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_291, n_170, n_294, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_283, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_293, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_290, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1279);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_292;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_291;
input n_170;
input n_294;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_283;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_293;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1279;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_315;
wire n_409;
wire n_295;
wire n_677;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_994;
wire n_930;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_303;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_948;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_335;
wire n_700;
wire n_534;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_405;
wire n_491;
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_200), .Y(n_295) );
INVxp67_ASAP7_75t_SL g296 ( .A(n_81), .Y(n_296) );
INVxp67_ASAP7_75t_L g297 ( .A(n_70), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_95), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_212), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_152), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_270), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_224), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_272), .Y(n_303) );
BUFx2_ASAP7_75t_L g304 ( .A(n_126), .Y(n_304) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_48), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_89), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_194), .Y(n_307) );
CKINVDCx20_ASAP7_75t_R g308 ( .A(n_244), .Y(n_308) );
INVx2_ASAP7_75t_SL g309 ( .A(n_149), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_273), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_210), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_239), .Y(n_312) );
OR2x2_ASAP7_75t_L g313 ( .A(n_197), .B(n_248), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_61), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_8), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_144), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_156), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_176), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_106), .Y(n_319) );
CKINVDCx20_ASAP7_75t_R g320 ( .A(n_142), .Y(n_320) );
INVxp33_ASAP7_75t_L g321 ( .A(n_76), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_255), .Y(n_322) );
INVx1_ASAP7_75t_SL g323 ( .A(n_181), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_31), .Y(n_324) );
CKINVDCx16_ASAP7_75t_R g325 ( .A(n_88), .Y(n_325) );
INVxp67_ASAP7_75t_L g326 ( .A(n_186), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_216), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_36), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_110), .Y(n_329) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_30), .Y(n_330) );
CKINVDCx20_ASAP7_75t_R g331 ( .A(n_16), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_21), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_96), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_242), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_283), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_141), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_73), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_154), .Y(n_338) );
BUFx6f_ASAP7_75t_L g339 ( .A(n_102), .Y(n_339) );
BUFx3_ASAP7_75t_L g340 ( .A(n_231), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_187), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_145), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_230), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_109), .Y(n_344) );
CKINVDCx16_ASAP7_75t_R g345 ( .A(n_207), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_53), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_278), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_123), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_228), .Y(n_349) );
INVxp67_ASAP7_75t_SL g350 ( .A(n_49), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_125), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_293), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_163), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_90), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_83), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_227), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_105), .Y(n_357) );
INVxp67_ASAP7_75t_L g358 ( .A(n_147), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_286), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_183), .Y(n_360) );
CKINVDCx20_ASAP7_75t_R g361 ( .A(n_213), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_249), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_172), .Y(n_363) );
CKINVDCx20_ASAP7_75t_R g364 ( .A(n_206), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_94), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_135), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_40), .Y(n_367) );
INVxp67_ASAP7_75t_SL g368 ( .A(n_294), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_82), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_215), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_288), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_18), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_205), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g374 ( .A(n_168), .Y(n_374) );
INVxp67_ASAP7_75t_SL g375 ( .A(n_75), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_177), .Y(n_376) );
INVxp33_ASAP7_75t_L g377 ( .A(n_0), .Y(n_377) );
CKINVDCx20_ASAP7_75t_R g378 ( .A(n_36), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_160), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_150), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_219), .Y(n_381) );
INVxp67_ASAP7_75t_SL g382 ( .A(n_280), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_37), .Y(n_383) );
CKINVDCx14_ASAP7_75t_R g384 ( .A(n_174), .Y(n_384) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_218), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_41), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_190), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_192), .Y(n_388) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_31), .Y(n_389) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_281), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_151), .Y(n_391) );
INVxp67_ASAP7_75t_SL g392 ( .A(n_50), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_71), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_41), .B(n_25), .Y(n_394) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_35), .Y(n_395) );
INVxp33_ASAP7_75t_L g396 ( .A(n_51), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_217), .Y(n_397) );
CKINVDCx5p33_ASAP7_75t_R g398 ( .A(n_185), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_26), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_112), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_241), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_100), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_166), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_139), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_265), .Y(n_405) );
INVxp67_ASAP7_75t_SL g406 ( .A(n_274), .Y(n_406) );
INVxp67_ASAP7_75t_SL g407 ( .A(n_140), .Y(n_407) );
CKINVDCx16_ASAP7_75t_R g408 ( .A(n_108), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_148), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_277), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_93), .Y(n_411) );
BUFx3_ASAP7_75t_L g412 ( .A(n_146), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_17), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_57), .Y(n_414) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_153), .Y(n_415) );
INVxp67_ASAP7_75t_L g416 ( .A(n_263), .Y(n_416) );
CKINVDCx16_ASAP7_75t_R g417 ( .A(n_53), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_268), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_47), .Y(n_419) );
INVxp67_ASAP7_75t_L g420 ( .A(n_276), .Y(n_420) );
INVxp33_ASAP7_75t_SL g421 ( .A(n_23), .Y(n_421) );
INVxp67_ASAP7_75t_SL g422 ( .A(n_107), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_236), .B(n_138), .Y(n_423) );
INVxp67_ASAP7_75t_SL g424 ( .A(n_232), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_19), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_59), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_4), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_119), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_291), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_223), .Y(n_430) );
CKINVDCx16_ASAP7_75t_R g431 ( .A(n_114), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_98), .Y(n_432) );
INVxp33_ASAP7_75t_L g433 ( .A(n_50), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_143), .Y(n_434) );
INVxp33_ASAP7_75t_SL g435 ( .A(n_24), .Y(n_435) );
CKINVDCx5p33_ASAP7_75t_R g436 ( .A(n_246), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_11), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_2), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_178), .Y(n_439) );
INVxp33_ASAP7_75t_L g440 ( .A(n_180), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_49), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_250), .Y(n_442) );
INVxp67_ASAP7_75t_SL g443 ( .A(n_67), .Y(n_443) );
INVxp33_ASAP7_75t_L g444 ( .A(n_68), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_162), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_377), .B(n_0), .Y(n_446) );
AND2x2_ASAP7_75t_SL g447 ( .A(n_304), .B(n_292), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_334), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_334), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_305), .B(n_1), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_348), .Y(n_451) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_339), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_372), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_372), .Y(n_454) );
BUFx2_ASAP7_75t_L g455 ( .A(n_395), .Y(n_455) );
AND2x2_ASAP7_75t_SL g456 ( .A(n_313), .B(n_72), .Y(n_456) );
CKINVDCx16_ASAP7_75t_R g457 ( .A(n_325), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_330), .Y(n_458) );
AND2x4_ASAP7_75t_L g459 ( .A(n_413), .B(n_1), .Y(n_459) );
AND2x4_ASAP7_75t_L g460 ( .A(n_413), .B(n_3), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_348), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_366), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_425), .Y(n_463) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_339), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_417), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_366), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_421), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_467) );
NOR2xp67_ASAP7_75t_L g468 ( .A(n_371), .B(n_5), .Y(n_468) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_339), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_425), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_298), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_299), .Y(n_472) );
CKINVDCx5p33_ASAP7_75t_R g473 ( .A(n_345), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_300), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_385), .B(n_6), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_301), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_302), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_428), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_303), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_428), .Y(n_480) );
BUFx6f_ASAP7_75t_L g481 ( .A(n_339), .Y(n_481) );
INVx4_ASAP7_75t_L g482 ( .A(n_459), .Y(n_482) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_481), .Y(n_483) );
NAND3x1_ASAP7_75t_L g484 ( .A(n_467), .B(n_394), .C(n_315), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_455), .B(n_377), .Y(n_485) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_457), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_452), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_471), .B(n_321), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_459), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_457), .B(n_321), .Y(n_490) );
INVx3_ASAP7_75t_L g491 ( .A(n_459), .Y(n_491) );
NAND2x1p5_ASAP7_75t_L g492 ( .A(n_456), .B(n_306), .Y(n_492) );
AND2x2_ASAP7_75t_SL g493 ( .A(n_456), .B(n_447), .Y(n_493) );
AND2x2_ASAP7_75t_SL g494 ( .A(n_456), .B(n_408), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_455), .B(n_396), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_460), .Y(n_496) );
BUFx10_ASAP7_75t_L g497 ( .A(n_473), .Y(n_497) );
INVx4_ASAP7_75t_L g498 ( .A(n_460), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_446), .B(n_396), .Y(n_499) );
INVx3_ASAP7_75t_L g500 ( .A(n_460), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_460), .Y(n_501) );
INVx4_ASAP7_75t_L g502 ( .A(n_447), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_448), .Y(n_503) );
INVx4_ASAP7_75t_L g504 ( .A(n_447), .Y(n_504) );
AND2x4_ASAP7_75t_L g505 ( .A(n_471), .B(n_405), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_452), .Y(n_506) );
AND2x6_ASAP7_75t_L g507 ( .A(n_446), .B(n_340), .Y(n_507) );
INVxp33_ASAP7_75t_L g508 ( .A(n_450), .Y(n_508) );
AND2x6_ASAP7_75t_L g509 ( .A(n_472), .B(n_340), .Y(n_509) );
INVx3_ASAP7_75t_L g510 ( .A(n_448), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_472), .B(n_433), .Y(n_511) );
BUFx6f_ASAP7_75t_L g512 ( .A(n_481), .Y(n_512) );
INVx5_ASAP7_75t_L g513 ( .A(n_481), .Y(n_513) );
AND2x6_ASAP7_75t_L g514 ( .A(n_474), .B(n_412), .Y(n_514) );
AND2x4_ASAP7_75t_L g515 ( .A(n_474), .B(n_415), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_449), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_476), .B(n_440), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_465), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_476), .B(n_440), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_449), .Y(n_520) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_481), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_477), .B(n_433), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_477), .B(n_309), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_479), .B(n_297), .Y(n_524) );
BUFx6f_ASAP7_75t_L g525 ( .A(n_481), .Y(n_525) );
INVx3_ASAP7_75t_L g526 ( .A(n_451), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_452), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_510), .Y(n_528) );
OR2x2_ASAP7_75t_SL g529 ( .A(n_518), .B(n_431), .Y(n_529) );
INVx5_ASAP7_75t_L g530 ( .A(n_509), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_505), .B(n_479), .Y(n_531) );
INVx4_ASAP7_75t_L g532 ( .A(n_507), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_503), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_503), .Y(n_534) );
BUFx3_ASAP7_75t_L g535 ( .A(n_497), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_510), .Y(n_536) );
INVx4_ASAP7_75t_L g537 ( .A(n_507), .Y(n_537) );
INVx2_ASAP7_75t_SL g538 ( .A(n_511), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_516), .Y(n_539) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_505), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_505), .B(n_475), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_516), .Y(n_542) );
INVx3_ASAP7_75t_L g543 ( .A(n_482), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_520), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_485), .B(n_399), .Y(n_545) );
OR2x6_ASAP7_75t_L g546 ( .A(n_502), .B(n_468), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_508), .B(n_468), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_520), .Y(n_548) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_509), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_505), .B(n_451), .Y(n_550) );
NAND2x1p5_ASAP7_75t_L g551 ( .A(n_515), .B(n_467), .Y(n_551) );
INVx2_ASAP7_75t_SL g552 ( .A(n_511), .Y(n_552) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_495), .Y(n_553) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_509), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_493), .A2(n_435), .B1(n_421), .B2(n_308), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_515), .B(n_488), .Y(n_556) );
AOI21xp33_ASAP7_75t_L g557 ( .A1(n_494), .A2(n_310), .B(n_307), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_515), .B(n_461), .Y(n_558) );
INVx2_ASAP7_75t_SL g559 ( .A(n_495), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_510), .Y(n_560) );
AND2x6_ASAP7_75t_SL g561 ( .A(n_490), .B(n_314), .Y(n_561) );
O2A1O1Ixp33_ASAP7_75t_L g562 ( .A1(n_489), .A2(n_454), .B(n_463), .C(n_453), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_515), .B(n_295), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_499), .B(n_444), .Y(n_564) );
INVx2_ASAP7_75t_SL g565 ( .A(n_499), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_510), .Y(n_566) );
INVx2_ASAP7_75t_SL g567 ( .A(n_522), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_517), .B(n_519), .Y(n_568) );
BUFx3_ASAP7_75t_L g569 ( .A(n_497), .Y(n_569) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_482), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_482), .B(n_498), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_526), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_482), .B(n_295), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_498), .B(n_461), .Y(n_574) );
AND2x4_ASAP7_75t_L g575 ( .A(n_498), .B(n_308), .Y(n_575) );
OAI22xp5_ASAP7_75t_SL g576 ( .A1(n_493), .A2(n_331), .B1(n_378), .B2(n_435), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_498), .B(n_326), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_496), .B(n_462), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_496), .B(n_462), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_526), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_501), .Y(n_581) );
INVx2_ASAP7_75t_SL g582 ( .A(n_497), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g583 ( .A1(n_501), .A2(n_478), .B(n_466), .Y(n_583) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_494), .B(n_311), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_491), .B(n_466), .Y(n_585) );
INVx2_ASAP7_75t_SL g586 ( .A(n_497), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_491), .B(n_478), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_491), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_500), .B(n_480), .Y(n_589) );
INVx5_ASAP7_75t_L g590 ( .A(n_509), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_502), .A2(n_384), .B1(n_444), .B2(n_324), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_526), .Y(n_592) );
AND2x6_ASAP7_75t_SL g593 ( .A(n_486), .B(n_332), .Y(n_593) );
AND2x4_ASAP7_75t_L g594 ( .A(n_502), .B(n_320), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_492), .B(n_399), .Y(n_595) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_509), .Y(n_596) );
AND2x4_ASAP7_75t_L g597 ( .A(n_502), .B(n_320), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_504), .A2(n_384), .B1(n_346), .B2(n_383), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_526), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_500), .Y(n_600) );
AND2x4_ASAP7_75t_L g601 ( .A(n_504), .B(n_361), .Y(n_601) );
OR2x2_ASAP7_75t_SL g602 ( .A(n_484), .B(n_378), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_500), .B(n_480), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_507), .B(n_317), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_507), .B(n_317), .Y(n_605) );
CKINVDCx5p33_ASAP7_75t_R g606 ( .A(n_504), .Y(n_606) );
INVx2_ASAP7_75t_SL g607 ( .A(n_507), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_507), .B(n_327), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_524), .B(n_509), .Y(n_609) );
NAND2xp33_ASAP7_75t_SL g610 ( .A(n_492), .B(n_361), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_567), .B(n_414), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_574), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_568), .B(n_523), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_545), .B(n_419), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_568), .B(n_509), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_551), .A2(n_484), .B1(n_514), .B2(n_374), .Y(n_616) );
NOR2xp33_ASAP7_75t_SL g617 ( .A(n_532), .B(n_364), .Y(n_617) );
A2O1A1Ixp33_ASAP7_75t_L g618 ( .A1(n_562), .A2(n_427), .B(n_438), .C(n_426), .Y(n_618) );
A2O1A1Ixp33_ASAP7_75t_L g619 ( .A1(n_562), .A2(n_441), .B(n_392), .C(n_350), .Y(n_619) );
AND2x4_ASAP7_75t_L g620 ( .A(n_535), .B(n_443), .Y(n_620) );
OAI21xp33_ASAP7_75t_L g621 ( .A1(n_531), .A2(n_454), .B(n_453), .Y(n_621) );
O2A1O1Ixp5_ASAP7_75t_L g622 ( .A1(n_573), .A2(n_368), .B(n_375), .C(n_296), .Y(n_622) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_540), .Y(n_623) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_549), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_543), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_574), .Y(n_626) );
BUFx12f_ASAP7_75t_L g627 ( .A(n_593), .Y(n_627) );
A2O1A1Ixp33_ASAP7_75t_SL g628 ( .A1(n_547), .A2(n_577), .B(n_598), .C(n_591), .Y(n_628) );
BUFx2_ASAP7_75t_L g629 ( .A(n_575), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_543), .Y(n_630) );
CKINVDCx5p33_ASAP7_75t_R g631 ( .A(n_569), .Y(n_631) );
BUFx3_ASAP7_75t_L g632 ( .A(n_565), .Y(n_632) );
INVx3_ASAP7_75t_L g633 ( .A(n_532), .Y(n_633) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_549), .Y(n_634) );
AND2x4_ASAP7_75t_L g635 ( .A(n_582), .B(n_364), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_540), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_585), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_551), .A2(n_514), .B1(n_445), .B2(n_374), .Y(n_638) );
INVx3_ASAP7_75t_L g639 ( .A(n_537), .Y(n_639) );
AOI21xp5_ASAP7_75t_L g640 ( .A1(n_609), .A2(n_406), .B(n_382), .Y(n_640) );
NOR2xp67_ASAP7_75t_L g641 ( .A(n_537), .B(n_74), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_556), .A2(n_514), .B1(n_445), .B2(n_419), .Y(n_642) );
OAI22xp5_ASAP7_75t_SL g643 ( .A1(n_602), .A2(n_437), .B1(n_328), .B2(n_386), .Y(n_643) );
CKINVDCx5p33_ASAP7_75t_R g644 ( .A(n_561), .Y(n_644) );
INVx1_ASAP7_75t_SL g645 ( .A(n_575), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_585), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_556), .B(n_514), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_559), .B(n_437), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_553), .B(n_367), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_557), .A2(n_552), .B1(n_538), .B2(n_541), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_541), .A2(n_398), .B1(n_403), .B2(n_327), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_600), .Y(n_652) );
INVx2_ASAP7_75t_SL g653 ( .A(n_564), .Y(n_653) );
NAND3xp33_ASAP7_75t_SL g654 ( .A(n_555), .B(n_436), .C(n_403), .Y(n_654) );
INVx2_ASAP7_75t_SL g655 ( .A(n_531), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_587), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g657 ( .A1(n_609), .A2(n_422), .B(n_407), .Y(n_657) );
BUFx6f_ASAP7_75t_L g658 ( .A(n_549), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_606), .A2(n_436), .B1(n_424), .B2(n_358), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_594), .B(n_470), .Y(n_660) );
BUFx2_ASAP7_75t_L g661 ( .A(n_594), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_595), .B(n_416), .Y(n_662) );
BUFx3_ASAP7_75t_L g663 ( .A(n_529), .Y(n_663) );
A2O1A1Ixp33_ASAP7_75t_L g664 ( .A1(n_581), .A2(n_316), .B(n_318), .C(n_312), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g665 ( .A1(n_557), .A2(n_514), .B1(n_322), .B2(n_333), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_588), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_587), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_550), .B(n_514), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_610), .A2(n_514), .B1(n_335), .B2(n_336), .Y(n_669) );
INVx5_ASAP7_75t_L g670 ( .A(n_554), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_550), .B(n_420), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_530), .B(n_329), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_584), .A2(n_330), .B1(n_389), .B2(n_337), .Y(n_673) );
OAI21xp33_ASAP7_75t_SL g674 ( .A1(n_533), .A2(n_338), .B(n_319), .Y(n_674) );
AOI21xp5_ASAP7_75t_L g675 ( .A1(n_571), .A2(n_342), .B(n_341), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_534), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_589), .Y(n_677) );
INVx4_ASAP7_75t_L g678 ( .A(n_554), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_589), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_597), .A2(n_330), .B1(n_389), .B2(n_347), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g681 ( .A1(n_571), .A2(n_349), .B(n_343), .Y(n_681) );
BUFx2_ASAP7_75t_L g682 ( .A(n_601), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_601), .B(n_389), .Y(n_683) );
INVx1_ASAP7_75t_SL g684 ( .A(n_558), .Y(n_684) );
INVx3_ASAP7_75t_L g685 ( .A(n_554), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_539), .Y(n_686) );
O2A1O1Ixp33_ASAP7_75t_SL g687 ( .A1(n_603), .A2(n_351), .B(n_353), .C(n_352), .Y(n_687) );
INVx4_ASAP7_75t_L g688 ( .A(n_596), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_603), .A2(n_355), .B(n_354), .Y(n_689) );
INVx2_ASAP7_75t_SL g690 ( .A(n_558), .Y(n_690) );
NOR2xp67_ASAP7_75t_SL g691 ( .A(n_530), .B(n_344), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_576), .A2(n_359), .B1(n_360), .B2(n_357), .Y(n_692) );
INVx1_ASAP7_75t_SL g693 ( .A(n_563), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_570), .B(n_356), .Y(n_694) );
INVx2_ASAP7_75t_SL g695 ( .A(n_586), .Y(n_695) );
O2A1O1Ixp33_ASAP7_75t_L g696 ( .A1(n_578), .A2(n_362), .B(n_369), .C(n_365), .Y(n_696) );
O2A1O1Ixp33_ASAP7_75t_L g697 ( .A1(n_578), .A2(n_370), .B(n_380), .C(n_373), .Y(n_697) );
A2O1A1Ixp33_ASAP7_75t_SL g698 ( .A1(n_528), .A2(n_423), .B(n_458), .C(n_487), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_579), .Y(n_699) );
O2A1O1Ixp33_ASAP7_75t_L g700 ( .A1(n_579), .A2(n_381), .B(n_388), .C(n_387), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_570), .Y(n_701) );
INVx2_ASAP7_75t_L g702 ( .A(n_542), .Y(n_702) );
BUFx3_ASAP7_75t_L g703 ( .A(n_546), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_544), .A2(n_400), .B1(n_401), .B2(n_397), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_548), .Y(n_705) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_604), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_536), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_560), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_583), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_566), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_546), .B(n_363), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g712 ( .A1(n_604), .A2(n_404), .B(n_402), .Y(n_712) );
OAI22x1_ASAP7_75t_L g713 ( .A1(n_607), .A2(n_376), .B1(n_391), .B2(n_379), .Y(n_713) );
A2O1A1Ixp33_ASAP7_75t_SL g714 ( .A1(n_572), .A2(n_580), .B(n_599), .C(n_592), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_608), .A2(n_410), .B1(n_411), .B2(n_409), .Y(n_715) );
AOI222xp33_ASAP7_75t_L g716 ( .A1(n_605), .A2(n_439), .B1(n_432), .B2(n_418), .C1(n_429), .C2(n_430), .Y(n_716) );
AND2x4_ASAP7_75t_L g717 ( .A(n_530), .B(n_412), .Y(n_717) );
INVx3_ASAP7_75t_L g718 ( .A(n_596), .Y(n_718) );
HAxp5_ASAP7_75t_L g719 ( .A(n_605), .B(n_6), .CON(n_719), .SN(n_719) );
CKINVDCx11_ASAP7_75t_R g720 ( .A(n_590), .Y(n_720) );
OR2x6_ASAP7_75t_L g721 ( .A(n_590), .B(n_434), .Y(n_721) );
AND2x4_ASAP7_75t_L g722 ( .A(n_590), .B(n_7), .Y(n_722) );
AOI21xp5_ASAP7_75t_L g723 ( .A1(n_590), .A2(n_442), .B(n_434), .Y(n_723) );
INVxp67_ASAP7_75t_L g724 ( .A(n_567), .Y(n_724) );
AND2x4_ASAP7_75t_SL g725 ( .A(n_575), .B(n_442), .Y(n_725) );
INVx3_ASAP7_75t_L g726 ( .A(n_543), .Y(n_726) );
BUFx2_ASAP7_75t_L g727 ( .A(n_575), .Y(n_727) );
CKINVDCx8_ASAP7_75t_R g728 ( .A(n_593), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_568), .B(n_393), .Y(n_729) );
AOI21xp5_ASAP7_75t_SL g730 ( .A1(n_532), .A2(n_390), .B(n_487), .Y(n_730) );
O2A1O1Ixp5_ASAP7_75t_SL g731 ( .A1(n_557), .A2(n_458), .B(n_464), .C(n_452), .Y(n_731) );
OR2x6_ASAP7_75t_L g732 ( .A(n_594), .B(n_390), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_556), .A2(n_323), .B1(n_458), .B2(n_390), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_574), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_568), .B(n_458), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_574), .Y(n_736) );
INVx3_ASAP7_75t_L g737 ( .A(n_678), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_699), .B(n_7), .Y(n_738) );
BUFx2_ASAP7_75t_L g739 ( .A(n_732), .Y(n_739) );
OAI21x1_ASAP7_75t_L g740 ( .A1(n_731), .A2(n_527), .B(n_506), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_655), .A2(n_390), .B1(n_464), .B2(n_469), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_653), .A2(n_464), .B1(n_469), .B2(n_481), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_612), .B(n_8), .Y(n_743) );
OR2x2_ASAP7_75t_L g744 ( .A(n_614), .B(n_9), .Y(n_744) );
AND2x4_ASAP7_75t_SL g745 ( .A(n_732), .B(n_464), .Y(n_745) );
BUFx8_ASAP7_75t_L g746 ( .A(n_627), .Y(n_746) );
A2O1A1Ixp33_ASAP7_75t_L g747 ( .A1(n_709), .A2(n_469), .B(n_464), .C(n_513), .Y(n_747) );
NAND2x1p5_ASAP7_75t_L g748 ( .A(n_670), .B(n_513), .Y(n_748) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_638), .A2(n_469), .B1(n_513), .B2(n_483), .Y(n_749) );
BUFx2_ASAP7_75t_L g750 ( .A(n_732), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_735), .Y(n_751) );
OAI21x1_ASAP7_75t_L g752 ( .A1(n_641), .A2(n_78), .B(n_77), .Y(n_752) );
NAND2x1p5_ASAP7_75t_L g753 ( .A(n_670), .B(n_513), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_638), .A2(n_469), .B1(n_513), .B2(n_483), .Y(n_754) );
BUFx6f_ASAP7_75t_L g755 ( .A(n_624), .Y(n_755) );
INVx6_ASAP7_75t_L g756 ( .A(n_670), .Y(n_756) );
AND2x4_ASAP7_75t_L g757 ( .A(n_703), .B(n_9), .Y(n_757) );
OAI21x1_ASAP7_75t_L g758 ( .A1(n_723), .A2(n_730), .B(n_712), .Y(n_758) );
INVx2_ASAP7_75t_L g759 ( .A(n_676), .Y(n_759) );
OR2x6_ASAP7_75t_L g760 ( .A(n_635), .B(n_10), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_616), .A2(n_513), .B1(n_483), .B2(n_525), .Y(n_761) );
OAI21x1_ASAP7_75t_L g762 ( .A1(n_675), .A2(n_80), .B(n_79), .Y(n_762) );
OAI21xp5_ASAP7_75t_L g763 ( .A1(n_615), .A2(n_483), .B(n_10), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_643), .A2(n_483), .B1(n_521), .B2(n_512), .Y(n_764) );
NOR2xp67_ASAP7_75t_SL g765 ( .A(n_728), .B(n_11), .Y(n_765) );
INVx2_ASAP7_75t_SL g766 ( .A(n_631), .Y(n_766) );
AND2x2_ASAP7_75t_L g767 ( .A(n_611), .B(n_12), .Y(n_767) );
OR2x6_ASAP7_75t_L g768 ( .A(n_635), .B(n_12), .Y(n_768) );
INVx2_ASAP7_75t_L g769 ( .A(n_686), .Y(n_769) );
AOI22x1_ASAP7_75t_L g770 ( .A1(n_681), .A2(n_525), .B1(n_521), .B2(n_512), .Y(n_770) );
AND2x2_ASAP7_75t_L g771 ( .A(n_724), .B(n_13), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_702), .Y(n_772) );
OAI21x1_ASAP7_75t_L g773 ( .A1(n_689), .A2(n_85), .B(n_84), .Y(n_773) );
AND2x4_ASAP7_75t_L g774 ( .A(n_695), .B(n_13), .Y(n_774) );
CKINVDCx8_ASAP7_75t_R g775 ( .A(n_644), .Y(n_775) );
NAND2x1p5_ASAP7_75t_L g776 ( .A(n_678), .B(n_14), .Y(n_776) );
OAI21xp5_ASAP7_75t_L g777 ( .A1(n_674), .A2(n_14), .B(n_15), .Y(n_777) );
OAI21x1_ASAP7_75t_L g778 ( .A1(n_705), .A2(n_87), .B(n_86), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_626), .B(n_15), .Y(n_779) );
OAI21x1_ASAP7_75t_SL g780 ( .A1(n_669), .A2(n_16), .B(n_17), .Y(n_780) );
HB1xp67_ASAP7_75t_L g781 ( .A(n_734), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_645), .B(n_18), .Y(n_782) );
INVx2_ASAP7_75t_L g783 ( .A(n_701), .Y(n_783) );
OAI21x1_ASAP7_75t_L g784 ( .A1(n_666), .A2(n_92), .B(n_91), .Y(n_784) );
CKINVDCx16_ASAP7_75t_R g785 ( .A(n_617), .Y(n_785) );
OAI21xp5_ASAP7_75t_L g786 ( .A1(n_674), .A2(n_19), .B(n_20), .Y(n_786) );
INVx6_ASAP7_75t_L g787 ( .A(n_688), .Y(n_787) );
A2O1A1Ixp33_ASAP7_75t_L g788 ( .A1(n_637), .A2(n_525), .B(n_521), .C(n_512), .Y(n_788) );
AO21x2_ASAP7_75t_L g789 ( .A1(n_698), .A2(n_521), .B(n_512), .Y(n_789) );
OAI21x1_ASAP7_75t_L g790 ( .A1(n_707), .A2(n_99), .B(n_97), .Y(n_790) );
INVx2_ASAP7_75t_L g791 ( .A(n_652), .Y(n_791) );
OAI22xp33_ASAP7_75t_L g792 ( .A1(n_617), .A2(n_20), .B1(n_21), .B2(n_22), .Y(n_792) );
NAND2x1p5_ASAP7_75t_L g793 ( .A(n_688), .B(n_22), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_683), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_645), .B(n_24), .Y(n_795) );
INVx4_ASAP7_75t_L g796 ( .A(n_720), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_660), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_623), .Y(n_798) );
O2A1O1Ixp33_ASAP7_75t_SL g799 ( .A1(n_628), .A2(n_167), .B(n_290), .C(n_289), .Y(n_799) );
AND2x2_ASAP7_75t_L g800 ( .A(n_629), .B(n_25), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_636), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_625), .Y(n_802) );
OAI21x1_ASAP7_75t_L g803 ( .A1(n_708), .A2(n_103), .B(n_101), .Y(n_803) );
OAI21x1_ASAP7_75t_L g804 ( .A1(n_672), .A2(n_639), .B(n_633), .Y(n_804) );
OAI21x1_ASAP7_75t_L g805 ( .A1(n_633), .A2(n_111), .B(n_104), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_690), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_736), .Y(n_807) );
OAI21x1_ASAP7_75t_L g808 ( .A1(n_639), .A2(n_115), .B(n_113), .Y(n_808) );
INVx4_ASAP7_75t_L g809 ( .A(n_722), .Y(n_809) );
CKINVDCx11_ASAP7_75t_R g810 ( .A(n_663), .Y(n_810) );
AO32x2_ASAP7_75t_L g811 ( .A1(n_680), .A2(n_26), .A3(n_27), .B1(n_28), .B2(n_29), .Y(n_811) );
OAI21x1_ASAP7_75t_L g812 ( .A1(n_710), .A2(n_117), .B(n_116), .Y(n_812) );
AND2x4_ASAP7_75t_L g813 ( .A(n_684), .B(n_27), .Y(n_813) );
INVx2_ASAP7_75t_L g814 ( .A(n_630), .Y(n_814) );
BUFx3_ASAP7_75t_L g815 ( .A(n_632), .Y(n_815) );
INVx3_ASAP7_75t_L g816 ( .A(n_624), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_646), .B(n_28), .Y(n_817) );
OA21x2_ASAP7_75t_L g818 ( .A1(n_621), .A2(n_521), .B(n_512), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_656), .B(n_29), .Y(n_819) );
BUFx3_ASAP7_75t_L g820 ( .A(n_620), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g821 ( .A1(n_616), .A2(n_525), .B1(n_521), .B2(n_512), .Y(n_821) );
NOR2xp33_ASAP7_75t_L g822 ( .A(n_661), .B(n_30), .Y(n_822) );
O2A1O1Ixp33_ASAP7_75t_SL g823 ( .A1(n_714), .A2(n_179), .B(n_287), .C(n_285), .Y(n_823) );
OAI21x1_ASAP7_75t_L g824 ( .A1(n_685), .A2(n_173), .B(n_284), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_643), .A2(n_525), .B1(n_33), .B2(n_34), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_667), .B(n_32), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_677), .Y(n_827) );
OAI21x1_ASAP7_75t_L g828 ( .A1(n_685), .A2(n_171), .B(n_282), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_679), .Y(n_829) );
OA21x2_ASAP7_75t_L g830 ( .A1(n_621), .A2(n_525), .B(n_170), .Y(n_830) );
BUFx3_ASAP7_75t_L g831 ( .A(n_620), .Y(n_831) );
O2A1O1Ixp33_ASAP7_75t_L g832 ( .A1(n_618), .A2(n_32), .B(n_33), .C(n_34), .Y(n_832) );
INVx2_ASAP7_75t_L g833 ( .A(n_726), .Y(n_833) );
OAI21x1_ASAP7_75t_SL g834 ( .A1(n_669), .A2(n_35), .B(n_37), .Y(n_834) );
OAI222xp33_ASAP7_75t_L g835 ( .A1(n_692), .A2(n_38), .B1(n_39), .B2(n_40), .C1(n_42), .C2(n_43), .Y(n_835) );
INVx2_ASAP7_75t_L g836 ( .A(n_726), .Y(n_836) );
OAI21xp5_ASAP7_75t_L g837 ( .A1(n_647), .A2(n_38), .B(n_39), .Y(n_837) );
OAI21x1_ASAP7_75t_L g838 ( .A1(n_718), .A2(n_182), .B(n_275), .Y(n_838) );
OA21x2_ASAP7_75t_L g839 ( .A1(n_664), .A2(n_665), .B(n_657), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_727), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_613), .Y(n_841) );
INVx3_ASAP7_75t_L g842 ( .A(n_624), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_682), .Y(n_843) );
AND2x2_ASAP7_75t_L g844 ( .A(n_692), .B(n_42), .Y(n_844) );
INVx2_ASAP7_75t_L g845 ( .A(n_722), .Y(n_845) );
OAI21x1_ASAP7_75t_L g846 ( .A1(n_733), .A2(n_184), .B(n_271), .Y(n_846) );
NOR2xp33_ASAP7_75t_L g847 ( .A(n_654), .B(n_43), .Y(n_847) );
NAND3xp33_ASAP7_75t_L g848 ( .A(n_716), .B(n_44), .C(n_45), .Y(n_848) );
OAI22xp5_ASAP7_75t_L g849 ( .A1(n_642), .A2(n_44), .B1(n_45), .B2(n_46), .Y(n_849) );
BUFx2_ASAP7_75t_SL g850 ( .A(n_717), .Y(n_850) );
OAI21x1_ASAP7_75t_L g851 ( .A1(n_668), .A2(n_188), .B(n_269), .Y(n_851) );
INVx2_ASAP7_75t_SL g852 ( .A(n_725), .Y(n_852) );
INVx3_ASAP7_75t_SL g853 ( .A(n_721), .Y(n_853) );
AND2x2_ASAP7_75t_L g854 ( .A(n_719), .B(n_46), .Y(n_854) );
OAI21xp5_ASAP7_75t_L g855 ( .A1(n_619), .A2(n_48), .B(n_51), .Y(n_855) );
OAI21x1_ASAP7_75t_L g856 ( .A1(n_622), .A2(n_640), .B(n_696), .Y(n_856) );
OAI21x1_ASAP7_75t_L g857 ( .A1(n_697), .A2(n_191), .B(n_267), .Y(n_857) );
OAI21xp5_ASAP7_75t_L g858 ( .A1(n_665), .A2(n_52), .B(n_54), .Y(n_858) );
INVxp33_ASAP7_75t_L g859 ( .A(n_642), .Y(n_859) );
OAI21x1_ASAP7_75t_L g860 ( .A1(n_700), .A2(n_189), .B(n_266), .Y(n_860) );
INVx2_ASAP7_75t_L g861 ( .A(n_717), .Y(n_861) );
OAI21x1_ASAP7_75t_L g862 ( .A1(n_673), .A2(n_175), .B(n_264), .Y(n_862) );
OAI21xp33_ASAP7_75t_SL g863 ( .A1(n_704), .A2(n_52), .B(n_54), .Y(n_863) );
INVx2_ASAP7_75t_L g864 ( .A(n_721), .Y(n_864) );
NAND3xp33_ASAP7_75t_L g865 ( .A(n_650), .B(n_55), .C(n_56), .Y(n_865) );
OAI21x1_ASAP7_75t_L g866 ( .A1(n_715), .A2(n_193), .B(n_262), .Y(n_866) );
OR2x6_ASAP7_75t_L g867 ( .A(n_721), .B(n_55), .Y(n_867) );
INVx4_ASAP7_75t_SL g868 ( .A(n_634), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_671), .Y(n_869) );
NAND2x1p5_ASAP7_75t_L g870 ( .A(n_634), .B(n_658), .Y(n_870) );
AO21x2_ASAP7_75t_L g871 ( .A1(n_687), .A2(n_169), .B(n_261), .Y(n_871) );
AND2x4_ASAP7_75t_L g872 ( .A(n_693), .B(n_56), .Y(n_872) );
OAI21xp5_ASAP7_75t_L g873 ( .A1(n_706), .A2(n_57), .B(n_58), .Y(n_873) );
INVx5_ASAP7_75t_L g874 ( .A(n_634), .Y(n_874) );
BUFx3_ASAP7_75t_L g875 ( .A(n_658), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_704), .Y(n_876) );
AOI21x1_ASAP7_75t_L g877 ( .A1(n_691), .A2(n_195), .B(n_260), .Y(n_877) );
AOI21xp5_ASAP7_75t_L g878 ( .A1(n_788), .A2(n_729), .B(n_658), .Y(n_878) );
OR2x2_ASAP7_75t_L g879 ( .A(n_841), .B(n_651), .Y(n_879) );
AND2x2_ASAP7_75t_L g880 ( .A(n_844), .B(n_662), .Y(n_880) );
OAI211xp5_ASAP7_75t_L g881 ( .A1(n_825), .A2(n_649), .B(n_648), .C(n_711), .Y(n_881) );
NOR4xp25_ASAP7_75t_L g882 ( .A(n_835), .B(n_659), .C(n_694), .D(n_60), .Y(n_882) );
A2O1A1Ixp33_ASAP7_75t_L g883 ( .A1(n_777), .A2(n_713), .B(n_59), .C(n_61), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_760), .A2(n_58), .B1(n_62), .B2(n_63), .Y(n_884) );
INVx5_ASAP7_75t_SL g885 ( .A(n_867), .Y(n_885) );
A2O1A1Ixp33_ASAP7_75t_L g886 ( .A1(n_777), .A2(n_62), .B(n_63), .C(n_64), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_760), .A2(n_64), .B1(n_65), .B2(n_66), .Y(n_887) );
AND2x2_ASAP7_75t_L g888 ( .A(n_760), .B(n_65), .Y(n_888) );
OAI22xp33_ASAP7_75t_L g889 ( .A1(n_768), .A2(n_66), .B1(n_67), .B2(n_68), .Y(n_889) );
AOI22xp33_ASAP7_75t_SL g890 ( .A1(n_785), .A2(n_69), .B1(n_118), .B2(n_120), .Y(n_890) );
AND2x2_ASAP7_75t_L g891 ( .A(n_768), .B(n_781), .Y(n_891) );
INVx8_ASAP7_75t_L g892 ( .A(n_867), .Y(n_892) );
OAI211xp5_ASAP7_75t_L g893 ( .A1(n_825), .A2(n_69), .B(n_121), .C(n_122), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_768), .A2(n_124), .B1(n_127), .B2(n_128), .Y(n_894) );
AND2x2_ASAP7_75t_L g895 ( .A(n_854), .B(n_129), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_876), .B(n_130), .Y(n_896) );
OAI21xp33_ASAP7_75t_L g897 ( .A1(n_848), .A2(n_131), .B(n_132), .Y(n_897) );
AOI221xp5_ASAP7_75t_L g898 ( .A1(n_869), .A2(n_133), .B1(n_134), .B2(n_136), .C(n_137), .Y(n_898) );
OA21x2_ASAP7_75t_L g899 ( .A1(n_747), .A2(n_155), .B(n_157), .Y(n_899) );
NAND2x1p5_ASAP7_75t_L g900 ( .A(n_809), .B(n_874), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_797), .B(n_158), .Y(n_901) );
OAI22xp5_ASAP7_75t_L g902 ( .A1(n_867), .A2(n_159), .B1(n_161), .B2(n_164), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_859), .A2(n_165), .B1(n_196), .B2(n_198), .Y(n_903) );
OAI211xp5_ASAP7_75t_L g904 ( .A1(n_863), .A2(n_199), .B(n_201), .C(n_202), .Y(n_904) );
OAI22xp5_ASAP7_75t_L g905 ( .A1(n_859), .A2(n_203), .B1(n_204), .B2(n_208), .Y(n_905) );
O2A1O1Ixp33_ASAP7_75t_L g906 ( .A1(n_849), .A2(n_209), .B(n_211), .C(n_214), .Y(n_906) );
BUFx4f_ASAP7_75t_SL g907 ( .A(n_746), .Y(n_907) );
BUFx8_ASAP7_75t_L g908 ( .A(n_766), .Y(n_908) );
AOI21xp5_ASAP7_75t_L g909 ( .A1(n_799), .A2(n_220), .B(n_221), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_798), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_801), .Y(n_911) );
AOI222xp33_ASAP7_75t_L g912 ( .A1(n_835), .A2(n_222), .B1(n_225), .B2(n_226), .C1(n_229), .C2(n_233), .Y(n_912) );
AOI21xp5_ASAP7_75t_L g913 ( .A1(n_789), .A2(n_234), .B(n_235), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_813), .A2(n_237), .B1(n_238), .B2(n_240), .Y(n_914) );
INVx2_ASAP7_75t_L g915 ( .A(n_807), .Y(n_915) );
OAI22xp33_ASAP7_75t_L g916 ( .A1(n_853), .A2(n_243), .B1(n_245), .B2(n_247), .Y(n_916) );
AOI21xp33_ASAP7_75t_L g917 ( .A1(n_761), .A2(n_279), .B(n_252), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_813), .A2(n_251), .B1(n_253), .B2(n_254), .Y(n_918) );
OR2x2_ASAP7_75t_L g919 ( .A(n_744), .B(n_256), .Y(n_919) );
INVx3_ASAP7_75t_L g920 ( .A(n_756), .Y(n_920) );
AOI22xp33_ASAP7_75t_SL g921 ( .A1(n_757), .A2(n_257), .B1(n_258), .B2(n_259), .Y(n_921) );
INVx2_ASAP7_75t_L g922 ( .A(n_827), .Y(n_922) );
INVx3_ASAP7_75t_L g923 ( .A(n_756), .Y(n_923) );
BUFx2_ASAP7_75t_L g924 ( .A(n_815), .Y(n_924) );
AOI221xp5_ASAP7_75t_L g925 ( .A1(n_849), .A2(n_843), .B1(n_840), .B2(n_822), .C(n_855), .Y(n_925) );
AOI221xp5_ASAP7_75t_L g926 ( .A1(n_822), .A2(n_855), .B1(n_829), .B2(n_832), .C(n_786), .Y(n_926) );
AO31x2_ASAP7_75t_L g927 ( .A1(n_747), .A2(n_821), .A3(n_754), .B(n_749), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_782), .A2(n_795), .B1(n_767), .B2(n_872), .Y(n_928) );
NAND4xp25_ASAP7_75t_L g929 ( .A(n_786), .B(n_847), .C(n_832), .D(n_873), .Y(n_929) );
NOR2x1_ASAP7_75t_SL g930 ( .A(n_809), .B(n_850), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_782), .A2(n_795), .B1(n_872), .B2(n_847), .Y(n_931) );
HB1xp67_ASAP7_75t_L g932 ( .A(n_757), .Y(n_932) );
INVx2_ASAP7_75t_L g933 ( .A(n_783), .Y(n_933) );
AOI221xp5_ASAP7_75t_SL g934 ( .A1(n_858), .A2(n_792), .B1(n_873), .B2(n_837), .C(n_754), .Y(n_934) );
OAI22xp33_ASAP7_75t_L g935 ( .A1(n_853), .A2(n_858), .B1(n_792), .B2(n_738), .Y(n_935) );
AND2x2_ASAP7_75t_L g936 ( .A(n_774), .B(n_800), .Y(n_936) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_749), .A2(n_738), .B1(n_779), .B2(n_743), .Y(n_937) );
AND2x2_ASAP7_75t_L g938 ( .A(n_774), .B(n_759), .Y(n_938) );
OAI22xp33_ASAP7_75t_L g939 ( .A1(n_796), .A2(n_779), .B1(n_743), .B2(n_817), .Y(n_939) );
OA21x2_ASAP7_75t_L g940 ( .A1(n_740), .A2(n_763), .B(n_778), .Y(n_940) );
AOI221xp5_ASAP7_75t_L g941 ( .A1(n_751), .A2(n_831), .B1(n_820), .B2(n_806), .C(n_771), .Y(n_941) );
AOI21xp5_ASAP7_75t_L g942 ( .A1(n_789), .A2(n_823), .B(n_770), .Y(n_942) );
AOI221xp5_ASAP7_75t_L g943 ( .A1(n_852), .A2(n_794), .B1(n_837), .B2(n_865), .C(n_819), .Y(n_943) );
AOI21xp33_ASAP7_75t_L g944 ( .A1(n_839), .A2(n_817), .B(n_826), .Y(n_944) );
AOI21xp5_ASAP7_75t_L g945 ( .A1(n_823), .A2(n_818), .B(n_763), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_769), .B(n_772), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_819), .B(n_826), .Y(n_947) );
OR2x6_ASAP7_75t_L g948 ( .A(n_796), .B(n_739), .Y(n_948) );
AOI22xp33_ASAP7_75t_SL g949 ( .A1(n_776), .A2(n_793), .B1(n_834), .B2(n_780), .Y(n_949) );
OAI221xp5_ASAP7_75t_L g950 ( .A1(n_764), .A2(n_865), .B1(n_776), .B2(n_793), .C(n_765), .Y(n_950) );
AOI221xp5_ASAP7_75t_L g951 ( .A1(n_764), .A2(n_845), .B1(n_750), .B2(n_861), .C(n_864), .Y(n_951) );
AND2x2_ASAP7_75t_L g952 ( .A(n_791), .B(n_811), .Y(n_952) );
AND2x2_ASAP7_75t_L g953 ( .A(n_811), .B(n_802), .Y(n_953) );
A2O1A1Ixp33_ASAP7_75t_L g954 ( .A1(n_856), .A2(n_860), .B(n_857), .C(n_745), .Y(n_954) );
AOI211xp5_ASAP7_75t_L g955 ( .A1(n_866), .A2(n_846), .B(n_836), .C(n_833), .Y(n_955) );
OAI22xp5_ASAP7_75t_L g956 ( .A1(n_839), .A2(n_741), .B1(n_874), .B2(n_787), .Y(n_956) );
INVx2_ASAP7_75t_L g957 ( .A(n_814), .Y(n_957) );
AND2x2_ASAP7_75t_L g958 ( .A(n_811), .B(n_810), .Y(n_958) );
CKINVDCx11_ASAP7_75t_R g959 ( .A(n_775), .Y(n_959) );
A2O1A1Ixp33_ASAP7_75t_L g960 ( .A1(n_758), .A2(n_762), .B(n_773), .C(n_851), .Y(n_960) );
AOI211xp5_ASAP7_75t_L g961 ( .A1(n_805), .A2(n_808), .B(n_812), .C(n_752), .Y(n_961) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_737), .B(n_787), .Y(n_962) );
OAI221xp5_ASAP7_75t_L g963 ( .A1(n_742), .A2(n_741), .B1(n_737), .B2(n_787), .C(n_756), .Y(n_963) );
INVx3_ASAP7_75t_L g964 ( .A(n_874), .Y(n_964) );
INVx2_ASAP7_75t_L g965 ( .A(n_824), .Y(n_965) );
INVx1_ASAP7_75t_L g966 ( .A(n_828), .Y(n_966) );
BUFx6f_ASAP7_75t_L g967 ( .A(n_755), .Y(n_967) );
BUFx2_ASAP7_75t_L g968 ( .A(n_748), .Y(n_968) );
OAI22xp5_ASAP7_75t_L g969 ( .A1(n_874), .A2(n_742), .B1(n_870), .B2(n_830), .Y(n_969) );
INVx3_ASAP7_75t_L g970 ( .A(n_748), .Y(n_970) );
AND2x2_ASAP7_75t_L g971 ( .A(n_753), .B(n_875), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_838), .Y(n_972) );
HB1xp67_ASAP7_75t_L g973 ( .A(n_753), .Y(n_973) );
AND2x2_ASAP7_75t_L g974 ( .A(n_868), .B(n_842), .Y(n_974) );
AOI22xp5_ASAP7_75t_L g975 ( .A1(n_871), .A2(n_842), .B1(n_816), .B2(n_755), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_784), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_871), .A2(n_816), .B1(n_755), .B2(n_804), .Y(n_977) );
OAI211xp5_ASAP7_75t_SL g978 ( .A1(n_877), .A2(n_790), .B(n_803), .C(n_862), .Y(n_978) );
CKINVDCx11_ASAP7_75t_R g979 ( .A(n_868), .Y(n_979) );
AND2x2_ASAP7_75t_L g980 ( .A(n_868), .B(n_870), .Y(n_980) );
OA21x2_ASAP7_75t_L g981 ( .A1(n_818), .A2(n_747), .B(n_788), .Y(n_981) );
A2O1A1Ixp33_ASAP7_75t_L g982 ( .A1(n_830), .A2(n_777), .B(n_786), .C(n_493), .Y(n_982) );
AOI21xp5_ASAP7_75t_L g983 ( .A1(n_788), .A2(n_799), .B(n_698), .Y(n_983) );
AOI21xp5_ASAP7_75t_L g984 ( .A1(n_788), .A2(n_799), .B(n_698), .Y(n_984) );
AOI21xp5_ASAP7_75t_L g985 ( .A1(n_788), .A2(n_799), .B(n_698), .Y(n_985) );
OAI221xp5_ASAP7_75t_L g986 ( .A1(n_841), .A2(n_551), .B1(n_692), .B2(n_643), .C(n_616), .Y(n_986) );
OA21x2_ASAP7_75t_L g987 ( .A1(n_747), .A2(n_788), .B(n_740), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_760), .A2(n_493), .B1(n_504), .B2(n_502), .Y(n_988) );
AO21x1_ASAP7_75t_L g989 ( .A1(n_821), .A2(n_792), .B(n_761), .Y(n_989) );
AO21x2_ASAP7_75t_L g990 ( .A1(n_747), .A2(n_788), .B(n_763), .Y(n_990) );
OAI22xp5_ASAP7_75t_L g991 ( .A1(n_781), .A2(n_493), .B1(n_638), .B2(n_504), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_841), .Y(n_992) );
INVx1_ASAP7_75t_L g993 ( .A(n_841), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_760), .A2(n_493), .B1(n_504), .B2(n_502), .Y(n_994) );
AOI21xp5_ASAP7_75t_L g995 ( .A1(n_788), .A2(n_799), .B(n_698), .Y(n_995) );
OAI321xp33_ASAP7_75t_L g996 ( .A1(n_792), .A2(n_777), .A3(n_786), .B1(n_849), .B2(n_848), .C(n_858), .Y(n_996) );
CKINVDCx5p33_ASAP7_75t_R g997 ( .A(n_746), .Y(n_997) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_841), .B(n_876), .Y(n_998) );
AND2x2_ASAP7_75t_L g999 ( .A(n_933), .B(n_915), .Y(n_999) );
BUFx2_ASAP7_75t_L g1000 ( .A(n_892), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_922), .B(n_998), .Y(n_1001) );
CKINVDCx5p33_ASAP7_75t_R g1002 ( .A(n_907), .Y(n_1002) );
OR2x2_ASAP7_75t_L g1003 ( .A(n_885), .B(n_891), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_986), .A2(n_880), .B1(n_892), .B2(n_994), .Y(n_1004) );
INVx2_ASAP7_75t_L g1005 ( .A(n_981), .Y(n_1005) );
INVxp67_ASAP7_75t_L g1006 ( .A(n_924), .Y(n_1006) );
INVx2_ASAP7_75t_L g1007 ( .A(n_987), .Y(n_1007) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_992), .B(n_993), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_911), .B(n_879), .Y(n_1009) );
BUFx3_ASAP7_75t_L g1010 ( .A(n_900), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_957), .B(n_946), .Y(n_1011) );
INVx1_ASAP7_75t_L g1012 ( .A(n_952), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_953), .Y(n_1013) );
AND2x2_ASAP7_75t_L g1014 ( .A(n_938), .B(n_882), .Y(n_1014) );
AND2x2_ASAP7_75t_L g1015 ( .A(n_882), .B(n_947), .Y(n_1015) );
AND2x4_ASAP7_75t_L g1016 ( .A(n_980), .B(n_974), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_973), .B(n_885), .Y(n_1017) );
INVx1_ASAP7_75t_L g1018 ( .A(n_966), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g1019 ( .A(n_910), .B(n_936), .Y(n_1019) );
NOR2xp33_ASAP7_75t_L g1020 ( .A(n_932), .B(n_892), .Y(n_1020) );
AND2x2_ASAP7_75t_L g1021 ( .A(n_885), .B(n_968), .Y(n_1021) );
INVx1_ASAP7_75t_L g1022 ( .A(n_972), .Y(n_1022) );
OR2x2_ASAP7_75t_L g1023 ( .A(n_929), .B(n_928), .Y(n_1023) );
OAI21xp33_ASAP7_75t_L g1024 ( .A1(n_929), .A2(n_912), .B(n_886), .Y(n_1024) );
INVx2_ASAP7_75t_L g1025 ( .A(n_976), .Y(n_1025) );
NAND2xp5_ASAP7_75t_L g1026 ( .A(n_925), .B(n_941), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_970), .B(n_971), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_896), .Y(n_1028) );
BUFx2_ASAP7_75t_L g1029 ( .A(n_927), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_982), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_965), .Y(n_1031) );
OAI22xp5_ASAP7_75t_L g1032 ( .A1(n_988), .A2(n_991), .B1(n_931), .B2(n_887), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_970), .B(n_926), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g1034 ( .A(n_888), .B(n_881), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_895), .B(n_964), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_964), .B(n_912), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g1037 ( .A1(n_958), .A2(n_939), .B1(n_935), .B2(n_950), .Y(n_1037) );
HB1xp67_ASAP7_75t_L g1038 ( .A(n_900), .Y(n_1038) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_883), .B(n_934), .Y(n_1039) );
INVx2_ASAP7_75t_L g1040 ( .A(n_940), .Y(n_1040) );
NAND2xp5_ASAP7_75t_L g1041 ( .A(n_930), .B(n_919), .Y(n_1041) );
BUFx2_ASAP7_75t_L g1042 ( .A(n_927), .Y(n_1042) );
INVx2_ASAP7_75t_L g1043 ( .A(n_940), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_934), .B(n_884), .Y(n_1044) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_949), .B(n_943), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_899), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_944), .B(n_937), .Y(n_1047) );
INVx2_ASAP7_75t_L g1048 ( .A(n_990), .Y(n_1048) );
INVx2_ASAP7_75t_L g1049 ( .A(n_927), .Y(n_1049) );
AND2x4_ASAP7_75t_L g1050 ( .A(n_967), .B(n_975), .Y(n_1050) );
OR2x2_ASAP7_75t_L g1051 ( .A(n_962), .B(n_937), .Y(n_1051) );
BUFx6f_ASAP7_75t_L g1052 ( .A(n_967), .Y(n_1052) );
INVx1_ASAP7_75t_L g1053 ( .A(n_989), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_889), .B(n_920), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_956), .Y(n_1055) );
INVx2_ASAP7_75t_L g1056 ( .A(n_967), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_951), .B(n_901), .Y(n_1057) );
OAI31xp33_ASAP7_75t_L g1058 ( .A1(n_893), .A2(n_897), .A3(n_904), .B(n_902), .Y(n_1058) );
AO21x2_ASAP7_75t_L g1059 ( .A1(n_945), .A2(n_942), .B(n_985), .Y(n_1059) );
NOR2xp33_ASAP7_75t_L g1060 ( .A(n_908), .B(n_948), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_956), .Y(n_1061) );
OR2x2_ASAP7_75t_L g1062 ( .A(n_948), .B(n_923), .Y(n_1062) );
BUFx2_ASAP7_75t_L g1063 ( .A(n_948), .Y(n_1063) );
BUFx2_ASAP7_75t_L g1064 ( .A(n_969), .Y(n_1064) );
INVx4_ASAP7_75t_L g1065 ( .A(n_979), .Y(n_1065) );
INVx2_ASAP7_75t_SL g1066 ( .A(n_920), .Y(n_1066) );
INVx2_ASAP7_75t_L g1067 ( .A(n_963), .Y(n_1067) );
INVx2_ASAP7_75t_L g1068 ( .A(n_923), .Y(n_1068) );
HB1xp67_ASAP7_75t_L g1069 ( .A(n_997), .Y(n_1069) );
OAI21x1_ASAP7_75t_L g1070 ( .A1(n_977), .A2(n_984), .B(n_995), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_921), .B(n_894), .Y(n_1071) );
OR2x2_ASAP7_75t_L g1072 ( .A(n_878), .B(n_960), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_890), .B(n_914), .Y(n_1073) );
AND2x4_ASAP7_75t_L g1074 ( .A(n_954), .B(n_913), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_918), .B(n_903), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_996), .Y(n_1076) );
INVx5_ASAP7_75t_L g1077 ( .A(n_916), .Y(n_1077) );
INVx1_ASAP7_75t_L g1078 ( .A(n_955), .Y(n_1078) );
INVxp67_ASAP7_75t_SL g1079 ( .A(n_961), .Y(n_1079) );
INVx2_ASAP7_75t_L g1080 ( .A(n_905), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_906), .B(n_955), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_898), .B(n_917), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_961), .B(n_983), .Y(n_1083) );
INVx2_ASAP7_75t_L g1084 ( .A(n_978), .Y(n_1084) );
AND2x4_ASAP7_75t_L g1085 ( .A(n_909), .B(n_959), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_933), .B(n_777), .Y(n_1086) );
AND2x2_ASAP7_75t_L g1087 ( .A(n_933), .B(n_777), .Y(n_1087) );
BUFx3_ASAP7_75t_L g1088 ( .A(n_900), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_933), .B(n_777), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_952), .Y(n_1090) );
INVx2_ASAP7_75t_L g1091 ( .A(n_981), .Y(n_1091) );
OR2x2_ASAP7_75t_L g1092 ( .A(n_1023), .B(n_1012), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_1012), .B(n_1013), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1094 ( .A(n_1013), .B(n_1090), .Y(n_1094) );
NAND2xp5_ASAP7_75t_L g1095 ( .A(n_1001), .B(n_1015), .Y(n_1095) );
BUFx2_ASAP7_75t_L g1096 ( .A(n_1050), .Y(n_1096) );
INVxp33_ASAP7_75t_L g1097 ( .A(n_1060), .Y(n_1097) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1018), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g1099 ( .A(n_1001), .B(n_1015), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_1090), .B(n_1053), .Y(n_1100) );
NAND2xp5_ASAP7_75t_L g1101 ( .A(n_999), .B(n_1011), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_1053), .B(n_1047), .Y(n_1102) );
NAND3xp33_ASAP7_75t_L g1103 ( .A(n_1076), .B(n_1024), .C(n_1034), .Y(n_1103) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1018), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_1029), .B(n_1042), .Y(n_1105) );
AND2x4_ASAP7_75t_L g1106 ( .A(n_1022), .B(n_1050), .Y(n_1106) );
INVx1_ASAP7_75t_L g1107 ( .A(n_1022), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1042), .B(n_1014), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1025), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1025), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_1014), .B(n_1030), .Y(n_1111) );
NAND3xp33_ASAP7_75t_L g1112 ( .A(n_1076), .B(n_1024), .C(n_1023), .Y(n_1112) );
OR2x2_ASAP7_75t_L g1113 ( .A(n_1051), .B(n_1009), .Y(n_1113) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_1030), .B(n_999), .Y(n_1114) );
AOI221xp5_ASAP7_75t_L g1115 ( .A1(n_1026), .A2(n_1045), .B1(n_1033), .B2(n_1039), .C(n_1004), .Y(n_1115) );
BUFx3_ASAP7_75t_L g1116 ( .A(n_1010), .Y(n_1116) );
AOI322xp5_ASAP7_75t_L g1117 ( .A1(n_1036), .A2(n_1000), .A3(n_1045), .B1(n_1037), .B2(n_1008), .C1(n_1039), .C2(n_1019), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_1086), .B(n_1087), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_1086), .B(n_1087), .Y(n_1119) );
HB1xp67_ASAP7_75t_L g1120 ( .A(n_1038), .Y(n_1120) );
INVx3_ASAP7_75t_SL g1121 ( .A(n_1002), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1031), .Y(n_1122) );
OAI22xp33_ASAP7_75t_L g1123 ( .A1(n_1065), .A2(n_1041), .B1(n_1010), .B2(n_1088), .Y(n_1123) );
HB1xp67_ASAP7_75t_L g1124 ( .A(n_1010), .Y(n_1124) );
NAND2xp5_ASAP7_75t_L g1125 ( .A(n_1027), .B(n_1089), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1049), .B(n_1051), .Y(n_1126) );
INVx3_ASAP7_75t_L g1127 ( .A(n_1052), .Y(n_1127) );
NOR2xp33_ASAP7_75t_L g1128 ( .A(n_1069), .B(n_1006), .Y(n_1128) );
NAND4xp25_ASAP7_75t_L g1129 ( .A(n_1054), .B(n_1032), .C(n_1065), .D(n_1044), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_1083), .B(n_1048), .Y(n_1130) );
INVx2_ASAP7_75t_L g1131 ( .A(n_1040), .Y(n_1131) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1031), .Y(n_1132) );
AO21x2_ASAP7_75t_L g1133 ( .A1(n_1084), .A2(n_1046), .B(n_1059), .Y(n_1133) );
AOI33xp33_ASAP7_75t_L g1134 ( .A1(n_1017), .A2(n_1067), .A3(n_1021), .B1(n_1078), .B2(n_1057), .B3(n_1027), .Y(n_1134) );
OAI22xp5_ASAP7_75t_L g1135 ( .A1(n_1088), .A2(n_1077), .B1(n_1063), .B2(n_1064), .Y(n_1135) );
OR2x2_ASAP7_75t_L g1136 ( .A(n_1003), .B(n_1067), .Y(n_1136) );
OAI31xp33_ASAP7_75t_L g1137 ( .A1(n_1073), .A2(n_1071), .A3(n_1088), .B(n_1075), .Y(n_1137) );
AOI21xp5_ASAP7_75t_SL g1138 ( .A1(n_1085), .A2(n_1079), .B(n_1080), .Y(n_1138) );
INVxp67_ASAP7_75t_SL g1139 ( .A(n_1056), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g1140 ( .A1(n_1077), .A2(n_1080), .B1(n_1028), .B2(n_1085), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1055), .B(n_1061), .Y(n_1141) );
OAI221xp5_ASAP7_75t_L g1142 ( .A1(n_1058), .A2(n_1028), .B1(n_1020), .B2(n_1062), .C(n_1065), .Y(n_1142) );
HB1xp67_ASAP7_75t_L g1143 ( .A(n_1035), .Y(n_1143) );
BUFx2_ASAP7_75t_L g1144 ( .A(n_1050), .Y(n_1144) );
HB1xp67_ASAP7_75t_L g1145 ( .A(n_1035), .Y(n_1145) );
NOR2xp33_ASAP7_75t_L g1146 ( .A(n_1097), .B(n_1065), .Y(n_1146) );
OR2x2_ASAP7_75t_L g1147 ( .A(n_1095), .B(n_1055), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1118), .B(n_1078), .Y(n_1148) );
INVx2_ASAP7_75t_L g1149 ( .A(n_1131), .Y(n_1149) );
HB1xp67_ASAP7_75t_L g1150 ( .A(n_1120), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1098), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1152 ( .A(n_1118), .B(n_1005), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_1119), .B(n_1091), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1104), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1104), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_1119), .B(n_1091), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1099), .B(n_1016), .Y(n_1157) );
AND2x4_ASAP7_75t_L g1158 ( .A(n_1130), .B(n_1050), .Y(n_1158) );
HB1xp67_ASAP7_75t_L g1159 ( .A(n_1143), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1102), .B(n_1091), .Y(n_1160) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1107), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1108), .B(n_1007), .Y(n_1162) );
NOR2xp33_ASAP7_75t_L g1163 ( .A(n_1128), .B(n_1066), .Y(n_1163) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1107), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1108), .B(n_1007), .Y(n_1165) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1122), .Y(n_1166) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1122), .Y(n_1167) );
NAND2xp5_ASAP7_75t_SL g1168 ( .A(n_1123), .B(n_1085), .Y(n_1168) );
NAND2xp5_ASAP7_75t_L g1169 ( .A(n_1101), .B(n_1093), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1093), .B(n_1068), .Y(n_1170) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1132), .Y(n_1171) );
INVxp67_ASAP7_75t_L g1172 ( .A(n_1124), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1132), .Y(n_1173) );
INVx1_ASAP7_75t_SL g1174 ( .A(n_1121), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1111), .B(n_1043), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1111), .B(n_1084), .Y(n_1176) );
OAI221xp5_ASAP7_75t_SL g1177 ( .A1(n_1137), .A2(n_1081), .B1(n_1072), .B2(n_1080), .C(n_1084), .Y(n_1177) );
NAND2xp5_ASAP7_75t_L g1178 ( .A(n_1094), .B(n_1068), .Y(n_1178) );
INVxp33_ASAP7_75t_L g1179 ( .A(n_1129), .Y(n_1179) );
NAND3xp33_ASAP7_75t_L g1180 ( .A(n_1112), .B(n_1103), .C(n_1117), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1126), .B(n_1059), .Y(n_1181) );
INVx3_ASAP7_75t_L g1182 ( .A(n_1133), .Y(n_1182) );
INVx3_ASAP7_75t_L g1183 ( .A(n_1133), .Y(n_1183) );
BUFx2_ASAP7_75t_SL g1184 ( .A(n_1116), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1126), .B(n_1059), .Y(n_1185) );
NAND2xp5_ASAP7_75t_L g1186 ( .A(n_1114), .B(n_1066), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1100), .B(n_1072), .Y(n_1187) );
AND2x4_ASAP7_75t_L g1188 ( .A(n_1106), .B(n_1074), .Y(n_1188) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1109), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1110), .Y(n_1190) );
INVx4_ASAP7_75t_L g1191 ( .A(n_1116), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1100), .B(n_1070), .Y(n_1192) );
INVx2_ASAP7_75t_SL g1193 ( .A(n_1116), .Y(n_1193) );
INVx2_ASAP7_75t_L g1194 ( .A(n_1149), .Y(n_1194) );
AND2x4_ASAP7_75t_L g1195 ( .A(n_1188), .B(n_1106), .Y(n_1195) );
AND2x4_ASAP7_75t_L g1196 ( .A(n_1188), .B(n_1106), .Y(n_1196) );
OR2x2_ASAP7_75t_L g1197 ( .A(n_1159), .B(n_1092), .Y(n_1197) );
INVx2_ASAP7_75t_SL g1198 ( .A(n_1191), .Y(n_1198) );
INVx3_ASAP7_75t_L g1199 ( .A(n_1191), .Y(n_1199) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1151), .Y(n_1200) );
NAND2xp5_ASAP7_75t_L g1201 ( .A(n_1148), .B(n_1112), .Y(n_1201) );
NAND3xp33_ASAP7_75t_L g1202 ( .A(n_1180), .B(n_1103), .C(n_1129), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1152), .B(n_1106), .Y(n_1203) );
NAND3xp33_ASAP7_75t_L g1204 ( .A(n_1180), .B(n_1117), .C(n_1115), .Y(n_1204) );
OR2x2_ASAP7_75t_L g1205 ( .A(n_1169), .B(n_1113), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1148), .B(n_1145), .Y(n_1206) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1154), .Y(n_1207) );
HB1xp67_ASAP7_75t_L g1208 ( .A(n_1150), .Y(n_1208) );
NAND2xp5_ASAP7_75t_L g1209 ( .A(n_1176), .B(n_1113), .Y(n_1209) );
OR2x6_ASAP7_75t_L g1210 ( .A(n_1184), .B(n_1138), .Y(n_1210) );
OAI31xp33_ASAP7_75t_L g1211 ( .A1(n_1179), .A2(n_1142), .A3(n_1135), .B(n_1140), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1212 ( .A(n_1176), .B(n_1114), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1213 ( .A(n_1147), .B(n_1125), .Y(n_1213) );
CKINVDCx16_ASAP7_75t_R g1214 ( .A(n_1174), .Y(n_1214) );
OAI21xp5_ASAP7_75t_L g1215 ( .A1(n_1168), .A2(n_1134), .B(n_1138), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1152), .B(n_1144), .Y(n_1216) );
NOR3xp33_ASAP7_75t_L g1217 ( .A(n_1146), .B(n_1082), .C(n_1136), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1153), .B(n_1144), .Y(n_1218) );
INVxp67_ASAP7_75t_SL g1219 ( .A(n_1182), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1155), .Y(n_1220) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1153), .B(n_1141), .Y(n_1221) );
AND2x4_ASAP7_75t_L g1222 ( .A(n_1188), .B(n_1096), .Y(n_1222) );
AND4x1_ASAP7_75t_L g1223 ( .A(n_1163), .B(n_1121), .C(n_1105), .D(n_1077), .Y(n_1223) );
INVx2_ASAP7_75t_L g1224 ( .A(n_1149), .Y(n_1224) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1161), .Y(n_1225) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1161), .Y(n_1226) );
NOR4xp25_ASAP7_75t_L g1227 ( .A(n_1202), .B(n_1177), .C(n_1172), .D(n_1186), .Y(n_1227) );
NAND2xp5_ASAP7_75t_L g1228 ( .A(n_1201), .B(n_1187), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1229 ( .A(n_1208), .B(n_1187), .Y(n_1229) );
AOI21xp33_ASAP7_75t_L g1230 ( .A1(n_1204), .A2(n_1211), .B(n_1215), .Y(n_1230) );
INVxp67_ASAP7_75t_L g1231 ( .A(n_1197), .Y(n_1231) );
NAND2xp5_ASAP7_75t_L g1232 ( .A(n_1221), .B(n_1181), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1221), .B(n_1158), .Y(n_1233) );
NAND2xp5_ASAP7_75t_L g1234 ( .A(n_1209), .B(n_1181), .Y(n_1234) );
OAI21xp5_ASAP7_75t_SL g1235 ( .A1(n_1217), .A2(n_1157), .B(n_1193), .Y(n_1235) );
AOI22xp5_ASAP7_75t_L g1236 ( .A1(n_1217), .A2(n_1158), .B1(n_1185), .B2(n_1192), .Y(n_1236) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1203), .B(n_1185), .Y(n_1237) );
A2O1A1Ixp33_ASAP7_75t_L g1238 ( .A1(n_1198), .A2(n_1184), .B(n_1188), .C(n_1077), .Y(n_1238) );
NOR2xp33_ASAP7_75t_L g1239 ( .A(n_1214), .B(n_1164), .Y(n_1239) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_1212), .B(n_1175), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1200), .Y(n_1241) );
AOI21xp5_ASAP7_75t_L g1242 ( .A1(n_1210), .A2(n_1191), .B(n_1139), .Y(n_1242) );
OAI21xp5_ASAP7_75t_SL g1243 ( .A1(n_1223), .A2(n_1165), .B(n_1162), .Y(n_1243) );
INVx2_ASAP7_75t_L g1244 ( .A(n_1194), .Y(n_1244) );
NAND2xp5_ASAP7_75t_L g1245 ( .A(n_1234), .B(n_1213), .Y(n_1245) );
OAI211xp5_ASAP7_75t_SL g1246 ( .A1(n_1230), .A2(n_1205), .B(n_1199), .C(n_1219), .Y(n_1246) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1229), .Y(n_1247) );
INVxp67_ASAP7_75t_L g1248 ( .A(n_1239), .Y(n_1248) );
OAI22xp5_ASAP7_75t_L g1249 ( .A1(n_1235), .A2(n_1210), .B1(n_1206), .B2(n_1222), .Y(n_1249) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1241), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g1251 ( .A(n_1228), .B(n_1216), .Y(n_1251) );
INVx2_ASAP7_75t_L g1252 ( .A(n_1244), .Y(n_1252) );
NOR2x1p5_ASAP7_75t_SL g1253 ( .A(n_1227), .B(n_1194), .Y(n_1253) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1231), .Y(n_1254) );
AOI22xp5_ASAP7_75t_L g1255 ( .A1(n_1236), .A2(n_1222), .B1(n_1195), .B2(n_1196), .Y(n_1255) );
AOI21xp5_ASAP7_75t_L g1256 ( .A1(n_1249), .A2(n_1243), .B(n_1238), .Y(n_1256) );
NAND2xp5_ASAP7_75t_L g1257 ( .A(n_1247), .B(n_1237), .Y(n_1257) );
OAI221xp5_ASAP7_75t_L g1258 ( .A1(n_1249), .A2(n_1242), .B1(n_1232), .B2(n_1219), .C(n_1240), .Y(n_1258) );
OAI21xp5_ASAP7_75t_L g1259 ( .A1(n_1246), .A2(n_1233), .B(n_1237), .Y(n_1259) );
AOI221x1_ASAP7_75t_L g1260 ( .A1(n_1254), .A2(n_1182), .B1(n_1183), .B2(n_1207), .C(n_1226), .Y(n_1260) );
AOI221xp5_ASAP7_75t_L g1261 ( .A1(n_1248), .A2(n_1203), .B1(n_1218), .B2(n_1225), .C(n_1220), .Y(n_1261) );
AOI222xp33_ASAP7_75t_L g1262 ( .A1(n_1253), .A2(n_1171), .B1(n_1173), .B2(n_1167), .C1(n_1166), .C2(n_1178), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1263 ( .A(n_1259), .B(n_1255), .Y(n_1263) );
OAI21xp33_ASAP7_75t_SL g1264 ( .A1(n_1262), .A2(n_1251), .B(n_1245), .Y(n_1264) );
OAI22xp33_ASAP7_75t_L g1265 ( .A1(n_1256), .A2(n_1245), .B1(n_1250), .B2(n_1252), .Y(n_1265) );
OAI221xp5_ASAP7_75t_R g1266 ( .A1(n_1258), .A2(n_1196), .B1(n_1195), .B2(n_1156), .C(n_1165), .Y(n_1266) );
OAI21xp33_ASAP7_75t_L g1267 ( .A1(n_1264), .A2(n_1261), .B(n_1257), .Y(n_1267) );
XNOR2x1_ASAP7_75t_L g1268 ( .A(n_1263), .B(n_1074), .Y(n_1268) );
OAI22xp5_ASAP7_75t_L g1269 ( .A1(n_1265), .A2(n_1170), .B1(n_1173), .B2(n_1162), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1268), .B(n_1269), .Y(n_1270) );
OR3x1_ASAP7_75t_L g1271 ( .A(n_1267), .B(n_1266), .C(n_1260), .Y(n_1271) );
AND4x2_ASAP7_75t_L g1272 ( .A(n_1271), .B(n_1133), .C(n_1074), .D(n_1127), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_1270), .B(n_1160), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1273), .Y(n_1274) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1274), .Y(n_1275) );
AO21x2_ASAP7_75t_L g1276 ( .A1(n_1275), .A2(n_1272), .B(n_1189), .Y(n_1276) );
AOI22xp33_ASAP7_75t_L g1277 ( .A1(n_1275), .A2(n_1074), .B1(n_1224), .B2(n_1190), .Y(n_1277) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1276), .Y(n_1278) );
AOI21xp5_ASAP7_75t_L g1279 ( .A1(n_1278), .A2(n_1277), .B(n_1056), .Y(n_1279) );
endmodule