module fake_netlist_5_527_n_1529 (n_137, n_294, n_318, n_380, n_82, n_194, n_316, n_389, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_244, n_47, n_173, n_198, n_247, n_314, n_368, n_8, n_321, n_292, n_100, n_212, n_385, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_341, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_13, n_371, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_267, n_297, n_156, n_5, n_225, n_377, n_219, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_361, n_363, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_359, n_117, n_326, n_233, n_205, n_366, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_391, n_175, n_262, n_238, n_99, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1529);

input n_137;
input n_294;
input n_318;
input n_380;
input n_82;
input n_194;
input n_316;
input n_389;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_368;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_385;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_341;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_13;
input n_371;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_363;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_391;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1529;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_1517;
wire n_976;
wire n_1449;
wire n_1078;
wire n_775;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_955;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_521;
wire n_845;
wire n_663;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_464;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1199;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1233;
wire n_526;
wire n_677;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_689;
wire n_738;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_1163;
wire n_906;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_396;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_486;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_815;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_950;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_507;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_681;
wire n_584;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1419;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_487;
wire n_665;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_1399;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_622;
wire n_1087;
wire n_994;
wire n_848;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1245;
wire n_846;
wire n_465;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_1402;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

INVx1_ASAP7_75t_L g394 ( 
.A(n_223),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_123),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_79),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_285),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_40),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_106),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_113),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_293),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_392),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_37),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_373),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_255),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_151),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_141),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_63),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_273),
.Y(n_409)
);

BUFx2_ASAP7_75t_SL g410 ( 
.A(n_382),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_152),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_101),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_96),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_8),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_221),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_375),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_282),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_367),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_127),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_144),
.Y(n_420)
);

BUFx5_ASAP7_75t_L g421 ( 
.A(n_166),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_24),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_83),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_53),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_388),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_214),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_122),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_391),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_45),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_38),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_107),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_74),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_354),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_84),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_194),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_238),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_341),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_25),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_201),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_37),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_71),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_5),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_350),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_321),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_260),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_43),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_345),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_115),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_234),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_118),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_323),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_253),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_338),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_177),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_167),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_67),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_381),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_126),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_92),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_374),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_0),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_147),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_239),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_209),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_212),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_268),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_163),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_358),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_322),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_91),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_356),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_3),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_332),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_274),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_185),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_328),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_364),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_76),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_376),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_304),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_35),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_237),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_217),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_362),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_288),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_94),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_8),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_219),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_44),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_15),
.Y(n_490)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_284),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_380),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_21),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_38),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_206),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_272),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_7),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_386),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_160),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_184),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_233),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_283),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_143),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_346),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_57),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_174),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_337),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_327),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_31),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_18),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_232),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_336),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_99),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_40),
.Y(n_514)
);

INVx1_ASAP7_75t_SL g515 ( 
.A(n_326),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_222),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_86),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_379),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_267),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_357),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_377),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_295),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_314),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_102),
.Y(n_524)
);

BUFx10_ASAP7_75t_L g525 ( 
.A(n_385),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_258),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_23),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_259),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_134),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g530 ( 
.A(n_80),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_138),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_309),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_378),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_56),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_43),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_306),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_4),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_271),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_352),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_41),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_266),
.Y(n_541)
);

BUFx10_ASAP7_75t_L g542 ( 
.A(n_13),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_11),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_12),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_131),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_299),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_182),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_244),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_162),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_1),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_55),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_192),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_54),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_81),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_4),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_132),
.Y(n_556)
);

BUFx10_ASAP7_75t_L g557 ( 
.A(n_246),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_0),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_130),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_333),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_75),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_110),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_303),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_307),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_108),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_220),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_216),
.Y(n_567)
);

CKINVDCx16_ASAP7_75t_R g568 ( 
.A(n_10),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_275),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_104),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_294),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_47),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_229),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_145),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_53),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_317),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_135),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_87),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_103),
.Y(n_579)
);

BUFx8_ASAP7_75t_SL g580 ( 
.A(n_30),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_360),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_189),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_12),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_264),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_172),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_170),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_225),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_363),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_35),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_77),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_218),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_207),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_197),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_121),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_575),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_414),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_575),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_398),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_403),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_442),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_537),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_461),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_405),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g604 ( 
.A(n_580),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_494),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_396),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_510),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_397),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_496),
.B(n_1),
.Y(n_609)
);

INVxp67_ASAP7_75t_SL g610 ( 
.A(n_576),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_514),
.Y(n_611)
);

NOR2xp67_ASAP7_75t_L g612 ( 
.A(n_550),
.B(n_2),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_555),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_583),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_399),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_400),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_421),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_407),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_408),
.Y(n_619)
);

INVxp67_ASAP7_75t_L g620 ( 
.A(n_542),
.Y(n_620)
);

INVxp67_ASAP7_75t_SL g621 ( 
.A(n_462),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_409),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_417),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_418),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_394),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_568),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_423),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_530),
.B(n_2),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_437),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_401),
.Y(n_630)
);

INVxp33_ASAP7_75t_SL g631 ( 
.A(n_422),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_402),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_426),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_404),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_427),
.Y(n_635)
);

INVxp67_ASAP7_75t_SL g636 ( 
.A(n_420),
.Y(n_636)
);

CKINVDCx16_ASAP7_75t_R g637 ( 
.A(n_432),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_406),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_433),
.Y(n_639)
);

INVxp67_ASAP7_75t_SL g640 ( 
.A(n_478),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_421),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_411),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_439),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_412),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_444),
.Y(n_645)
);

INVxp33_ASAP7_75t_L g646 ( 
.A(n_542),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_445),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_421),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_413),
.B(n_3),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_448),
.Y(n_650)
);

INVxp67_ASAP7_75t_SL g651 ( 
.A(n_569),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_415),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_449),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_451),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_416),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_425),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_452),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_456),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_424),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_457),
.Y(n_660)
);

NOR2xp67_ASAP7_75t_L g661 ( 
.A(n_429),
.B(n_5),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_434),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_471),
.Y(n_663)
);

CKINVDCx16_ASAP7_75t_R g664 ( 
.A(n_498),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_436),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_508),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_443),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_447),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_458),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_460),
.Y(n_670)
);

CKINVDCx14_ASAP7_75t_R g671 ( 
.A(n_525),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_450),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_430),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_453),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_454),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_455),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_525),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_470),
.Y(n_678)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_522),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_463),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_477),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_419),
.B(n_6),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_421),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_464),
.Y(n_684)
);

INVxp67_ASAP7_75t_SL g685 ( 
.A(n_482),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_557),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_465),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_466),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_483),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_488),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_467),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_547),
.Y(n_692)
);

INVxp67_ASAP7_75t_SL g693 ( 
.A(n_492),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_495),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_504),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_395),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_421),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_468),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_628),
.B(n_428),
.Y(n_699)
);

BUFx2_ASAP7_75t_L g700 ( 
.A(n_626),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_696),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_696),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_696),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_625),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_630),
.Y(n_705)
);

HB1xp67_ASAP7_75t_L g706 ( 
.A(n_659),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_632),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_696),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_601),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_634),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_617),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_638),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_598),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_599),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_685),
.B(n_693),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_617),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_642),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_641),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_644),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_641),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_652),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_648),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_600),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_655),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_656),
.B(n_469),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_601),
.Y(n_726)
);

OA21x2_ASAP7_75t_L g727 ( 
.A1(n_648),
.A2(n_512),
.B(n_511),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_636),
.B(n_431),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_662),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_665),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_667),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_640),
.B(n_557),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_602),
.Y(n_733)
);

AND2x6_ASAP7_75t_L g734 ( 
.A(n_683),
.B(n_395),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_628),
.B(n_438),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_605),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_668),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_672),
.Y(n_738)
);

BUFx2_ASAP7_75t_L g739 ( 
.A(n_677),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_674),
.B(n_473),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_675),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_651),
.B(n_441),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_607),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_683),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_676),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_611),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_697),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_678),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_681),
.Y(n_749)
);

HB1xp67_ASAP7_75t_L g750 ( 
.A(n_620),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_677),
.B(n_548),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_686),
.B(n_565),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_649),
.B(n_440),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_689),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_613),
.Y(n_755)
);

BUFx2_ASAP7_75t_L g756 ( 
.A(n_686),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_614),
.Y(n_757)
);

OA21x2_ASAP7_75t_L g758 ( 
.A1(n_697),
.A2(n_521),
.B(n_518),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_690),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_596),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_694),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_695),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_606),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_595),
.B(n_523),
.Y(n_764)
);

CKINVDCx8_ASAP7_75t_R g765 ( 
.A(n_664),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_673),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_608),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_609),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_612),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_610),
.Y(n_770)
);

BUFx8_ASAP7_75t_L g771 ( 
.A(n_671),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_609),
.B(n_474),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_621),
.B(n_594),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_SL g774 ( 
.A1(n_646),
.A2(n_481),
.B1(n_472),
.B2(n_446),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_649),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_682),
.Y(n_776)
);

AND2x4_ASAP7_75t_L g777 ( 
.A(n_597),
.B(n_524),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_682),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_615),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_616),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_661),
.B(n_487),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_618),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_619),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_622),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_623),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_760),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_742),
.B(n_637),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_760),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_711),
.B(n_421),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_751),
.B(n_577),
.Y(n_790)
);

INVx4_ASAP7_75t_L g791 ( 
.A(n_762),
.Y(n_791)
);

INVx6_ASAP7_75t_L g792 ( 
.A(n_771),
.Y(n_792)
);

BUFx4f_ASAP7_75t_L g793 ( 
.A(n_782),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_704),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_732),
.B(n_624),
.Y(n_795)
);

NAND2xp33_ASAP7_75t_L g796 ( 
.A(n_768),
.B(n_627),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_699),
.B(n_633),
.Y(n_797)
);

INVxp67_ASAP7_75t_L g798 ( 
.A(n_750),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_699),
.B(n_635),
.Y(n_799)
);

CKINVDCx8_ASAP7_75t_R g800 ( 
.A(n_783),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_703),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_705),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_772),
.B(n_639),
.Y(n_803)
);

AND2x4_ASAP7_75t_L g804 ( 
.A(n_751),
.B(n_528),
.Y(n_804)
);

INVx5_ASAP7_75t_L g805 ( 
.A(n_734),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_772),
.B(n_643),
.Y(n_806)
);

INVx4_ASAP7_75t_L g807 ( 
.A(n_762),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_703),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_702),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_702),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_707),
.Y(n_811)
);

OAI22xp33_ASAP7_75t_L g812 ( 
.A1(n_775),
.A2(n_490),
.B1(n_493),
.B2(n_489),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_780),
.B(n_631),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_739),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_701),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_756),
.Y(n_816)
);

OAI221xp5_ASAP7_75t_L g817 ( 
.A1(n_768),
.A2(n_516),
.B1(n_515),
.B2(n_491),
.C(n_531),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_710),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_702),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_780),
.B(n_645),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_701),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_784),
.B(n_647),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_708),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_708),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_706),
.B(n_650),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_712),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_711),
.B(n_653),
.Y(n_827)
);

INVxp33_ASAP7_75t_L g828 ( 
.A(n_750),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_776),
.A2(n_410),
.B1(n_435),
.B2(n_395),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_706),
.B(n_654),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_702),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_716),
.B(n_657),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_766),
.B(n_658),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_778),
.B(n_660),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_723),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_716),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_717),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_735),
.A2(n_435),
.B1(n_459),
.B2(n_395),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_719),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_771),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_721),
.Y(n_841)
);

INVxp67_ASAP7_75t_SL g842 ( 
.A(n_727),
.Y(n_842)
);

BUFx10_ASAP7_75t_L g843 ( 
.A(n_752),
.Y(n_843)
);

CKINVDCx20_ASAP7_75t_R g844 ( 
.A(n_765),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_715),
.B(n_728),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_763),
.B(n_669),
.Y(n_846)
);

NAND3xp33_ASAP7_75t_L g847 ( 
.A(n_715),
.B(n_534),
.C(n_532),
.Y(n_847)
);

INVx4_ASAP7_75t_L g848 ( 
.A(n_762),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_724),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_SL g850 ( 
.A(n_774),
.B(n_497),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_763),
.B(n_670),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_735),
.A2(n_527),
.B1(n_535),
.B2(n_509),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_718),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_700),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_784),
.B(n_680),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_723),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_779),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_770),
.B(n_684),
.Y(n_858)
);

NAND2xp33_ASAP7_75t_SL g859 ( 
.A(n_753),
.B(n_540),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_729),
.Y(n_860)
);

BUFx10_ASAP7_75t_L g861 ( 
.A(n_752),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_718),
.B(n_687),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_720),
.B(n_688),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_785),
.B(n_545),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_753),
.A2(n_544),
.B1(n_558),
.B2(n_543),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_730),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_731),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_728),
.B(n_691),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_764),
.A2(n_459),
.B1(n_541),
.B2(n_435),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_720),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_769),
.B(n_698),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_773),
.B(n_475),
.Y(n_872)
);

BUFx4f_ASAP7_75t_L g873 ( 
.A(n_779),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_722),
.B(n_553),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_722),
.A2(n_559),
.B(n_567),
.C(n_556),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_744),
.B(n_570),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_785),
.B(n_604),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_744),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_737),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_794),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_803),
.B(n_773),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_836),
.Y(n_882)
);

AO22x2_ASAP7_75t_L g883 ( 
.A1(n_797),
.A2(n_777),
.B1(n_764),
.B2(n_781),
.Y(n_883)
);

NAND2x1p5_ASAP7_75t_L g884 ( 
.A(n_873),
.B(n_767),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_802),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_811),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_818),
.Y(n_887)
);

CKINVDCx20_ASAP7_75t_R g888 ( 
.A(n_844),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_826),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_837),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_873),
.B(n_725),
.Y(n_891)
);

AO22x2_ASAP7_75t_L g892 ( 
.A1(n_799),
.A2(n_777),
.B1(n_781),
.B2(n_579),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_853),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_787),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_806),
.B(n_725),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_795),
.B(n_740),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_798),
.B(n_740),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_845),
.A2(n_629),
.B1(n_663),
.B2(n_603),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_842),
.B(n_762),
.Y(n_899)
);

AO22x2_ASAP7_75t_L g900 ( 
.A1(n_834),
.A2(n_582),
.B1(n_584),
.B2(n_574),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_839),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_841),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_820),
.B(n_747),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_822),
.B(n_855),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_849),
.Y(n_905)
);

AO22x2_ASAP7_75t_L g906 ( 
.A1(n_847),
.A2(n_587),
.B1(n_592),
.B2(n_586),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_870),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_786),
.B(n_788),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_860),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_866),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_828),
.B(n_666),
.Y(n_911)
);

NAND2x1p5_ASAP7_75t_L g912 ( 
.A(n_868),
.B(n_709),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_878),
.Y(n_913)
);

AO22x2_ASAP7_75t_L g914 ( 
.A1(n_847),
.A2(n_741),
.B1(n_745),
.B2(n_738),
.Y(n_914)
);

BUFx8_ASAP7_75t_L g915 ( 
.A(n_825),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_867),
.Y(n_916)
);

NAND2x1p5_ASAP7_75t_L g917 ( 
.A(n_816),
.B(n_793),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_879),
.Y(n_918)
);

OAI221xp5_ASAP7_75t_L g919 ( 
.A1(n_817),
.A2(n_754),
.B1(n_761),
.B2(n_749),
.C(n_748),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_815),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_821),
.Y(n_921)
);

INVxp67_ASAP7_75t_L g922 ( 
.A(n_854),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_804),
.B(n_679),
.Y(n_923)
);

AO22x2_ASAP7_75t_L g924 ( 
.A1(n_790),
.A2(n_692),
.B1(n_9),
.B2(n_6),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_800),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_823),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_830),
.B(n_709),
.Y(n_927)
);

AO22x2_ASAP7_75t_L g928 ( 
.A1(n_790),
.A2(n_10),
.B1(n_7),
.B2(n_9),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_872),
.B(n_747),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_827),
.B(n_727),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_824),
.Y(n_931)
);

AO22x2_ASAP7_75t_L g932 ( 
.A1(n_814),
.A2(n_833),
.B1(n_864),
.B2(n_804),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_864),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_801),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_827),
.B(n_727),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_808),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_793),
.A2(n_479),
.B1(n_480),
.B2(n_476),
.Y(n_937)
);

OAI221xp5_ASAP7_75t_L g938 ( 
.A1(n_852),
.A2(n_759),
.B1(n_713),
.B2(n_757),
.C(n_733),
.Y(n_938)
);

BUFx8_ASAP7_75t_L g939 ( 
.A(n_871),
.Y(n_939)
);

AO22x2_ASAP7_75t_L g940 ( 
.A1(n_858),
.A2(n_14),
.B1(n_11),
.B2(n_13),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_832),
.B(n_862),
.Y(n_941)
);

NAND2x1p5_ASAP7_75t_L g942 ( 
.A(n_846),
.B(n_726),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_789),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_789),
.Y(n_944)
);

NAND2x1p5_ASAP7_75t_L g945 ( 
.A(n_851),
.B(n_726),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_874),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_832),
.B(n_714),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_796),
.A2(n_485),
.B1(n_486),
.B2(n_484),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_810),
.Y(n_949)
);

AO22x2_ASAP7_75t_L g950 ( 
.A1(n_850),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_862),
.B(n_758),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_874),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_876),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_829),
.A2(n_500),
.B1(n_501),
.B2(n_499),
.Y(n_954)
);

AO22x2_ASAP7_75t_L g955 ( 
.A1(n_812),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_863),
.B(n_758),
.Y(n_956)
);

AO22x2_ASAP7_75t_L g957 ( 
.A1(n_863),
.A2(n_20),
.B1(n_17),
.B2(n_19),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_859),
.A2(n_503),
.B1(n_505),
.B2(n_502),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_876),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_813),
.B(n_835),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_810),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_843),
.Y(n_962)
);

NAND2xp33_ASAP7_75t_L g963 ( 
.A(n_838),
.B(n_506),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_857),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_809),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_835),
.B(n_758),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_843),
.Y(n_967)
);

AO22x2_ASAP7_75t_L g968 ( 
.A1(n_852),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_968)
);

OAI221xp5_ASAP7_75t_L g969 ( 
.A1(n_865),
.A2(n_746),
.B1(n_589),
.B2(n_572),
.C(n_736),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_861),
.Y(n_970)
);

BUFx8_ASAP7_75t_L g971 ( 
.A(n_792),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_861),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_831),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_809),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_856),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_856),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_865),
.A2(n_746),
.B(n_513),
.C(n_517),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_809),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_819),
.Y(n_979)
);

NAND2xp33_ASAP7_75t_SL g980 ( 
.A(n_904),
.B(n_840),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_908),
.B(n_877),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_881),
.B(n_895),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_941),
.B(n_805),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_897),
.B(n_805),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_927),
.B(n_805),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_946),
.B(n_791),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_947),
.B(n_791),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_960),
.B(n_807),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_896),
.B(n_807),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_894),
.B(n_848),
.Y(n_990)
);

NAND2xp33_ASAP7_75t_SL g991 ( 
.A(n_925),
.B(n_869),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_884),
.B(n_848),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_952),
.B(n_723),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_953),
.B(n_723),
.Y(n_994)
);

NAND2xp33_ASAP7_75t_SL g995 ( 
.A(n_964),
.B(n_962),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_959),
.B(n_736),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_933),
.B(n_736),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_903),
.B(n_819),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_891),
.B(n_736),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_917),
.B(n_743),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_880),
.B(n_743),
.Y(n_1001)
);

NAND2xp33_ASAP7_75t_SL g1002 ( 
.A(n_967),
.B(n_507),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_885),
.B(n_743),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_886),
.B(n_743),
.Y(n_1004)
);

NAND2xp33_ASAP7_75t_SL g1005 ( 
.A(n_970),
.B(n_519),
.Y(n_1005)
);

NAND2xp33_ASAP7_75t_SL g1006 ( 
.A(n_972),
.B(n_520),
.Y(n_1006)
);

NAND2xp33_ASAP7_75t_SL g1007 ( 
.A(n_923),
.B(n_526),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_887),
.B(n_755),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_889),
.B(n_755),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_890),
.B(n_755),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_901),
.B(n_902),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_905),
.B(n_755),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_909),
.B(n_819),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_943),
.B(n_529),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_910),
.B(n_916),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_911),
.B(n_792),
.Y(n_1016)
);

NAND2xp33_ASAP7_75t_SL g1017 ( 
.A(n_888),
.B(n_533),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_918),
.B(n_536),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_898),
.B(n_538),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_944),
.B(n_899),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_922),
.B(n_539),
.Y(n_1021)
);

NAND2xp33_ASAP7_75t_SL g1022 ( 
.A(n_930),
.B(n_546),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_912),
.B(n_549),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_977),
.B(n_551),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_948),
.B(n_552),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_958),
.B(n_554),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_929),
.B(n_560),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_942),
.B(n_561),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_945),
.B(n_562),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_937),
.B(n_563),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_934),
.B(n_564),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_935),
.B(n_566),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_936),
.B(n_571),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_932),
.B(n_578),
.Y(n_1034)
);

NAND2xp33_ASAP7_75t_SL g1035 ( 
.A(n_951),
.B(n_581),
.Y(n_1035)
);

AND3x1_ASAP7_75t_L g1036 ( 
.A(n_924),
.B(n_875),
.C(n_22),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_954),
.B(n_585),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_956),
.B(n_588),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_932),
.B(n_590),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_882),
.B(n_591),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_893),
.B(n_593),
.Y(n_1041)
);

NAND2xp33_ASAP7_75t_SL g1042 ( 
.A(n_965),
.B(n_435),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_907),
.B(n_459),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_883),
.B(n_734),
.Y(n_1044)
);

NAND2xp33_ASAP7_75t_SL g1045 ( 
.A(n_974),
.B(n_459),
.Y(n_1045)
);

NAND2xp33_ASAP7_75t_SL g1046 ( 
.A(n_978),
.B(n_541),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_914),
.B(n_22),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_883),
.B(n_734),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_913),
.B(n_58),
.Y(n_1049)
);

NAND2xp33_ASAP7_75t_SL g1050 ( 
.A(n_979),
.B(n_541),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_921),
.B(n_541),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_926),
.B(n_573),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_931),
.B(n_573),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_914),
.B(n_734),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_966),
.B(n_573),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_982),
.A2(n_938),
.B(n_969),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_981),
.B(n_1016),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_1020),
.A2(n_976),
.B(n_975),
.Y(n_1058)
);

INVx2_ASAP7_75t_SL g1059 ( 
.A(n_981),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_L g1060 ( 
.A1(n_1055),
.A2(n_961),
.B(n_949),
.Y(n_1060)
);

AO31x2_ASAP7_75t_L g1061 ( 
.A1(n_1044),
.A2(n_973),
.A3(n_920),
.B(n_892),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_1011),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1014),
.B(n_892),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_991),
.A2(n_919),
.B(n_963),
.C(n_900),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_1015),
.B(n_939),
.Y(n_1065)
);

CKINVDCx8_ASAP7_75t_R g1066 ( 
.A(n_1049),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_1019),
.B(n_915),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_1021),
.B(n_971),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_1055),
.A2(n_906),
.B(n_900),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_1034),
.B(n_928),
.Y(n_1070)
);

CKINVDCx20_ASAP7_75t_R g1071 ( 
.A(n_1017),
.Y(n_1071)
);

NOR3xp33_ASAP7_75t_SL g1072 ( 
.A(n_980),
.B(n_940),
.C(n_968),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1049),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1027),
.B(n_906),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_998),
.Y(n_1075)
);

INVx3_ASAP7_75t_SL g1076 ( 
.A(n_1047),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_986),
.A2(n_940),
.B1(n_928),
.B2(n_968),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1032),
.B(n_955),
.Y(n_1078)
);

AO21x2_ASAP7_75t_L g1079 ( 
.A1(n_1038),
.A2(n_957),
.B(n_955),
.Y(n_1079)
);

NAND3xp33_ASAP7_75t_SL g1080 ( 
.A(n_1039),
.B(n_950),
.C(n_957),
.Y(n_1080)
);

HB1xp67_ASAP7_75t_L g1081 ( 
.A(n_997),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_1054),
.A2(n_60),
.B(n_59),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_SL g1083 ( 
.A1(n_992),
.A2(n_573),
.B(n_734),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_988),
.A2(n_950),
.B(n_62),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_1048),
.A2(n_64),
.B(n_61),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_SL g1086 ( 
.A1(n_989),
.A2(n_66),
.B(n_65),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_1031),
.Y(n_1087)
);

NAND2xp33_ASAP7_75t_L g1088 ( 
.A(n_1028),
.B(n_68),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_983),
.A2(n_70),
.B(n_69),
.Y(n_1089)
);

AOI221xp5_ASAP7_75t_L g1090 ( 
.A1(n_1036),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.C(n_26),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_987),
.B(n_26),
.Y(n_1091)
);

AOI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_993),
.A2(n_73),
.B1(n_78),
.B2(n_72),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_985),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_994),
.B(n_27),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_996),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_999),
.A2(n_85),
.B(n_82),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1018),
.B(n_27),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_1013),
.A2(n_1003),
.B(n_1001),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1022),
.A2(n_89),
.B(n_88),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1035),
.A2(n_93),
.B(n_90),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_995),
.B(n_95),
.Y(n_1101)
);

OA21x2_ASAP7_75t_L g1102 ( 
.A1(n_1024),
.A2(n_98),
.B(n_97),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1037),
.A2(n_105),
.B(n_100),
.Y(n_1103)
);

AOI221xp5_ASAP7_75t_SL g1104 ( 
.A1(n_984),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.C(n_31),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_990),
.B(n_28),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_1004),
.A2(n_111),
.B(n_109),
.Y(n_1106)
);

NAND3x1_ASAP7_75t_L g1107 ( 
.A(n_1007),
.B(n_29),
.C(n_32),
.Y(n_1107)
);

NOR3xp33_ASAP7_75t_L g1108 ( 
.A(n_1002),
.B(n_32),
.C(n_33),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_SL g1109 ( 
.A(n_1000),
.B(n_112),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_1023),
.B(n_114),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1029),
.B(n_33),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1025),
.A2(n_247),
.B1(n_390),
.B2(n_389),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1033),
.B(n_34),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1040),
.B(n_34),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1008),
.B(n_36),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_1005),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1041),
.B(n_36),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1030),
.A2(n_117),
.B(n_116),
.Y(n_1118)
);

BUFx3_ASAP7_75t_L g1119 ( 
.A(n_1059),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_1060),
.A2(n_1010),
.B(n_1009),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_SL g1121 ( 
.A1(n_1084),
.A2(n_1012),
.B(n_1046),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_1073),
.B(n_1026),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_1057),
.B(n_1006),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_1064),
.A2(n_1050),
.B(n_1053),
.C(n_1051),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_1076),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_1066),
.Y(n_1126)
);

OA21x2_ASAP7_75t_L g1127 ( 
.A1(n_1058),
.A2(n_1052),
.B(n_1043),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1089),
.A2(n_1045),
.B(n_1042),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_1062),
.Y(n_1129)
);

INVx1_ASAP7_75t_SL g1130 ( 
.A(n_1078),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_1093),
.B(n_119),
.Y(n_1131)
);

NAND3xp33_ASAP7_75t_L g1132 ( 
.A(n_1090),
.B(n_39),
.C(n_41),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1075),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_1093),
.B(n_120),
.Y(n_1134)
);

NAND4xp25_ASAP7_75t_L g1135 ( 
.A(n_1068),
.B(n_39),
.C(n_42),
.D(n_44),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1096),
.A2(n_1082),
.B(n_1098),
.Y(n_1136)
);

OR2x2_ASAP7_75t_L g1137 ( 
.A(n_1074),
.B(n_42),
.Y(n_1137)
);

NOR2xp67_ASAP7_75t_L g1138 ( 
.A(n_1087),
.B(n_124),
.Y(n_1138)
);

INVxp67_ASAP7_75t_L g1139 ( 
.A(n_1065),
.Y(n_1139)
);

OA21x2_ASAP7_75t_L g1140 ( 
.A1(n_1056),
.A2(n_128),
.B(n_125),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1070),
.B(n_45),
.Y(n_1141)
);

AND2x4_ASAP7_75t_L g1142 ( 
.A(n_1065),
.B(n_129),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1063),
.B(n_46),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1106),
.A2(n_136),
.B(n_133),
.Y(n_1144)
);

OA21x2_ASAP7_75t_L g1145 ( 
.A1(n_1056),
.A2(n_139),
.B(n_137),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_1071),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1115),
.B(n_1072),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1081),
.Y(n_1148)
);

INVx3_ASAP7_75t_L g1149 ( 
.A(n_1061),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1077),
.B(n_46),
.Y(n_1150)
);

AOI21xp33_ASAP7_75t_L g1151 ( 
.A1(n_1079),
.A2(n_47),
.B(n_48),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1095),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1069),
.A2(n_142),
.B(n_140),
.Y(n_1153)
);

BUFx12f_ASAP7_75t_L g1154 ( 
.A(n_1116),
.Y(n_1154)
);

OR2x6_ASAP7_75t_L g1155 ( 
.A(n_1086),
.B(n_146),
.Y(n_1155)
);

O2A1O1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1108),
.A2(n_48),
.B(n_49),
.C(n_50),
.Y(n_1156)
);

AO21x1_ASAP7_75t_L g1157 ( 
.A1(n_1085),
.A2(n_49),
.B(n_50),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1099),
.A2(n_149),
.B(n_148),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1079),
.B(n_51),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1100),
.A2(n_153),
.B(n_150),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1061),
.Y(n_1161)
);

NOR2xp67_ASAP7_75t_L g1162 ( 
.A(n_1091),
.B(n_154),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1061),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_1103),
.A2(n_51),
.B(n_52),
.C(n_155),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_1105),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1094),
.A2(n_157),
.B(n_156),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1080),
.A2(n_52),
.B1(n_158),
.B2(n_159),
.Y(n_1167)
);

BUFx3_ASAP7_75t_L g1168 ( 
.A(n_1067),
.Y(n_1168)
);

INVx2_ASAP7_75t_SL g1169 ( 
.A(n_1111),
.Y(n_1169)
);

INVx1_ASAP7_75t_SL g1170 ( 
.A(n_1114),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1102),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1097),
.B(n_393),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_1113),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1117),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1118),
.A2(n_161),
.B(n_164),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_1110),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1101),
.B(n_165),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1163),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1133),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1129),
.Y(n_1180)
);

O2A1O1Ixp33_ASAP7_75t_SL g1181 ( 
.A1(n_1164),
.A2(n_1112),
.B(n_1092),
.C(n_1104),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_1131),
.Y(n_1182)
);

OR2x2_ASAP7_75t_L g1183 ( 
.A(n_1130),
.B(n_1102),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1152),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1143),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1143),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_1119),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1161),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1149),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1141),
.B(n_1104),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1148),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1159),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1174),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1130),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1170),
.B(n_1107),
.Y(n_1195)
);

INVx4_ASAP7_75t_L g1196 ( 
.A(n_1126),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_1146),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1170),
.B(n_1092),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1136),
.A2(n_1083),
.B(n_1088),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1165),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1169),
.Y(n_1201)
);

AO21x2_ASAP7_75t_L g1202 ( 
.A1(n_1171),
.A2(n_1109),
.B(n_168),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1137),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1147),
.B(n_1109),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1131),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_1126),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_1154),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1122),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1122),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1149),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1150),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1134),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_1176),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1140),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1134),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1162),
.Y(n_1216)
);

BUFx8_ASAP7_75t_SL g1217 ( 
.A(n_1126),
.Y(n_1217)
);

AOI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1120),
.A2(n_1121),
.B(n_1127),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1140),
.Y(n_1219)
);

OR2x2_ASAP7_75t_L g1220 ( 
.A(n_1173),
.B(n_169),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1123),
.B(n_387),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_1142),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1145),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1162),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1132),
.A2(n_171),
.B1(n_173),
.B2(n_175),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1145),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1138),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_1125),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1138),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1142),
.B(n_176),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1153),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1157),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1124),
.A2(n_178),
.B(n_179),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_1127),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_1139),
.Y(n_1235)
);

OR2x6_ASAP7_75t_L g1236 ( 
.A(n_1155),
.B(n_180),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_1155),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1144),
.Y(n_1238)
);

OA21x2_ASAP7_75t_L g1239 ( 
.A1(n_1151),
.A2(n_181),
.B(n_183),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_1168),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1132),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1158),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1160),
.Y(n_1243)
);

AOI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1128),
.A2(n_186),
.B(n_187),
.Y(n_1244)
);

INVxp67_ASAP7_75t_L g1245 ( 
.A(n_1172),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_1155),
.Y(n_1246)
);

INVxp67_ASAP7_75t_R g1247 ( 
.A(n_1175),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1177),
.Y(n_1248)
);

NAND2xp33_ASAP7_75t_R g1249 ( 
.A(n_1197),
.B(n_1166),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1204),
.B(n_1167),
.Y(n_1250)
);

NAND2xp33_ASAP7_75t_R g1251 ( 
.A(n_1197),
.B(n_1166),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_R g1252 ( 
.A(n_1207),
.B(n_188),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_R g1253 ( 
.A(n_1207),
.B(n_190),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_R g1254 ( 
.A(n_1206),
.B(n_191),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1203),
.B(n_1208),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_R g1256 ( 
.A(n_1206),
.B(n_193),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_1182),
.B(n_195),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1211),
.B(n_1156),
.Y(n_1258)
);

NAND2xp33_ASAP7_75t_R g1259 ( 
.A(n_1187),
.B(n_196),
.Y(n_1259)
);

NAND2xp33_ASAP7_75t_R g1260 ( 
.A(n_1228),
.B(n_198),
.Y(n_1260)
);

INVxp67_ASAP7_75t_L g1261 ( 
.A(n_1201),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_1240),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1182),
.B(n_1205),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1185),
.B(n_1135),
.Y(n_1264)
);

XNOR2xp5_ASAP7_75t_L g1265 ( 
.A(n_1240),
.B(n_1135),
.Y(n_1265)
);

BUFx3_ASAP7_75t_L g1266 ( 
.A(n_1217),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1205),
.B(n_199),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1209),
.B(n_1151),
.Y(n_1268)
);

OR2x6_ASAP7_75t_L g1269 ( 
.A(n_1236),
.B(n_1237),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1245),
.B(n_200),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1194),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_1212),
.B(n_202),
.Y(n_1272)
);

OR2x6_ASAP7_75t_L g1273 ( 
.A(n_1236),
.B(n_203),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_R g1274 ( 
.A(n_1222),
.B(n_204),
.Y(n_1274)
);

INVxp67_ASAP7_75t_L g1275 ( 
.A(n_1180),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1186),
.B(n_205),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1188),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1188),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1245),
.B(n_208),
.Y(n_1279)
);

INVx3_ASAP7_75t_L g1280 ( 
.A(n_1196),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1198),
.B(n_210),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_R g1282 ( 
.A(n_1222),
.B(n_211),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1192),
.B(n_213),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1217),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1193),
.B(n_215),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_SL g1286 ( 
.A(n_1221),
.B(n_224),
.Y(n_1286)
);

NAND2xp33_ASAP7_75t_R g1287 ( 
.A(n_1230),
.B(n_1246),
.Y(n_1287)
);

CKINVDCx12_ASAP7_75t_R g1288 ( 
.A(n_1220),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1227),
.B(n_1229),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1222),
.B(n_226),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1184),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1196),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_R g1293 ( 
.A(n_1222),
.B(n_1246),
.Y(n_1293)
);

NAND2xp33_ASAP7_75t_R g1294 ( 
.A(n_1236),
.B(n_227),
.Y(n_1294)
);

NAND2xp33_ASAP7_75t_SL g1295 ( 
.A(n_1225),
.B(n_228),
.Y(n_1295)
);

NAND2xp33_ASAP7_75t_R g1296 ( 
.A(n_1235),
.B(n_230),
.Y(n_1296)
);

NAND2xp33_ASAP7_75t_R g1297 ( 
.A(n_1195),
.B(n_231),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1191),
.Y(n_1298)
);

XNOR2xp5_ASAP7_75t_L g1299 ( 
.A(n_1213),
.B(n_384),
.Y(n_1299)
);

NAND2xp33_ASAP7_75t_R g1300 ( 
.A(n_1190),
.B(n_235),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1215),
.B(n_236),
.Y(n_1301)
);

INVxp67_ASAP7_75t_L g1302 ( 
.A(n_1200),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1248),
.B(n_240),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1241),
.B(n_241),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1178),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1213),
.B(n_242),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1184),
.B(n_243),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1179),
.B(n_1196),
.Y(n_1308)
);

INVxp67_ASAP7_75t_L g1309 ( 
.A(n_1216),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1237),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1224),
.B(n_245),
.Y(n_1311)
);

CKINVDCx8_ASAP7_75t_R g1312 ( 
.A(n_1237),
.Y(n_1312)
);

INVx1_ASAP7_75t_SL g1313 ( 
.A(n_1262),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1277),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1278),
.Y(n_1315)
);

AND2x4_ASAP7_75t_SL g1316 ( 
.A(n_1269),
.B(n_1237),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1302),
.B(n_1232),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1275),
.B(n_1183),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1255),
.B(n_1242),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1308),
.B(n_1242),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1305),
.B(n_1189),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1271),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1298),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1264),
.B(n_1178),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1261),
.Y(n_1325)
);

NAND2x1_ASAP7_75t_L g1326 ( 
.A(n_1269),
.B(n_1189),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1268),
.B(n_1210),
.Y(n_1327)
);

INVxp67_ASAP7_75t_SL g1328 ( 
.A(n_1309),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1291),
.Y(n_1329)
);

INVx1_ASAP7_75t_SL g1330 ( 
.A(n_1292),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1289),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1263),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1258),
.B(n_1234),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1281),
.B(n_1210),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1295),
.A2(n_1225),
.B1(n_1250),
.B2(n_1273),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1293),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1306),
.B(n_1234),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1310),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1285),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1263),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1273),
.A2(n_1239),
.B1(n_1233),
.B2(n_1202),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1304),
.B(n_1214),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1312),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_L g1344 ( 
.A(n_1287),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1270),
.B(n_1239),
.Y(n_1345)
);

INVx1_ASAP7_75t_SL g1346 ( 
.A(n_1265),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1307),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1280),
.B(n_1214),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1283),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1279),
.B(n_1299),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1276),
.B(n_1219),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1303),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1311),
.B(n_1219),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1301),
.B(n_1239),
.Y(n_1354)
);

NOR2x1_ASAP7_75t_L g1355 ( 
.A(n_1266),
.B(n_1202),
.Y(n_1355)
);

OR2x6_ASAP7_75t_SL g1356 ( 
.A(n_1294),
.B(n_1243),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1288),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1286),
.A2(n_1181),
.B1(n_1226),
.B2(n_1223),
.Y(n_1358)
);

BUFx8_ASAP7_75t_L g1359 ( 
.A(n_1284),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1272),
.B(n_1223),
.Y(n_1360)
);

CKINVDCx20_ASAP7_75t_R g1361 ( 
.A(n_1252),
.Y(n_1361)
);

INVx2_ASAP7_75t_SL g1362 ( 
.A(n_1322),
.Y(n_1362)
);

INVxp67_ASAP7_75t_L g1363 ( 
.A(n_1325),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1323),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1315),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1315),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1320),
.B(n_1226),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1335),
.A2(n_1344),
.B1(n_1352),
.B2(n_1349),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_1359),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1319),
.B(n_1218),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1359),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1323),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1337),
.B(n_1243),
.Y(n_1373)
);

INVx2_ASAP7_75t_SL g1374 ( 
.A(n_1322),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1314),
.Y(n_1375)
);

NOR2xp67_ASAP7_75t_L g1376 ( 
.A(n_1344),
.B(n_1231),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1345),
.B(n_1247),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1314),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1335),
.A2(n_1249),
.B1(n_1251),
.B2(n_1300),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1327),
.B(n_1238),
.Y(n_1380)
);

AOI33xp33_ASAP7_75t_L g1381 ( 
.A1(n_1339),
.A2(n_1181),
.A3(n_1301),
.B1(n_1272),
.B2(n_1297),
.B3(n_1257),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1314),
.B(n_1238),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1329),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1329),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1356),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1332),
.B(n_1244),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1332),
.B(n_1340),
.Y(n_1387)
);

AND2x4_ASAP7_75t_SL g1388 ( 
.A(n_1336),
.B(n_1257),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1321),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1325),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1317),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1333),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1321),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1321),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1385),
.B(n_1340),
.Y(n_1395)
);

AND2x4_ASAP7_75t_SL g1396 ( 
.A(n_1380),
.B(n_1336),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1392),
.B(n_1318),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_1392),
.B(n_1363),
.Y(n_1398)
);

AND2x4_ASAP7_75t_L g1399 ( 
.A(n_1385),
.B(n_1328),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1389),
.B(n_1393),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1387),
.B(n_1357),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1387),
.B(n_1313),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1389),
.B(n_1338),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1365),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1393),
.B(n_1330),
.Y(n_1405)
);

NOR2x1_ASAP7_75t_SL g1406 ( 
.A(n_1362),
.B(n_1331),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1394),
.B(n_1331),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1394),
.B(n_1354),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1390),
.B(n_1362),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1364),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1391),
.B(n_1342),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1364),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1374),
.B(n_1351),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1372),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1391),
.B(n_1324),
.Y(n_1415)
);

OAI221xp5_ASAP7_75t_L g1416 ( 
.A1(n_1415),
.A2(n_1379),
.B1(n_1368),
.B2(n_1260),
.C(n_1296),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1410),
.Y(n_1417)
);

AND2x4_ASAP7_75t_SL g1418 ( 
.A(n_1399),
.B(n_1361),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1399),
.B(n_1370),
.Y(n_1419)
);

OAI221xp5_ASAP7_75t_L g1420 ( 
.A1(n_1415),
.A2(n_1259),
.B1(n_1411),
.B2(n_1397),
.C(n_1346),
.Y(n_1420)
);

NOR2x1_ASAP7_75t_L g1421 ( 
.A(n_1399),
.B(n_1369),
.Y(n_1421)
);

AO221x2_ASAP7_75t_L g1422 ( 
.A1(n_1411),
.A2(n_1343),
.B1(n_1412),
.B2(n_1414),
.C(n_1406),
.Y(n_1422)
);

NOR2x1_ASAP7_75t_L g1423 ( 
.A(n_1398),
.B(n_1369),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1395),
.B(n_1371),
.Y(n_1424)
);

AO221x2_ASAP7_75t_L g1425 ( 
.A1(n_1404),
.A2(n_1372),
.B1(n_1381),
.B2(n_1371),
.C(n_1378),
.Y(n_1425)
);

OAI31xp33_ASAP7_75t_SL g1426 ( 
.A1(n_1395),
.A2(n_1350),
.A3(n_1355),
.B(n_1377),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1407),
.B(n_1402),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_SL g1428 ( 
.A(n_1405),
.B(n_1376),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1425),
.B(n_1401),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1416),
.A2(n_1341),
.B1(n_1396),
.B2(n_1388),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1419),
.B(n_1427),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1423),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1422),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1425),
.B(n_1413),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1417),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1418),
.B(n_1359),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1421),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1424),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1428),
.Y(n_1439)
);

OAI21xp33_ASAP7_75t_SL g1440 ( 
.A1(n_1426),
.A2(n_1374),
.B(n_1403),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1420),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1425),
.B(n_1408),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1425),
.B(n_1409),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1435),
.Y(n_1444)
);

OAI222xp33_ASAP7_75t_L g1445 ( 
.A1(n_1433),
.A2(n_1377),
.B1(n_1341),
.B2(n_1358),
.C1(n_1400),
.C2(n_1353),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1441),
.B(n_1396),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1432),
.A2(n_1361),
.B(n_1388),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1431),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1438),
.B(n_1404),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1434),
.B(n_1383),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1443),
.B(n_1370),
.Y(n_1451)
);

INVx3_ASAP7_75t_L g1452 ( 
.A(n_1437),
.Y(n_1452)
);

CKINVDCx16_ASAP7_75t_R g1453 ( 
.A(n_1448),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1452),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1444),
.Y(n_1455)
);

NOR2xp33_ASAP7_75t_L g1456 ( 
.A(n_1447),
.B(n_1436),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1449),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1450),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1452),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1453),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1455),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1457),
.B(n_1446),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1456),
.B(n_1439),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1454),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1458),
.Y(n_1465)
);

INVx4_ASAP7_75t_L g1466 ( 
.A(n_1459),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1460),
.B(n_1451),
.Y(n_1467)
);

NAND4xp25_ASAP7_75t_L g1468 ( 
.A(n_1463),
.B(n_1430),
.C(n_1429),
.D(n_1442),
.Y(n_1468)
);

OAI211xp5_ASAP7_75t_L g1469 ( 
.A1(n_1464),
.A2(n_1440),
.B(n_1253),
.C(n_1256),
.Y(n_1469)
);

O2A1O1Ixp33_ASAP7_75t_L g1470 ( 
.A1(n_1461),
.A2(n_1445),
.B(n_1440),
.C(n_1290),
.Y(n_1470)
);

AOI221x1_ASAP7_75t_L g1471 ( 
.A1(n_1466),
.A2(n_1465),
.B1(n_1462),
.B2(n_1267),
.C(n_1384),
.Y(n_1471)
);

OAI221xp5_ASAP7_75t_L g1472 ( 
.A1(n_1466),
.A2(n_1358),
.B1(n_1326),
.B2(n_1347),
.C(n_1384),
.Y(n_1472)
);

A2O1A1Ixp33_ASAP7_75t_L g1473 ( 
.A1(n_1460),
.A2(n_1316),
.B(n_1386),
.C(n_1383),
.Y(n_1473)
);

NOR3x1_ASAP7_75t_L g1474 ( 
.A(n_1464),
.B(n_1254),
.C(n_1360),
.Y(n_1474)
);

AOI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1460),
.A2(n_1316),
.B(n_1386),
.Y(n_1475)
);

NOR2x1_ASAP7_75t_L g1476 ( 
.A(n_1467),
.B(n_1468),
.Y(n_1476)
);

AOI221x1_ASAP7_75t_L g1477 ( 
.A1(n_1475),
.A2(n_1267),
.B1(n_1375),
.B2(n_1378),
.C(n_1365),
.Y(n_1477)
);

OAI211xp5_ASAP7_75t_SL g1478 ( 
.A1(n_1470),
.A2(n_1347),
.B(n_1375),
.C(n_1366),
.Y(n_1478)
);

OAI211xp5_ASAP7_75t_SL g1479 ( 
.A1(n_1473),
.A2(n_1366),
.B(n_1282),
.C(n_1274),
.Y(n_1479)
);

INVx1_ASAP7_75t_SL g1480 ( 
.A(n_1471),
.Y(n_1480)
);

OAI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1469),
.A2(n_1334),
.B(n_1348),
.Y(n_1481)
);

AND4x1_ASAP7_75t_L g1482 ( 
.A(n_1474),
.B(n_1373),
.C(n_1380),
.D(n_1367),
.Y(n_1482)
);

OAI211xp5_ASAP7_75t_SL g1483 ( 
.A1(n_1472),
.A2(n_248),
.B(n_249),
.C(n_250),
.Y(n_1483)
);

XOR2x2_ASAP7_75t_L g1484 ( 
.A(n_1476),
.B(n_251),
.Y(n_1484)
);

NOR2x1_ASAP7_75t_L g1485 ( 
.A(n_1480),
.B(n_1483),
.Y(n_1485)
);

XOR2xp5_ASAP7_75t_L g1486 ( 
.A(n_1481),
.B(n_252),
.Y(n_1486)
);

AOI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1479),
.A2(n_1373),
.B1(n_1348),
.B2(n_1382),
.Y(n_1487)
);

AO22x1_ASAP7_75t_L g1488 ( 
.A1(n_1478),
.A2(n_1348),
.B1(n_1382),
.B2(n_1367),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1482),
.Y(n_1489)
);

NAND4xp75_ASAP7_75t_L g1490 ( 
.A(n_1477),
.B(n_254),
.C(n_256),
.D(n_257),
.Y(n_1490)
);

NOR2x1p5_ASAP7_75t_L g1491 ( 
.A(n_1476),
.B(n_261),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1485),
.B(n_262),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1491),
.B(n_263),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_SL g1494 ( 
.A(n_1484),
.B(n_1199),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1489),
.B(n_265),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_R g1496 ( 
.A(n_1486),
.B(n_269),
.Y(n_1496)
);

NOR3xp33_ASAP7_75t_SL g1497 ( 
.A(n_1490),
.B(n_270),
.C(n_276),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_R g1498 ( 
.A(n_1488),
.B(n_277),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1487),
.B(n_278),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1493),
.B(n_279),
.Y(n_1500)
);

O2A1O1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1492),
.A2(n_280),
.B(n_281),
.C(n_286),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1495),
.B(n_287),
.Y(n_1502)
);

AOI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1494),
.A2(n_1199),
.B1(n_290),
.B2(n_291),
.Y(n_1503)
);

AO22x1_ASAP7_75t_L g1504 ( 
.A1(n_1499),
.A2(n_289),
.B1(n_292),
.B2(n_296),
.Y(n_1504)
);

OAI22xp33_ASAP7_75t_R g1505 ( 
.A1(n_1496),
.A2(n_297),
.B1(n_298),
.B2(n_300),
.Y(n_1505)
);

AND2x2_ASAP7_75t_SL g1506 ( 
.A(n_1497),
.B(n_301),
.Y(n_1506)
);

AOI211xp5_ASAP7_75t_L g1507 ( 
.A1(n_1498),
.A2(n_302),
.B(n_305),
.C(n_308),
.Y(n_1507)
);

AOI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1505),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1506),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1507),
.B(n_1504),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1502),
.A2(n_313),
.B1(n_315),
.B2(n_316),
.Y(n_1511)
);

XNOR2xp5_ASAP7_75t_L g1512 ( 
.A(n_1500),
.B(n_318),
.Y(n_1512)
);

AOI22x1_ASAP7_75t_SL g1513 ( 
.A1(n_1501),
.A2(n_319),
.B1(n_320),
.B2(n_324),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1503),
.B(n_325),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1509),
.Y(n_1515)
);

NAND3xp33_ASAP7_75t_SL g1516 ( 
.A(n_1508),
.B(n_329),
.C(n_330),
.Y(n_1516)
);

AOI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1510),
.A2(n_331),
.B(n_334),
.Y(n_1517)
);

AOI22x1_ASAP7_75t_SL g1518 ( 
.A1(n_1513),
.A2(n_1512),
.B1(n_1514),
.B2(n_1511),
.Y(n_1518)
);

AOI31xp33_ASAP7_75t_L g1519 ( 
.A1(n_1515),
.A2(n_335),
.A3(n_339),
.B(n_340),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1517),
.A2(n_1518),
.B1(n_1516),
.B2(n_344),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1519),
.B(n_342),
.Y(n_1521)
);

AOI221x1_ASAP7_75t_L g1522 ( 
.A1(n_1520),
.A2(n_343),
.B1(n_347),
.B2(n_348),
.C(n_349),
.Y(n_1522)
);

AOI221xp5_ASAP7_75t_L g1523 ( 
.A1(n_1521),
.A2(n_383),
.B1(n_353),
.B2(n_355),
.C(n_359),
.Y(n_1523)
);

AOI31xp33_ASAP7_75t_L g1524 ( 
.A1(n_1522),
.A2(n_351),
.A3(n_361),
.B(n_365),
.Y(n_1524)
);

XNOR2xp5_ASAP7_75t_L g1525 ( 
.A(n_1521),
.B(n_366),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1525),
.Y(n_1526)
);

INVx4_ASAP7_75t_L g1527 ( 
.A(n_1524),
.Y(n_1527)
);

AOI221xp5_ASAP7_75t_L g1528 ( 
.A1(n_1527),
.A2(n_1523),
.B1(n_368),
.B2(n_369),
.C(n_370),
.Y(n_1528)
);

AOI211xp5_ASAP7_75t_L g1529 ( 
.A1(n_1528),
.A2(n_1526),
.B(n_371),
.C(n_372),
.Y(n_1529)
);


endmodule