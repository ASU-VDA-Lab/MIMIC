module fake_ibex_509_n_18 (n_4, n_2, n_5, n_6, n_0, n_3, n_1, n_18);

input n_4;
input n_2;
input n_5;
input n_6;
input n_0;
input n_3;
input n_1;

output n_18;

wire n_13;
wire n_7;
wire n_11;
wire n_15;
wire n_8;
wire n_17;
wire n_14;
wire n_10;
wire n_9;
wire n_16;
wire n_12;

OR2x6_ASAP7_75t_L g7 ( 
.A(n_3),
.B(n_5),
.Y(n_7)
);

OAI21xp33_ASAP7_75t_L g8 ( 
.A1(n_3),
.A2(n_4),
.B(n_1),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_1),
.B(n_6),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

OA21x2_ASAP7_75t_L g12 ( 
.A1(n_11),
.A2(n_0),
.B(n_2),
.Y(n_12)
);

AOI22xp33_ASAP7_75t_L g13 ( 
.A1(n_12),
.A2(n_11),
.B1(n_9),
.B2(n_7),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_13),
.B(n_9),
.Y(n_14)
);

OAI211xp5_ASAP7_75t_SL g15 ( 
.A1(n_14),
.A2(n_8),
.B(n_10),
.C(n_7),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_15),
.B(n_7),
.Y(n_16)
);

OAI221xp5_ASAP7_75t_L g17 ( 
.A1(n_15),
.A2(n_7),
.B1(n_12),
.B2(n_0),
.C(n_6),
.Y(n_17)
);

AO22x1_ASAP7_75t_L g18 ( 
.A1(n_16),
.A2(n_2),
.B1(n_5),
.B2(n_17),
.Y(n_18)
);


endmodule