module fake_jpeg_7621_n_295 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_43),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_25),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_45),
.B1(n_26),
.B2(n_35),
.Y(n_56)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_25),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_47),
.B(n_51),
.Y(n_83)
);

CKINVDCx6p67_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_48),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_25),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_61),
.C(n_20),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_22),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_53),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_22),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_62),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_36),
.B1(n_34),
.B2(n_19),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_59),
.B(n_60),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_31),
.B1(n_26),
.B2(n_18),
.Y(n_73)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVxp67_ASAP7_75t_SL g97 ( 
.A(n_58),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_27),
.B1(n_29),
.B2(n_36),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_27),
.B1(n_29),
.B2(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_27),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_18),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_18),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_34),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_39),
.A2(n_28),
.B(n_19),
.C(n_33),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_28),
.B(n_33),
.C(n_32),
.Y(n_84)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_17),
.Y(n_95)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_44),
.B1(n_42),
.B2(n_29),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_71),
.A2(n_73),
.B1(n_88),
.B2(n_67),
.Y(n_128)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_72),
.B(n_75),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_36),
.B1(n_34),
.B2(n_31),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_77),
.B(n_90),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_44),
.B1(n_34),
.B2(n_31),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_79),
.A2(n_67),
.B1(n_46),
.B2(n_57),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_81),
.Y(n_118)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_85),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_84),
.B(n_100),
.Y(n_109)
);

NOR3xp33_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_32),
.C(n_30),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_L g86 ( 
.A1(n_50),
.A2(n_15),
.B(n_16),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_86),
.A2(n_98),
.B1(n_107),
.B2(n_67),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_46),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_93),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_56),
.A2(n_44),
.B1(n_43),
.B2(n_26),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_89),
.Y(n_123)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_92),
.B(n_96),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_46),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_64),
.A2(n_21),
.B1(n_20),
.B2(n_43),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_61),
.A2(n_43),
.B(n_23),
.Y(n_99)
);

NOR3xp33_ASAP7_75t_SL g110 ( 
.A(n_99),
.B(n_23),
.C(n_24),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_49),
.B(n_21),
.Y(n_100)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_102),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_49),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_103),
.B(n_0),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_0),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_108),
.Y(n_120)
);

O2A1O1Ixp33_ASAP7_75t_SL g107 ( 
.A1(n_68),
.A2(n_38),
.B(n_23),
.C(n_17),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_69),
.B(n_38),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_110),
.A2(n_129),
.B(n_133),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_108),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_121),
.Y(n_145)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_24),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_130),
.Y(n_139)
);

HAxp5_ASAP7_75t_SL g152 ( 
.A(n_125),
.B(n_80),
.CON(n_152),
.SN(n_152)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_126),
.Y(n_150)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_132),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_128),
.A2(n_138),
.B1(n_70),
.B2(n_89),
.Y(n_161)
);

NOR2x1_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_66),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_90),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_66),
.Y(n_132)
);

AOI32xp33_ASAP7_75t_L g134 ( 
.A1(n_76),
.A2(n_30),
.A3(n_23),
.B1(n_58),
.B2(n_6),
.Y(n_134)
);

XNOR2x1_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_104),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_137),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_L g138 ( 
.A1(n_103),
.A2(n_58),
.B1(n_23),
.B2(n_30),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_128),
.A2(n_76),
.B1(n_80),
.B2(n_88),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_142),
.A2(n_158),
.B1(n_161),
.B2(n_162),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_130),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_144),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_109),
.B(n_83),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_109),
.B(n_83),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_149),
.Y(n_171)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_148),
.Y(n_177)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_78),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_155),
.Y(n_185)
);

AO21x1_ASAP7_75t_L g184 ( 
.A1(n_152),
.A2(n_116),
.B(n_91),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_121),
.A2(n_78),
.B1(n_99),
.B2(n_71),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_153),
.A2(n_139),
.B1(n_149),
.B2(n_142),
.Y(n_187)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_77),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_157),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_72),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_125),
.A2(n_129),
.B1(n_110),
.B2(n_112),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_118),
.B(n_104),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_133),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_163),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_93),
.B1(n_87),
.B2(n_101),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_164),
.B(n_166),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_81),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_165),
.B(n_106),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_112),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_117),
.A2(n_82),
.B1(n_107),
.B2(n_105),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_168),
.B1(n_106),
.B2(n_105),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_117),
.A2(n_122),
.B1(n_111),
.B2(n_113),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_169),
.Y(n_213)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_175),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_153),
.A2(n_134),
.B1(n_123),
.B2(n_131),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_173),
.A2(n_192),
.B1(n_150),
.B2(n_161),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_154),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_176),
.Y(n_212)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_143),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_181),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_166),
.B(n_118),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_182),
.B(n_183),
.Y(n_214)
);

AOI322xp5_ASAP7_75t_L g183 ( 
.A1(n_159),
.A2(n_116),
.A3(n_107),
.B1(n_131),
.B2(n_97),
.C1(n_58),
.C2(n_136),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_184),
.A2(n_190),
.B(n_196),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_187),
.A2(n_150),
.B1(n_140),
.B2(n_137),
.Y(n_220)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_188),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_189),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_144),
.B(n_13),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_139),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_193),
.A2(n_160),
.B1(n_147),
.B2(n_164),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_194),
.Y(n_197)
);

AOI322xp5_ASAP7_75t_SL g195 ( 
.A1(n_168),
.A2(n_12),
.A3(n_4),
.B1(n_5),
.B2(n_7),
.C1(n_9),
.C2(n_10),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_146),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_141),
.A2(n_136),
.B(n_137),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_156),
.C(n_157),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_201),
.C(n_202),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_158),
.C(n_141),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_155),
.C(n_151),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_177),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_206),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_172),
.A2(n_167),
.B(n_148),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_204),
.A2(n_208),
.B1(n_209),
.B2(n_181),
.Y(n_225)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_215),
.Y(n_224)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_178),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_209),
.B(n_211),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_171),
.B(n_170),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_190),
.C(n_194),
.Y(n_235)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_191),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_177),
.Y(n_217)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_218),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_220),
.A2(n_185),
.B1(n_183),
.B2(n_182),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_206),
.A2(n_179),
.B1(n_175),
.B2(n_186),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_221),
.A2(n_226),
.B1(n_233),
.B2(n_199),
.Y(n_250)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_225),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_211),
.A2(n_186),
.B1(n_176),
.B2(n_196),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_204),
.A2(n_192),
.B1(n_174),
.B2(n_171),
.Y(n_227)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_227),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_173),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_236),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_229),
.A2(n_232),
.B1(n_230),
.B2(n_200),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_220),
.A2(n_170),
.B1(n_184),
.B2(n_180),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_215),
.A2(n_184),
.B1(n_188),
.B2(n_185),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_237),
.C(n_205),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_198),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_58),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_140),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_239),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_9),
.Y(n_239)
);

NOR3xp33_ASAP7_75t_SL g240 ( 
.A(n_234),
.B(n_207),
.C(n_224),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_252),
.Y(n_261)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_248),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_243),
.A2(n_245),
.B1(n_229),
.B2(n_235),
.Y(n_256)
);

OA21x2_ASAP7_75t_L g244 ( 
.A1(n_226),
.A2(n_216),
.B(n_205),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_244),
.A2(n_231),
.B(n_236),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_232),
.A2(n_212),
.B1(n_197),
.B2(n_213),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_1),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_202),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_1),
.C(n_4),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_221),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_237),
.B(n_199),
.Y(n_249)
);

XNOR2x1_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_228),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_250),
.A2(n_219),
.B1(n_197),
.B2(n_238),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_233),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_239),
.Y(n_253)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_253),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_256),
.B(n_259),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_265),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_222),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_258),
.A2(n_244),
.B(n_246),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_245),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_264),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_262),
.A2(n_258),
.B(n_257),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_255),
.A2(n_249),
.B1(n_244),
.B2(n_243),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_254),
.C(n_251),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_268),
.A2(n_269),
.B(n_270),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_260),
.A2(n_240),
.B(n_247),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_254),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_272),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_266),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_274),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_263),
.Y(n_278)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_278),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_275),
.A2(n_262),
.B1(n_265),
.B2(n_251),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_279),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_268),
.A2(n_267),
.B1(n_7),
.B2(n_12),
.Y(n_281)
);

A2O1A1Ixp33_ASAP7_75t_L g288 ( 
.A1(n_281),
.A2(n_282),
.B(n_15),
.C(n_279),
.Y(n_288)
);

OAI221xp5_ASAP7_75t_L g282 ( 
.A1(n_274),
.A2(n_5),
.B1(n_7),
.B2(n_13),
.C(n_14),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_280),
.A2(n_276),
.B(n_14),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_288),
.Y(n_291)
);

MAJx2_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_5),
.C(n_14),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_281),
.C(n_283),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_285),
.C(n_15),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_287),
.Y(n_290)
);

BUFx24_ASAP7_75t_SL g293 ( 
.A(n_290),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_292),
.B(n_291),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_293),
.Y(n_295)
);


endmodule