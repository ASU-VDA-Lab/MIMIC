module real_jpeg_4348_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_2),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_2),
.A2(n_44),
.B1(n_76),
.B2(n_81),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_2),
.A2(n_44),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_2),
.A2(n_44),
.B1(n_207),
.B2(n_209),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_3),
.A2(n_50),
.B1(n_55),
.B2(n_56),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_3),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_3),
.A2(n_55),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_3),
.A2(n_25),
.B1(n_55),
.B2(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_3),
.B(n_132),
.Y(n_231)
);

O2A1O1Ixp33_ASAP7_75t_L g254 ( 
.A1(n_3),
.A2(n_255),
.B(n_257),
.C(n_263),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_3),
.B(n_22),
.C(n_64),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_3),
.B(n_86),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_3),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_3),
.B(n_67),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_4),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_4),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_4),
.A2(n_141),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_4),
.A2(n_141),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_4),
.A2(n_141),
.B1(n_292),
.B2(n_294),
.Y(n_291)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_5),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_6),
.Y(n_309)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_7),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_7),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_7),
.Y(n_133)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_7),
.Y(n_162)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_8),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_9),
.Y(n_116)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_9),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_9),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_9),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_9),
.Y(n_140)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_9),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_9),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_9),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_10),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_10),
.A2(n_21),
.B1(n_188),
.B2(n_190),
.Y(n_187)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_11),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_222),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_220),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_194),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_16),
.B(n_194),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_147),
.C(n_175),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_17),
.B(n_175),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_84),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_18),
.B(n_113),
.C(n_145),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_47),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_19),
.B(n_47),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_30),
.B(n_36),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_20),
.A2(n_153),
.B(n_155),
.Y(n_152)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_23),
.Y(n_295)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx4_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_29),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_31),
.B(n_40),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_31),
.A2(n_180),
.B(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_31),
.B(n_180),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_31),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_34),
.Y(n_178)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_36),
.B(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_36),
.B(n_290),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_39),
.Y(n_154)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_39),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g315 ( 
.A(n_46),
.Y(n_315)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_74),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_48),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_58),
.Y(n_48)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_49),
.Y(n_247)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_54),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_55),
.B(n_143),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_55),
.A2(n_165),
.B(n_203),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_L g257 ( 
.A1(n_55),
.A2(n_258),
.B(n_260),
.Y(n_257)
);

INVx4_ASAP7_75t_SL g192 ( 
.A(n_56),
.Y(n_192)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_58),
.B(n_75),
.Y(n_193)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_58),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_58),
.B(n_270),
.Y(n_269)
);

NOR2x1_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_67),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_62),
.Y(n_271)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_66),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_67),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_67),
.B(n_270),
.Y(n_286)
);

AO22x1_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_70),
.Y(n_293)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_74),
.A2(n_187),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_74),
.B(n_269),
.Y(n_297)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_88),
.B1(n_91),
.B2(n_92),
.Y(n_87)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_80),
.Y(n_274)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_113),
.B1(n_145),
.B2(n_146),
.Y(n_84)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_95),
.B(n_106),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_86),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_86),
.B(n_172),
.Y(n_244)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_87),
.B(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_90),
.Y(n_259)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_95),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_95),
.B(n_106),
.Y(n_211)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_96),
.B(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_100),
.B1(n_103),
.B2(n_104),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_99),
.Y(n_256)
);

AO22x1_ASAP7_75t_SL g132 ( 
.A1(n_100),
.A2(n_133),
.B1(n_134),
.B2(n_136),
.Y(n_132)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_102),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp33_ASAP7_75t_SL g166 ( 
.A(n_105),
.B(n_133),
.Y(n_166)
);

INVxp67_ASAP7_75t_SL g170 ( 
.A(n_106),
.Y(n_170)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_111),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_138),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_120),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_132),
.Y(n_149)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_139),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_120),
.B(n_202),
.Y(n_238)
);

NOR2x1_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_132),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_127),
.B2(n_130),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_132),
.B(n_202),
.Y(n_201)
);

INVx6_ASAP7_75t_SL g134 ( 
.A(n_135),
.Y(n_134)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_138),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_147),
.B(n_353),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.C(n_167),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_148),
.B(n_167),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_150),
.B(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_151),
.B(n_350),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_156),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_152),
.B(n_156),
.Y(n_235)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

AOI32xp33_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_160),
.A3(n_163),
.B1(n_164),
.B2(n_166),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVxp33_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_171),
.B(n_205),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_185),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_185),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_184),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_177),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_178),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_184),
.B(n_306),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B(n_193),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_186),
.A2(n_217),
.B(n_247),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_186),
.B(n_247),
.Y(n_268)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_193),
.B(n_286),
.Y(n_330)
);

BUFx24_ASAP7_75t_SL g359 ( 
.A(n_194),
.Y(n_359)
);

FAx1_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_212),
.CI(n_219),
.CON(n_194),
.SN(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_204),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_211),
.Y(n_204)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_206),
.Y(n_243)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_210),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_211),
.B(n_244),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_215),
.B1(n_216),
.B2(n_218),
.Y(n_212)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_213),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_213),
.A2(n_218),
.B1(n_254),
.B2(n_333),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_342),
.B(n_355),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_275),
.B(n_341),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_249),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_225),
.B(n_249),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_236),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_234),
.B2(n_235),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_228),
.B(n_234),
.C(n_236),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.C(n_232),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_251),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_232),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_233),
.B(n_307),
.Y(n_318)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_237),
.B(n_240),
.C(n_246),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_245),
.B1(n_246),
.B2(n_248),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_240),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_244),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_253),
.C(n_265),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_250),
.B(n_337),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_253),
.A2(n_265),
.B1(n_266),
.B2(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_253),
.Y(n_338)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_254),
.Y(n_333)
);

INVx8_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_262),
.Y(n_283)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_269),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_335),
.B(n_340),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_325),
.B(n_334),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_301),
.B(n_324),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_287),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_279),
.B(n_287),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_285),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_280),
.A2(n_281),
.B1(n_285),
.B2(n_304),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_285),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_296),
.Y(n_287)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_288),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_308),
.Y(n_307)
);

INVx6_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_297),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_298),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_298),
.B(n_299),
.C(n_327),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_310),
.B(n_323),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_305),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_303),
.B(n_305),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_319),
.B(n_322),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_318),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_316),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_321),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_328),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_326),
.B(n_328),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_332),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_330),
.B(n_331),
.C(n_332),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_339),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_336),
.B(n_339),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_351),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_344),
.B(n_345),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_349),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_347),
.B(n_348),
.C(n_349),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_351),
.A2(n_356),
.B(n_357),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_352),
.B(n_354),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_352),
.B(n_354),
.Y(n_357)
);


endmodule