module fake_jpeg_31252_n_411 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_411);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_411;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_292;
wire n_213;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx2_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_11),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_46),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_17),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_47),
.A2(n_40),
.B1(n_33),
.B2(n_21),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_49),
.Y(n_116)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_25),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_53),
.Y(n_94)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_58),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_60),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_25),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_65),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_15),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_29),
.B(n_14),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_72),
.Y(n_107)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

BUFx16f_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_69),
.Y(n_91)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_25),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_75),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_17),
.B(n_14),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_77),
.Y(n_110)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_78),
.B(n_80),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_27),
.B(n_12),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_35),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_25),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_81),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_82),
.Y(n_114)
);

BUFx12f_ASAP7_75t_SL g83 ( 
.A(n_19),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_26),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_76),
.A2(n_78),
.B1(n_73),
.B2(n_61),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_84),
.A2(n_86),
.B1(n_102),
.B2(n_108),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_54),
.A2(n_24),
.B1(n_32),
.B2(n_35),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_83),
.A2(n_32),
.B1(n_27),
.B2(n_34),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_SL g137 ( 
.A1(n_92),
.A2(n_113),
.B(n_126),
.C(n_127),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_93),
.B(n_119),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_96),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_63),
.A2(n_16),
.B1(n_40),
.B2(n_20),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_57),
.A2(n_34),
.B1(n_16),
.B2(n_19),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_44),
.B(n_0),
.Y(n_115)
);

OR2x2_ASAP7_75t_SL g165 ( 
.A(n_115),
.B(n_31),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_50),
.B(n_12),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_55),
.A2(n_39),
.B1(n_37),
.B2(n_41),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_123),
.B1(n_124),
.B2(n_46),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_56),
.A2(n_39),
.B1(n_41),
.B2(n_20),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_58),
.A2(n_39),
.B1(n_41),
.B2(n_33),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_62),
.B(n_26),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_125),
.B(n_41),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_74),
.A2(n_21),
.B1(n_31),
.B2(n_38),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_47),
.A2(n_38),
.B1(n_25),
.B2(n_31),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_131),
.B(n_139),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_132),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_133),
.Y(n_213)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_135),
.Y(n_177)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_138),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_26),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_146),
.Y(n_184)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

INVx11_ASAP7_75t_L g206 ( 
.A(n_141),
.Y(n_206)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_144),
.Y(n_196)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_106),
.A2(n_68),
.B1(n_71),
.B2(n_70),
.Y(n_146)
);

INVx6_ASAP7_75t_SL g147 ( 
.A(n_91),
.Y(n_147)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_147),
.Y(n_203)
);

HAxp5_ASAP7_75t_SL g148 ( 
.A(n_96),
.B(n_69),
.CON(n_148),
.SN(n_148)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_148),
.Y(n_187)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_149),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_L g150 ( 
.A1(n_128),
.A2(n_60),
.B1(n_81),
.B2(n_59),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_150),
.A2(n_156),
.B1(n_160),
.B2(n_87),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_93),
.B(n_38),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_151),
.B(n_155),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_106),
.B(n_38),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_153),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_106),
.B(n_38),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_99),
.B(n_26),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_154),
.B(n_157),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_107),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_45),
.B1(n_69),
.B2(n_49),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_26),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_100),
.Y(n_159)
);

INVx3_ASAP7_75t_SL g186 ( 
.A(n_159),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_89),
.A2(n_49),
.B1(n_48),
.B2(n_41),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_89),
.Y(n_161)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_161),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_85),
.Y(n_162)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_162),
.Y(n_211)
);

BUFx10_ASAP7_75t_L g163 ( 
.A(n_91),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_163),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_115),
.B(n_82),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_164),
.B(n_102),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_166),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_115),
.A2(n_48),
.B1(n_82),
.B2(n_10),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_166),
.A2(n_84),
.B1(n_95),
.B2(n_103),
.Y(n_191)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_100),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_85),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_169),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_92),
.B(n_98),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_109),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_170),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_98),
.B(n_0),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_174),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_95),
.A2(n_31),
.B1(n_2),
.B2(n_3),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_121),
.Y(n_173)
);

INVxp33_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_111),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_121),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_112),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_176),
.B(n_195),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_143),
.B(n_158),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_178),
.B(n_163),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_179),
.B(n_31),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_188),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_191),
.A2(n_150),
.B1(n_120),
.B2(n_161),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_163),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_152),
.B(n_104),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_200),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_153),
.B(n_126),
.Y(n_200)
);

AO22x1_ASAP7_75t_L g202 ( 
.A1(n_137),
.A2(n_126),
.B1(n_104),
.B2(n_114),
.Y(n_202)
);

AO21x1_ASAP7_75t_L g243 ( 
.A1(n_202),
.A2(n_208),
.B(n_141),
.Y(n_243)
);

AND2x6_ASAP7_75t_L g208 ( 
.A(n_137),
.B(n_148),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_158),
.B(n_112),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_211),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_214),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_162),
.B(n_126),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_173),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_200),
.A2(n_137),
.B(n_146),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_216),
.A2(n_211),
.B(n_178),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_184),
.A2(n_137),
.B(n_147),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_217),
.A2(n_220),
.B(n_240),
.Y(n_262)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_218),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_190),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_227),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_202),
.A2(n_165),
.B(n_134),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_202),
.A2(n_128),
.B1(n_120),
.B2(n_103),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_222),
.A2(n_225),
.B1(n_244),
.B2(n_246),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_223),
.A2(n_232),
.B1(n_248),
.B2(n_249),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_224),
.B(n_234),
.Y(n_258)
);

OAI21xp33_ASAP7_75t_SL g225 ( 
.A1(n_204),
.A2(n_163),
.B(n_144),
.Y(n_225)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_177),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_228),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_229),
.B(n_236),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_230),
.A2(n_201),
.B(n_192),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_136),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_233),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_184),
.A2(n_129),
.B1(n_135),
.B2(n_170),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_197),
.B(n_142),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_180),
.B(n_193),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_179),
.B(n_159),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_181),
.Y(n_237)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_167),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_239),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_176),
.B(n_149),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_184),
.A2(n_174),
.B(n_116),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_180),
.B(n_132),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_245),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_243),
.B(n_247),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_208),
.A2(n_129),
.B1(n_97),
.B2(n_117),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_193),
.B(n_133),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_188),
.A2(n_97),
.B1(n_117),
.B2(n_101),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_97),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_191),
.A2(n_101),
.B1(n_130),
.B2(n_111),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_207),
.A2(n_116),
.B1(n_97),
.B2(n_4),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_181),
.Y(n_250)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_250),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_252),
.B(n_281),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_195),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_257),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_226),
.A2(n_204),
.B1(n_187),
.B2(n_210),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_259),
.A2(n_276),
.B1(n_278),
.B2(n_223),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_260),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_218),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_266),
.Y(n_298)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_237),
.Y(n_267)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_267),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_226),
.A2(n_183),
.B1(n_189),
.B2(n_209),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_269),
.A2(n_247),
.B(n_238),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_241),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_277),
.Y(n_284)
);

FAx1_ASAP7_75t_SL g272 ( 
.A(n_221),
.B(n_203),
.CI(n_183),
.CON(n_272),
.SN(n_272)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_272),
.B(n_227),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_236),
.B(n_185),
.C(n_199),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_274),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_229),
.B(n_185),
.C(n_199),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_217),
.A2(n_209),
.B1(n_186),
.B2(n_205),
.Y(n_276)
);

OA22x2_ASAP7_75t_L g277 ( 
.A1(n_248),
.A2(n_203),
.B1(n_205),
.B2(n_190),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_222),
.A2(n_186),
.B1(n_182),
.B2(n_206),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_221),
.B(n_182),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_280),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_231),
.B(n_203),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_235),
.B(n_194),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_271),
.Y(n_282)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_282),
.Y(n_321)
);

NAND3xp33_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_235),
.C(n_233),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_286),
.B(n_304),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_239),
.Y(n_287)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_287),
.Y(n_330)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_256),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_292),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_290),
.B(n_291),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_256),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_265),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_294),
.B(n_296),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_295),
.A2(n_297),
.B1(n_255),
.B2(n_262),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_252),
.B(n_240),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_251),
.A2(n_216),
.B1(n_243),
.B2(n_232),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_265),
.B(n_243),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_300),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_264),
.B(n_244),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_302),
.B(n_303),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_264),
.B(n_246),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_253),
.Y(n_304)
);

NOR4xp25_ASAP7_75t_L g305 ( 
.A(n_275),
.B(n_220),
.C(n_249),
.D(n_219),
.Y(n_305)
);

NOR3xp33_ASAP7_75t_SL g318 ( 
.A(n_305),
.B(n_275),
.C(n_272),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_253),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_306),
.B(n_307),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_272),
.B(n_219),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_261),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_308),
.A2(n_269),
.B1(n_261),
.B2(n_263),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_310),
.B(n_292),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_311),
.A2(n_314),
.B1(n_299),
.B2(n_284),
.Y(n_341)
);

BUFx24_ASAP7_75t_SL g313 ( 
.A(n_301),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_313),
.B(n_296),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_297),
.A2(n_255),
.B1(n_262),
.B2(n_280),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_268),
.C(n_273),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_315),
.B(n_317),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_288),
.B(n_268),
.C(n_274),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_318),
.A2(n_331),
.B1(n_290),
.B2(n_307),
.Y(n_339)
);

INVxp33_ASAP7_75t_SL g320 ( 
.A(n_293),
.Y(n_320)
);

INVx13_ASAP7_75t_L g332 ( 
.A(n_320),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_285),
.B(n_260),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_324),
.B(n_325),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_285),
.B(n_279),
.C(n_259),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_300),
.B(n_254),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_326),
.B(n_327),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_302),
.B(n_251),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_284),
.A2(n_276),
.B1(n_278),
.B2(n_277),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_329),
.A2(n_295),
.B1(n_327),
.B2(n_291),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_301),
.A2(n_277),
.B1(n_267),
.B2(n_263),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_334),
.B(n_337),
.Y(n_352)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_309),
.Y(n_335)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_335),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_321),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_309),
.Y(n_338)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_338),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_339),
.A2(n_330),
.B1(n_289),
.B2(n_324),
.Y(n_357)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_329),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_340),
.B(n_346),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_341),
.A2(n_335),
.B1(n_338),
.B2(n_319),
.Y(n_353)
);

NOR2xp67_ASAP7_75t_L g342 ( 
.A(n_322),
.B(n_287),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_342),
.B(n_347),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_315),
.B(n_294),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_344),
.B(n_317),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_345),
.A2(n_349),
.B1(n_350),
.B2(n_298),
.Y(n_365)
);

BUFx12_ASAP7_75t_L g346 ( 
.A(n_318),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_316),
.A2(n_305),
.B(n_303),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_328),
.Y(n_348)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_348),
.Y(n_361)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_312),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_353),
.A2(n_355),
.B1(n_357),
.B2(n_345),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_354),
.B(n_344),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_341),
.A2(n_323),
.B1(n_330),
.B2(n_311),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_336),
.B(n_326),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_356),
.B(n_364),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_336),
.B(n_325),
.C(n_314),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_358),
.B(n_333),
.C(n_343),
.Y(n_373)
);

BUFx24_ASAP7_75t_SL g362 ( 
.A(n_348),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_362),
.B(n_365),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_350),
.A2(n_321),
.B(n_308),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_347),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_366),
.B(n_332),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_360),
.B(n_346),
.Y(n_368)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_368),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_363),
.A2(n_343),
.B1(n_306),
.B2(n_304),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_369),
.B(n_356),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_371),
.A2(n_370),
.B1(n_375),
.B2(n_364),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_372),
.B(n_375),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_373),
.B(n_378),
.C(n_354),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_361),
.A2(n_333),
.B1(n_283),
.B2(n_298),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_282),
.Y(n_387)
);

AO21x1_ASAP7_75t_L g375 ( 
.A1(n_351),
.A2(n_346),
.B(n_332),
.Y(n_375)
);

NOR3xp33_ASAP7_75t_L g376 ( 
.A(n_352),
.B(n_277),
.C(n_283),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_376),
.B(n_353),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_377),
.A2(n_250),
.B(n_213),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_358),
.B(n_282),
.C(n_271),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_374),
.B(n_355),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_379),
.A2(n_380),
.B(n_389),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_367),
.B(n_359),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_382),
.B(n_383),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_385),
.B(n_373),
.C(n_372),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_386),
.A2(n_387),
.B1(n_1),
.B2(n_2),
.Y(n_397)
);

NOR2xp67_ASAP7_75t_SL g388 ( 
.A(n_378),
.B(n_213),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_388),
.A2(n_206),
.B(n_196),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_390),
.B(n_392),
.C(n_396),
.Y(n_404)
);

AOI21xp33_ASAP7_75t_L g391 ( 
.A1(n_384),
.A2(n_386),
.B(n_380),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_391),
.A2(n_394),
.B(n_6),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_381),
.B(n_370),
.C(n_228),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_393),
.B(n_397),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_379),
.A2(n_196),
.B(n_186),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_385),
.B(n_196),
.C(n_2),
.Y(n_396)
);

AOI322xp5_ASAP7_75t_L g399 ( 
.A1(n_395),
.A2(n_1),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_399),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_395),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_400)
);

CKINVDCx14_ASAP7_75t_R g407 ( 
.A(n_400),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_398),
.B(n_6),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_401),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_406),
.A2(n_404),
.B(n_403),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_408),
.B(n_409),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_405),
.A2(n_402),
.B(n_407),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_410),
.B(n_7),
.Y(n_411)
);


endmodule