module real_jpeg_17349_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_524),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_0),
.B(n_525),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_1),
.A2(n_70),
.B1(n_72),
.B2(n_77),
.Y(n_69)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_1),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_1),
.A2(n_77),
.B1(n_174),
.B2(n_177),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_1),
.A2(n_77),
.B1(n_236),
.B2(n_239),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_1),
.A2(n_77),
.B1(n_348),
.B2(n_351),
.Y(n_347)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_2),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_2),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_2),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g390 ( 
.A(n_2),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_3),
.Y(n_127)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_3),
.Y(n_327)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_4),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_4),
.Y(n_225)
);

BUFx5_ASAP7_75t_L g423 ( 
.A(n_4),
.Y(n_423)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_5),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_5),
.A2(n_22),
.B1(n_107),
.B2(n_110),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_5),
.B(n_143),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_5),
.A2(n_22),
.B1(n_226),
.B2(n_231),
.Y(n_230)
);

OAI32xp33_ASAP7_75t_L g374 ( 
.A1(n_5),
.A2(n_375),
.A3(n_378),
.B1(n_379),
.B2(n_384),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_5),
.B(n_125),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_5),
.B(n_421),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_5),
.B(n_253),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_6),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_6),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_6),
.Y(n_109)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_6),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_6),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_6),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_6),
.Y(n_213)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_6),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_7),
.A2(n_45),
.B1(n_49),
.B2(n_50),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_7),
.A2(n_49),
.B1(n_118),
.B2(n_122),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_7),
.A2(n_49),
.B1(n_206),
.B2(n_210),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_7),
.B(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_8),
.A2(n_268),
.B1(n_271),
.B2(n_272),
.Y(n_267)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_8),
.Y(n_271)
);

OAI22x1_ASAP7_75t_L g294 ( 
.A1(n_8),
.A2(n_271),
.B1(n_295),
.B2(n_298),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_8),
.A2(n_271),
.B1(n_337),
.B2(n_338),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_L g400 ( 
.A1(n_8),
.A2(n_271),
.B1(n_401),
.B2(n_404),
.Y(n_400)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_9),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_12),
.Y(n_86)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_12),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_12),
.Y(n_260)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx8_ASAP7_75t_L g76 ( 
.A(n_13),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_13),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_158),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_157),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_64),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_19),
.B(n_64),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_42),
.Y(n_19)
);

NAND2xp33_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_30),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_21),
.B(n_53),
.Y(n_168)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_21),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B(n_27),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_22),
.B(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_22),
.B(n_31),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_22),
.B(n_174),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_22),
.B(n_380),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_27),
.A2(n_317),
.B1(n_354),
.B2(n_355),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_30),
.B(n_44),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_30),
.B(n_267),
.Y(n_364)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AND2x4_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_54),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_31),
.A2(n_150),
.B1(n_246),
.B2(n_266),
.Y(n_265)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_33),
.Y(n_136)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_33),
.Y(n_144)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_34),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_34),
.Y(n_139)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_34),
.Y(n_176)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_37),
.Y(n_361)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_39),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_40),
.Y(n_123)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_41),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g180 ( 
.A(n_41),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_SL g67 ( 
.A1(n_42),
.A2(n_68),
.B(n_69),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_43),
.B(n_364),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_53),
.Y(n_43)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_SL g305 ( 
.A1(n_49),
.A2(n_256),
.B(n_306),
.C(n_308),
.Y(n_305)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_52),
.Y(n_272)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_53),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_53),
.B(n_267),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_58),
.B1(n_61),
.B2(n_63),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_57),
.Y(n_357)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_148),
.C(n_152),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_65),
.B(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_78),
.C(n_115),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_66),
.A2(n_67),
.B1(n_163),
.B2(n_166),
.Y(n_162)
);

INVxp33_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_68),
.A2(n_150),
.B(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_69),
.A2(n_150),
.B(n_151),
.Y(n_149)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_78),
.A2(n_115),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_78),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_78),
.B(n_171),
.C(n_172),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_78),
.A2(n_165),
.B1(n_172),
.B2(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_78),
.A2(n_165),
.B1(n_366),
.B2(n_367),
.Y(n_365)
);

OA21x2_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_92),
.B(n_106),
.Y(n_78)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_79),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_79),
.B(n_205),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_79),
.B(n_336),
.Y(n_392)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_85),
.B1(n_87),
.B2(n_91),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_86),
.Y(n_232)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_86),
.Y(n_383)
);

INVx5_ASAP7_75t_L g403 ( 
.A(n_86),
.Y(n_403)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_89),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_90),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_92),
.B(n_205),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_92),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_92),
.B(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_92),
.B(n_106),
.Y(n_393)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_96),
.B1(n_99),
.B2(n_103),
.Y(n_93)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_94),
.Y(n_339)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_95),
.Y(n_238)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_103),
.Y(n_337)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_104),
.Y(n_377)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_106),
.Y(n_202)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_113),
.Y(n_241)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_140),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_116),
.B(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_124),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_117),
.B(n_125),
.Y(n_181)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_123),
.Y(n_297)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_123),
.Y(n_300)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_124),
.B(n_294),
.Y(n_293)
);

NOR2x1p5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_133),
.Y(n_124)
);

NAND2xp33_ASAP7_75t_SL g140 ( 
.A(n_125),
.B(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_125),
.A2(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_125),
.B(n_294),
.Y(n_368)
);

AO22x2_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_128),
.B1(n_130),
.B2(n_131),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_131),
.A2(n_134),
.B1(n_137),
.B2(n_138),
.Y(n_133)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_140),
.B(n_293),
.Y(n_463)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI32xp33_ASAP7_75t_L g315 ( 
.A1(n_145),
.A2(n_316),
.A3(n_319),
.B1(n_322),
.B2(n_328),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_149),
.A2(n_152),
.B1(n_153),
.B2(n_184),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_149),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_151),
.B(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_153),
.A2(n_476),
.B1(n_477),
.B2(n_478),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_153),
.Y(n_476)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_153),
.Y(n_497)
);

AOI21x1_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B(n_156),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_155),
.A2(n_173),
.B(n_181),
.Y(n_172)
);

NOR2x1_ASAP7_75t_L g264 ( 
.A(n_155),
.B(n_156),
.Y(n_264)
);

OAI21x1_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_185),
.B(n_522),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_182),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_161),
.B(n_182),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_167),
.C(n_169),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_162),
.A2(n_167),
.B1(n_171),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_162),
.Y(n_284)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_163),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_165),
.B(n_363),
.C(n_367),
.Y(n_485)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_167),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_167),
.A2(n_171),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_168),
.B(n_364),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_170),
.B(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_172),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_SL g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_181),
.Y(n_263)
);

NAND2xp33_ASAP7_75t_SL g292 ( 
.A(n_181),
.B(n_293),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_287),
.B(n_519),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_281),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_247),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_188),
.B(n_247),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_214),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_195),
.B2(n_196),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_191),
.Y(n_286)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_195),
.B(n_214),
.C(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

OA21x2_ASAP7_75t_L g273 ( 
.A1(n_196),
.A2(n_197),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_200),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_201),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_203),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_204),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_204),
.B(n_441),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_244),
.B(n_245),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_215),
.A2(n_216),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_233),
.Y(n_216)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_217),
.A2(n_244),
.B1(n_245),
.B2(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_217),
.B(n_315),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_217),
.A2(n_244),
.B1(n_315),
.B2(n_446),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_217),
.A2(n_233),
.B1(n_244),
.B2(n_500),
.Y(n_499)
);

OA21x2_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_221),
.B(n_229),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_218),
.A2(n_229),
.B(n_255),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_220),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_222),
.B(n_230),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_222),
.B(n_400),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_222),
.A2(n_347),
.B(n_474),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_226),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_228),
.Y(n_307)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_228),
.Y(n_419)
);

AO21x1_ASAP7_75t_L g395 ( 
.A1(n_229),
.A2(n_396),
.B(n_399),
.Y(n_395)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_233),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_242),
.B(n_243),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NAND2xp33_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_243),
.B(n_335),
.Y(n_408)
);

NAND2xp67_ASAP7_75t_L g472 ( 
.A(n_243),
.B(n_393),
.Y(n_472)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_245),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_273),
.C(n_275),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_248),
.B(n_510),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_261),
.C(n_265),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_250),
.B(n_502),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B(n_254),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_251),
.B(n_252),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_254),
.B(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_255),
.Y(n_352)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_260),
.Y(n_350)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_260),
.Y(n_406)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_262),
.B(n_265),
.Y(n_502)
);

NOR2x1_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_264),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_273),
.A2(n_276),
.B1(n_277),
.B2(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_273),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_281),
.A2(n_520),
.B(n_521),
.Y(n_519)
);

NOR2x1_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_285),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_282),
.B(n_285),
.Y(n_521)
);

AO221x1_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_457),
.B1(n_512),
.B2(n_517),
.C(n_518),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_369),
.B(n_456),
.Y(n_288)
);

NOR2xp67_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_340),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_290),
.B(n_340),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_314),
.C(n_332),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_291),
.B(n_452),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_301),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_292),
.B(n_302),
.C(n_313),
.Y(n_343)
);

INVx2_ASAP7_75t_SL g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx8_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_312),
.B2(n_313),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_304),
.B(n_425),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_305),
.B(n_399),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_305),
.Y(n_474)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

OAI21xp33_ASAP7_75t_SL g346 ( 
.A1(n_308),
.A2(n_347),
.B(n_352),
.Y(n_346)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_311),
.Y(n_398)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_314),
.A2(n_332),
.B1(n_333),
.B2(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_314),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_315),
.Y(n_446)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx6_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_320),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_321),
.Y(n_331)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_362),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_342),
.A2(n_343),
.B1(n_344),
.B2(n_345),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_342),
.B(n_345),
.C(n_362),
.Y(n_488)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_353),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_346),
.B(n_353),
.Y(n_462)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_349),
.Y(n_351)
);

INVx5_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_352),
.B(n_432),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_358),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_365),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_368),
.B(n_444),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_370),
.A2(n_450),
.B(n_455),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_371),
.A2(n_436),
.B(n_449),
.Y(n_370)
);

AOI21x1_ASAP7_75t_L g371 ( 
.A1(n_372),
.A2(n_412),
.B(n_435),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_394),
.Y(n_372)
);

NOR2xp67_ASAP7_75t_L g435 ( 
.A(n_373),
.B(n_394),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_391),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_374),
.B(n_391),
.Y(n_433)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_387),
.Y(n_384)
);

INVx5_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_393),
.Y(n_391)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_392),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_407),
.Y(n_394)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_395),
.Y(n_448)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_397),
.B(n_400),
.Y(n_425)
);

INVx4_ASAP7_75t_SL g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_408),
.A2(n_409),
.B1(n_410),
.B2(n_411),
.Y(n_407)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_408),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_409),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_409),
.B(n_410),
.C(n_448),
.Y(n_447)
);

OAI21x1_ASAP7_75t_SL g412 ( 
.A1(n_413),
.A2(n_430),
.B(n_434),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_426),
.B(n_429),
.Y(n_413)
);

NOR2x1_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_424),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_420),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_425),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_427),
.B(n_428),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_427),
.B(n_428),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_433),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_431),
.B(n_433),
.Y(n_434)
);

NOR2xp67_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_447),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_437),
.B(n_447),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_445),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_439),
.A2(n_440),
.B1(n_442),
.B2(n_443),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_439),
.B(n_443),
.C(n_445),
.Y(n_454)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVxp67_ASAP7_75t_SL g442 ( 
.A(n_443),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_451),
.B(n_454),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_451),
.B(n_454),
.Y(n_455)
);

NOR3xp33_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_491),
.C(n_505),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_459),
.B(n_487),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_459),
.B(n_515),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_479),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_460),
.B(n_479),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_467),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_461),
.B(n_468),
.C(n_493),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_463),
.C(n_464),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_482),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_463),
.A2(n_464),
.B1(n_465),
.B2(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_463),
.Y(n_483)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_470),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_470),
.Y(n_493)
);

XNOR2x1_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_475),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_471),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_473),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_472),
.B(n_473),
.Y(n_486)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_477),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_478),
.B(n_496),
.C(n_497),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_484),
.C(n_486),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_481),
.B(n_490),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_485),
.B(n_486),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_489),
.Y(n_487)
);

NOR2xp67_ASAP7_75t_L g515 ( 
.A(n_488),
.B(n_489),
.Y(n_515)
);

A2O1A1Ixp33_ASAP7_75t_L g512 ( 
.A1(n_491),
.A2(n_513),
.B(n_514),
.C(n_516),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_494),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_492),
.B(n_494),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_498),
.Y(n_494)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_495),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_499),
.A2(n_501),
.B1(n_503),
.B2(n_504),
.Y(n_498)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_499),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_499),
.B(n_507),
.C(n_508),
.Y(n_506)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_501),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_504),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_505),
.Y(n_517)
);

NOR2x1_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_509),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_506),
.B(n_509),
.Y(n_518)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);


endmodule