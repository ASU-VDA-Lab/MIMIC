module real_jpeg_27701_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_105;
wire n_40;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_18;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_278;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_97;
wire n_75;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_244;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_273;
wire n_253;
wire n_89;

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_0),
.A2(n_76),
.B1(n_77),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_0),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_0),
.A2(n_46),
.B1(n_47),
.B2(n_102),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_0),
.A2(n_27),
.B1(n_29),
.B2(n_102),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_0),
.A2(n_32),
.B1(n_35),
.B2(n_102),
.Y(n_221)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_1),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_2),
.A2(n_27),
.B1(n_29),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_2),
.A2(n_42),
.B1(n_76),
.B2(n_77),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_2),
.A2(n_32),
.B1(n_35),
.B2(n_42),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_2),
.A2(n_42),
.B1(n_46),
.B2(n_47),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_3),
.A2(n_28),
.B1(n_32),
.B2(n_35),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_3),
.A2(n_28),
.B1(n_76),
.B2(n_77),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_3),
.A2(n_28),
.B1(n_46),
.B2(n_47),
.Y(n_122)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_5),
.A2(n_46),
.B1(n_47),
.B2(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_5),
.A2(n_27),
.B1(n_29),
.B2(n_55),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_5),
.A2(n_32),
.B1(n_35),
.B2(n_55),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_7),
.A2(n_76),
.B1(n_77),
.B2(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_7),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_7),
.A2(n_46),
.B1(n_47),
.B2(n_147),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_7),
.A2(n_27),
.B1(n_29),
.B2(n_147),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_7),
.A2(n_32),
.B1(n_35),
.B2(n_147),
.Y(n_234)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_8),
.Y(n_77)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_9),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_9),
.B(n_79),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_9),
.B(n_46),
.Y(n_186)
);

AOI21xp33_ASAP7_75t_L g190 ( 
.A1(n_9),
.A2(n_46),
.B(n_186),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_9),
.A2(n_27),
.B1(n_29),
.B2(n_145),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_9),
.A2(n_32),
.B(n_36),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_9),
.B(n_95),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_9),
.A2(n_60),
.B1(n_63),
.B2(n_234),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_10),
.A2(n_27),
.B1(n_29),
.B2(n_53),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_10),
.A2(n_32),
.B1(n_35),
.B2(n_53),
.Y(n_161)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_12),
.A2(n_76),
.B1(n_77),
.B2(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_12),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_12),
.A2(n_46),
.B1(n_47),
.B2(n_127),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_12),
.A2(n_27),
.B1(n_29),
.B2(n_127),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_12),
.A2(n_32),
.B1(n_35),
.B2(n_127),
.Y(n_226)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_45)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_14),
.A2(n_27),
.B1(n_29),
.B2(n_49),
.Y(n_50)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_14),
.Y(n_185)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_15),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_129),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_128),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_105),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_20),
.B(n_105),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_85),
.B2(n_104),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_57),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_43),
.B(n_56),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_24),
.B(n_43),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_37),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_25),
.A2(n_39),
.B(n_194),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_26),
.Y(n_138)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_29),
.B1(n_34),
.B2(n_36),
.Y(n_40)
);

NAND2xp33_ASAP7_75t_SL g187 ( 
.A(n_27),
.B(n_184),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_L g212 ( 
.A1(n_27),
.A2(n_34),
.B(n_145),
.C(n_213),
.Y(n_212)
);

AOI32xp33_ASAP7_75t_L g182 ( 
.A1(n_29),
.A2(n_47),
.A3(n_183),
.B1(n_186),
.B2(n_187),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_30),
.B(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_31),
.A2(n_39),
.B1(n_68),
.B2(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_31),
.A2(n_37),
.B(n_93),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_31),
.A2(n_39),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_31),
.A2(n_39),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_31),
.A2(n_39),
.B1(n_193),
.B2(n_211),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_31),
.B(n_145),
.Y(n_232)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_32),
.Y(n_35)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_35),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_39),
.A2(n_68),
.B(n_69),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_39),
.A2(n_69),
.B(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_50),
.B1(n_51),
.B2(n_54),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_44),
.B(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_44),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_44),
.A2(n_50),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_44),
.A2(n_50),
.B1(n_141),
.B2(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_44),
.A2(n_50),
.B1(n_170),
.B2(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_50),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_47),
.B1(n_74),
.B2(n_75),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_46),
.B(n_74),
.Y(n_159)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_47),
.A2(n_78),
.B1(n_144),
.B2(n_159),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_50),
.B(n_97),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_50),
.B(n_122),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_52),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_70),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_67),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_71),
.B1(n_72),
.B2(n_84),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_59),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_59),
.A2(n_67),
.B1(n_84),
.B2(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_64),
.B(n_65),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_60),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_60),
.A2(n_63),
.B1(n_115),
.B2(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_60),
.A2(n_91),
.B(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_60),
.A2(n_226),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_61),
.A2(n_66),
.B(n_117),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_61),
.A2(n_62),
.B1(n_225),
.B2(n_227),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_66),
.Y(n_91)
);

INVx11_ASAP7_75t_L g235 ( 
.A(n_62),
.Y(n_235)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_64),
.B(n_90),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_64),
.A2(n_88),
.B(n_161),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_67),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_80),
.B(n_81),
.Y(n_72)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_73),
.A2(n_79),
.B1(n_144),
.B2(n_146),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_76),
.B(n_78),
.C(n_79),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_76),
.Y(n_78)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

HAxp5_ASAP7_75t_SL g144 ( 
.A(n_76),
.B(n_145),
.CON(n_144),
.SN(n_144)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_79),
.B(n_80),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_82),
.A2(n_100),
.B1(n_101),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_82),
.A2(n_100),
.B1(n_126),
.B2(n_152),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_85),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_94),
.C(n_98),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_87),
.B(n_92),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_94),
.A2(n_98),
.B1(n_99),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_94),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_101),
.B(n_103),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.C(n_112),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_106),
.A2(n_107),
.B1(n_110),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_110),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_112),
.B(n_277),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_119),
.C(n_124),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_113),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_118),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_119),
.A2(n_124),
.B1(n_125),
.B2(n_270),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_119),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B(n_123),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_120),
.A2(n_155),
.B(n_156),
.Y(n_154)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_274),
.B(n_279),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_174),
.B(n_260),
.C(n_273),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_162),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_132),
.B(n_162),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_148),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_134),
.B(n_135),
.C(n_148),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.C(n_143),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_136),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_143),
.B(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_145),
.B(n_240),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_146),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_157),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_153),
.B2(n_154),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_150),
.B(n_154),
.C(n_157),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_160),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.C(n_168),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_163),
.A2(n_164),
.B1(n_255),
.B2(n_257),
.Y(n_254)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_168),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.C(n_173),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_173),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_259),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_252),
.B(n_258),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_204),
.B(n_251),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_195),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_178),
.B(n_195),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_188),
.C(n_191),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_179),
.A2(n_180),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_182),
.Y(n_202)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_188),
.A2(n_189),
.B1(n_191),
.B2(n_192),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_200),
.B2(n_201),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_196),
.B(n_202),
.C(n_203),
.Y(n_253)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_245),
.B(n_250),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_222),
.B(n_244),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_214),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_207),
.B(n_214),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_212),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_208),
.A2(n_209),
.B1(n_212),
.B2(n_229),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_212),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_220),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_219),
.C(n_220),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_221),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_230),
.B(n_243),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_228),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_224),
.B(n_228),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_236),
.B(n_242),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_232),
.B(n_233),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_246),
.B(n_247),
.Y(n_250)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_253),
.B(n_254),
.Y(n_258)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_255),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_261),
.B(n_262),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_271),
.B2(n_272),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_268),
.C(n_272),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_271),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_275),
.B(n_276),
.Y(n_279)
);


endmodule