module real_aes_2301_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g586 ( .A(n_0), .B(n_187), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_1), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g145 ( .A(n_2), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_3), .B(n_548), .Y(n_547) );
NAND2xp33_ASAP7_75t_SL g629 ( .A(n_4), .B(n_174), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_5), .B(n_154), .Y(n_178) );
INVx1_ASAP7_75t_L g622 ( .A(n_6), .Y(n_622) );
INVx1_ASAP7_75t_L g200 ( .A(n_7), .Y(n_200) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_8), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_9), .Y(n_216) );
AND2x2_ASAP7_75t_L g545 ( .A(n_10), .B(n_231), .Y(n_545) );
INVx2_ASAP7_75t_L g153 ( .A(n_11), .Y(n_153) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_12), .Y(n_114) );
INVx1_ASAP7_75t_L g188 ( .A(n_13), .Y(n_188) );
AOI221x1_ASAP7_75t_L g625 ( .A1(n_14), .A2(n_205), .B1(n_550), .B2(n_626), .C(n_628), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_15), .B(n_548), .Y(n_609) );
NOR2xp33_ASAP7_75t_SL g109 ( .A(n_16), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g512 ( .A(n_16), .Y(n_512) );
INVx1_ASAP7_75t_L g185 ( .A(n_17), .Y(n_185) );
INVx1_ASAP7_75t_SL g260 ( .A(n_18), .Y(n_260) );
INVxp33_ASAP7_75t_L g837 ( .A(n_19), .Y(n_837) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_20), .B(n_165), .Y(n_164) );
AOI22xp5_ASAP7_75t_L g822 ( .A1(n_21), .A2(n_823), .B1(n_824), .B2(n_825), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_21), .Y(n_823) );
AOI33xp33_ASAP7_75t_L g237 ( .A1(n_22), .A2(n_52), .A3(n_142), .B1(n_160), .B2(n_238), .B3(n_239), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_23), .A2(n_550), .B(n_551), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_24), .B(n_187), .Y(n_552) );
AOI221xp5_ASAP7_75t_SL g596 ( .A1(n_25), .A2(n_41), .B1(n_548), .B2(n_550), .C(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g209 ( .A(n_26), .Y(n_209) );
OAI22x1_ASAP7_75t_R g503 ( .A1(n_27), .A2(n_65), .B1(n_504), .B2(n_505), .Y(n_503) );
INVx1_ASAP7_75t_L g505 ( .A(n_27), .Y(n_505) );
OA21x2_ASAP7_75t_L g152 ( .A1(n_28), .A2(n_93), .B(n_153), .Y(n_152) );
OR2x2_ASAP7_75t_L g155 ( .A(n_28), .B(n_93), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_29), .B(n_190), .Y(n_613) );
INVxp67_ASAP7_75t_L g624 ( .A(n_30), .Y(n_624) );
AND2x2_ASAP7_75t_L g571 ( .A(n_31), .B(n_230), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_32), .B(n_198), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_33), .A2(n_550), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_34), .B(n_190), .Y(n_598) );
AND2x2_ASAP7_75t_L g148 ( .A(n_35), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g159 ( .A(n_35), .Y(n_159) );
AND2x2_ASAP7_75t_L g174 ( .A(n_35), .B(n_145), .Y(n_174) );
NOR3xp33_ASAP7_75t_L g111 ( .A(n_36), .B(n_112), .C(n_114), .Y(n_111) );
OR2x6_ASAP7_75t_L g510 ( .A(n_36), .B(n_511), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_37), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_38), .B(n_198), .Y(n_224) );
AOI22xp5_ASAP7_75t_L g138 ( .A1(n_39), .A2(n_139), .B1(n_151), .B2(n_154), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_40), .B(n_171), .Y(n_170) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_42), .A2(n_83), .B1(n_157), .B2(n_550), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_43), .B(n_165), .Y(n_261) );
AOI22xp5_ASAP7_75t_SL g826 ( .A1(n_44), .A2(n_74), .B1(n_827), .B2(n_828), .Y(n_826) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_44), .Y(n_828) );
CKINVDCx20_ASAP7_75t_R g832 ( .A(n_45), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_46), .B(n_187), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_47), .B(n_176), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_48), .B(n_165), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_49), .Y(n_150) );
AND2x2_ASAP7_75t_L g589 ( .A(n_50), .B(n_230), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_51), .B(n_230), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_53), .B(n_165), .Y(n_228) );
INVx1_ASAP7_75t_L g143 ( .A(n_54), .Y(n_143) );
INVx1_ASAP7_75t_L g167 ( .A(n_54), .Y(n_167) );
XOR2x2_ASAP7_75t_L g825 ( .A(n_55), .B(n_826), .Y(n_825) );
AND2x2_ASAP7_75t_L g229 ( .A(n_56), .B(n_230), .Y(n_229) );
AOI221xp5_ASAP7_75t_L g197 ( .A1(n_57), .A2(n_76), .B1(n_157), .B2(n_198), .C(n_199), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_58), .B(n_198), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_59), .B(n_548), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_60), .B(n_151), .Y(n_218) );
AOI21xp5_ASAP7_75t_SL g248 ( .A1(n_61), .A2(n_157), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g562 ( .A(n_62), .B(n_230), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_63), .B(n_190), .Y(n_587) );
INVx1_ASAP7_75t_L g181 ( .A(n_64), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_65), .Y(n_504) );
AND2x2_ASAP7_75t_SL g614 ( .A(n_65), .B(n_231), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_66), .B(n_187), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_67), .A2(n_550), .B(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g227 ( .A(n_68), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_69), .B(n_190), .Y(n_553) );
AND2x2_ASAP7_75t_SL g578 ( .A(n_70), .B(n_176), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_71), .A2(n_157), .B(n_226), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g126 ( .A1(n_72), .A2(n_91), .B1(n_127), .B2(n_128), .Y(n_126) );
INVx1_ASAP7_75t_L g128 ( .A(n_72), .Y(n_128) );
INVx1_ASAP7_75t_L g149 ( .A(n_73), .Y(n_149) );
INVx1_ASAP7_75t_L g169 ( .A(n_73), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g827 ( .A(n_74), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_75), .B(n_198), .Y(n_240) );
AND2x2_ASAP7_75t_L g262 ( .A(n_77), .B(n_205), .Y(n_262) );
INVx1_ASAP7_75t_L g182 ( .A(n_78), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_79), .A2(n_157), .B(n_259), .Y(n_258) );
A2O1A1Ixp33_ASAP7_75t_L g156 ( .A1(n_80), .A2(n_157), .B(n_163), .C(n_175), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_81), .B(n_548), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_82), .A2(n_86), .B1(n_198), .B2(n_548), .Y(n_576) );
INVx1_ASAP7_75t_L g110 ( .A(n_84), .Y(n_110) );
AND2x2_ASAP7_75t_SL g246 ( .A(n_85), .B(n_205), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_87), .A2(n_157), .B1(n_235), .B2(n_236), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_88), .B(n_187), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_89), .B(n_187), .Y(n_599) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_90), .A2(n_125), .B1(n_126), .B2(n_129), .Y(n_124) );
INVx1_ASAP7_75t_L g129 ( .A(n_90), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_91), .Y(n_127) );
NOR3xp33_ASAP7_75t_L g526 ( .A(n_91), .B(n_132), .C(n_473), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_92), .A2(n_550), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g250 ( .A(n_94), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_95), .B(n_190), .Y(n_559) );
AND2x2_ASAP7_75t_L g241 ( .A(n_96), .B(n_205), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_97), .A2(n_207), .B(n_208), .C(n_210), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_98), .B(n_548), .Y(n_588) );
INVxp67_ASAP7_75t_L g627 ( .A(n_99), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_100), .B(n_190), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_101), .A2(n_550), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g522 ( .A(n_102), .Y(n_522) );
BUFx2_ASAP7_75t_SL g120 ( .A(n_103), .Y(n_120) );
BUFx2_ASAP7_75t_L g513 ( .A(n_103), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_104), .B(n_165), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_115), .B(n_836), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_SL g838 ( .A(n_107), .Y(n_838) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_SL g108 ( .A(n_109), .B(n_111), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_110), .B(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_114), .B(n_509), .Y(n_508) );
OR2x2_ASAP7_75t_L g521 ( .A(n_114), .B(n_510), .Y(n_521) );
AND2x6_ASAP7_75t_SL g537 ( .A(n_114), .B(n_510), .Y(n_537) );
OR2x6_ASAP7_75t_SL g821 ( .A(n_114), .B(n_509), .Y(n_821) );
AO21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_514), .B(n_831), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_121), .B(n_507), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
CKINVDCx11_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
CKINVDCx8_ASAP7_75t_R g119 ( .A(n_120), .Y(n_119) );
OAI22xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_502), .B1(n_503), .B2(n_506), .Y(n_121) );
INVx2_ASAP7_75t_L g506 ( .A(n_122), .Y(n_506) );
XNOR2x1_ASAP7_75t_L g122 ( .A(n_123), .B(n_130), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_127), .A2(n_529), .B(n_530), .Y(n_528) );
AOI21xp5_ASAP7_75t_SL g531 ( .A1(n_127), .A2(n_532), .B(n_533), .Y(n_531) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_436), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_359), .Y(n_131) );
INVxp67_ASAP7_75t_L g530 ( .A(n_132), .Y(n_530) );
NAND3xp33_ASAP7_75t_L g132 ( .A(n_133), .B(n_306), .C(n_339), .Y(n_132) );
AOI211xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_263), .B(n_272), .C(n_296), .Y(n_133) );
OAI21xp33_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_192), .B(n_242), .Y(n_134) );
OR2x2_ASAP7_75t_L g316 ( .A(n_135), .B(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g471 ( .A(n_135), .B(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AOI22xp33_ASAP7_75t_SL g361 ( .A1(n_136), .A2(n_362), .B1(n_366), .B2(n_368), .Y(n_361) );
AND2x2_ASAP7_75t_L g398 ( .A(n_136), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_177), .Y(n_136) );
INVx1_ASAP7_75t_L g295 ( .A(n_137), .Y(n_295) );
AND2x4_ASAP7_75t_L g312 ( .A(n_137), .B(n_293), .Y(n_312) );
INVx2_ASAP7_75t_L g334 ( .A(n_137), .Y(n_334) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_137), .Y(n_417) );
AND2x2_ASAP7_75t_L g488 ( .A(n_137), .B(n_245), .Y(n_488) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_156), .Y(n_137) );
NOR3xp33_ASAP7_75t_L g139 ( .A(n_140), .B(n_146), .C(n_150), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x4_ASAP7_75t_L g198 ( .A(n_141), .B(n_147), .Y(n_198) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
OR2x6_ASAP7_75t_L g172 ( .A(n_142), .B(n_161), .Y(n_172) );
INVxp33_ASAP7_75t_L g238 ( .A(n_142), .Y(n_238) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g162 ( .A(n_143), .B(n_145), .Y(n_162) );
AND2x4_ASAP7_75t_L g190 ( .A(n_143), .B(n_168), .Y(n_190) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x6_ASAP7_75t_L g550 ( .A(n_148), .B(n_162), .Y(n_550) );
INVx2_ASAP7_75t_L g161 ( .A(n_149), .Y(n_161) );
AND2x6_ASAP7_75t_L g187 ( .A(n_149), .B(n_166), .Y(n_187) );
INVx4_ASAP7_75t_L g205 ( .A(n_151), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_151), .B(n_215), .Y(n_214) );
AOI21x1_ASAP7_75t_L g582 ( .A1(n_151), .A2(n_583), .B(n_589), .Y(n_582) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx4f_ASAP7_75t_L g176 ( .A(n_152), .Y(n_176) );
AND2x4_ASAP7_75t_L g154 ( .A(n_153), .B(n_155), .Y(n_154) );
AND2x2_ASAP7_75t_SL g231 ( .A(n_153), .B(n_155), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_154), .B(n_173), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_154), .A2(n_248), .B(n_252), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_154), .A2(n_547), .B(n_549), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_154), .B(n_622), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_154), .B(n_624), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_154), .B(n_627), .Y(n_626) );
NOR3xp33_ASAP7_75t_L g628 ( .A(n_154), .B(n_183), .C(n_629), .Y(n_628) );
INVxp67_ASAP7_75t_L g217 ( .A(n_157), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_157), .A2(n_198), .B1(n_621), .B2(n_623), .Y(n_620) );
AND2x4_ASAP7_75t_L g157 ( .A(n_158), .B(n_162), .Y(n_157) );
NOR2x1p5_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
INVx1_ASAP7_75t_L g239 ( .A(n_160), .Y(n_239) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_170), .B(n_173), .Y(n_163) );
INVx1_ASAP7_75t_L g183 ( .A(n_165), .Y(n_183) );
AND2x4_ASAP7_75t_L g548 ( .A(n_165), .B(n_174), .Y(n_548) );
AND2x4_ASAP7_75t_L g165 ( .A(n_166), .B(n_168), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
OAI22xp5_ASAP7_75t_L g180 ( .A1(n_172), .A2(n_181), .B1(n_182), .B2(n_183), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_SL g199 ( .A1(n_172), .A2(n_173), .B(n_200), .C(n_201), .Y(n_199) );
INVxp67_ASAP7_75t_L g207 ( .A(n_172), .Y(n_207) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_172), .A2(n_173), .B(n_227), .C(n_228), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_172), .A2(n_173), .B(n_250), .C(n_251), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_SL g259 ( .A1(n_172), .A2(n_173), .B(n_260), .C(n_261), .Y(n_259) );
INVx1_ASAP7_75t_L g235 ( .A(n_173), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_173), .A2(n_552), .B(n_553), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_173), .A2(n_559), .B(n_560), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_173), .A2(n_568), .B(n_569), .Y(n_567) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_173), .A2(n_586), .B(n_587), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_173), .A2(n_598), .B(n_599), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_173), .A2(n_612), .B(n_613), .Y(n_611) );
INVx5_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_174), .Y(n_210) );
AO21x2_ASAP7_75t_L g232 ( .A1(n_175), .A2(n_233), .B(n_241), .Y(n_232) );
AO21x2_ASAP7_75t_L g277 ( .A1(n_175), .A2(n_233), .B(n_241), .Y(n_277) );
AOI21x1_ASAP7_75t_L g574 ( .A1(n_175), .A2(n_575), .B(n_578), .Y(n_574) );
INVx2_ASAP7_75t_SL g175 ( .A(n_176), .Y(n_175) );
OA21x2_ASAP7_75t_L g196 ( .A1(n_176), .A2(n_197), .B(n_202), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_176), .A2(n_609), .B(n_610), .Y(n_608) );
AND2x2_ASAP7_75t_L g253 ( .A(n_177), .B(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g282 ( .A(n_177), .Y(n_282) );
INVx3_ASAP7_75t_L g293 ( .A(n_177), .Y(n_293) );
AND2x4_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
OAI21xp5_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_184), .B(n_191), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_183), .B(n_209), .Y(n_208) );
OAI22xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B1(n_188), .B2(n_189), .Y(n_184) );
INVxp67_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVxp67_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_192), .A2(n_483), .B1(n_485), .B2(n_487), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_192), .B(n_494), .Y(n_493) );
INVx2_ASAP7_75t_SL g192 ( .A(n_193), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_220), .Y(n_193) );
INVx3_ASAP7_75t_L g266 ( .A(n_194), .Y(n_266) );
AND2x2_ASAP7_75t_L g274 ( .A(n_194), .B(n_275), .Y(n_274) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_194), .Y(n_304) );
NAND2x1_ASAP7_75t_SL g498 ( .A(n_194), .B(n_265), .Y(n_498) );
AND2x4_ASAP7_75t_L g194 ( .A(n_195), .B(n_203), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g271 ( .A(n_196), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_196), .B(n_277), .Y(n_289) );
AND2x2_ASAP7_75t_L g302 ( .A(n_196), .B(n_203), .Y(n_302) );
AND2x4_ASAP7_75t_L g309 ( .A(n_196), .B(n_310), .Y(n_309) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_196), .Y(n_358) );
INVxp67_ASAP7_75t_L g365 ( .A(n_196), .Y(n_365) );
INVx1_ASAP7_75t_L g370 ( .A(n_196), .Y(n_370) );
INVx1_ASAP7_75t_L g219 ( .A(n_198), .Y(n_219) );
INVx1_ASAP7_75t_L g269 ( .A(n_203), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_203), .B(n_279), .Y(n_288) );
INVx2_ASAP7_75t_L g356 ( .A(n_203), .Y(n_356) );
INVx1_ASAP7_75t_L g395 ( .A(n_203), .Y(n_395) );
OR2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_213), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B1(n_211), .B2(n_212), .Y(n_204) );
INVx3_ASAP7_75t_L g212 ( .A(n_205), .Y(n_212) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_212), .A2(n_223), .B(n_229), .Y(n_222) );
AO21x2_ASAP7_75t_L g279 ( .A1(n_212), .A2(n_223), .B(n_229), .Y(n_279) );
OAI22xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_217), .B1(n_218), .B2(n_219), .Y(n_213) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g325 ( .A(n_220), .B(n_302), .Y(n_325) );
AND2x2_ASAP7_75t_L g393 ( .A(n_220), .B(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g407 ( .A(n_220), .B(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_220), .B(n_422), .Y(n_421) );
AND2x4_ASAP7_75t_L g220 ( .A(n_221), .B(n_232), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NOR2x1_ASAP7_75t_L g270 ( .A(n_222), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g363 ( .A(n_222), .B(n_356), .Y(n_363) );
AND2x2_ASAP7_75t_L g454 ( .A(n_222), .B(n_276), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_230), .Y(n_255) );
OA21x2_ASAP7_75t_L g595 ( .A1(n_230), .A2(n_596), .B(n_600), .Y(n_595) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g265 ( .A(n_232), .Y(n_265) );
INVx2_ASAP7_75t_L g310 ( .A(n_232), .Y(n_310) );
AND2x2_ASAP7_75t_L g355 ( .A(n_232), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_234), .B(n_240), .Y(n_233) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_253), .Y(n_243) );
AND2x2_ASAP7_75t_L g397 ( .A(n_244), .B(n_398), .Y(n_397) );
OR2x6_ASAP7_75t_L g456 ( .A(n_244), .B(n_457), .Y(n_456) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx4_ASAP7_75t_L g286 ( .A(n_245), .Y(n_286) );
AND2x4_ASAP7_75t_L g294 ( .A(n_245), .B(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g329 ( .A(n_245), .B(n_254), .Y(n_329) );
INVx2_ASAP7_75t_L g378 ( .A(n_245), .Y(n_378) );
NAND2xp5_ASAP7_75t_SL g427 ( .A(n_245), .B(n_352), .Y(n_427) );
AND2x2_ASAP7_75t_L g464 ( .A(n_245), .B(n_282), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_245), .B(n_347), .Y(n_472) );
OR2x6_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
AND2x2_ASAP7_75t_L g305 ( .A(n_253), .B(n_294), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_253), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_SL g444 ( .A(n_253), .B(n_332), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_253), .B(n_345), .Y(n_466) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_254), .Y(n_284) );
AND2x2_ASAP7_75t_L g292 ( .A(n_254), .B(n_293), .Y(n_292) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_254), .Y(n_315) );
INVx2_ASAP7_75t_L g318 ( .A(n_254), .Y(n_318) );
INVx1_ASAP7_75t_L g351 ( .A(n_254), .Y(n_351) );
INVx1_ASAP7_75t_L g399 ( .A(n_254), .Y(n_399) );
AO21x2_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_256), .B(n_262), .Y(n_254) );
AO21x2_ASAP7_75t_L g555 ( .A1(n_255), .A2(n_556), .B(n_562), .Y(n_555) );
AO21x2_ASAP7_75t_L g564 ( .A1(n_255), .A2(n_565), .B(n_571), .Y(n_564) );
AO21x2_ASAP7_75t_L g603 ( .A1(n_255), .A2(n_565), .B(n_571), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
NAND2xp33_ASAP7_75t_L g263 ( .A(n_264), .B(n_267), .Y(n_263) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_265), .B(n_268), .Y(n_341) );
OR2x2_ASAP7_75t_L g413 ( .A(n_265), .B(n_414), .Y(n_413) );
AND4x1_ASAP7_75t_SL g459 ( .A(n_265), .B(n_441), .C(n_460), .D(n_461), .Y(n_459) );
OR2x2_ASAP7_75t_L g483 ( .A(n_266), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
AND2x2_ASAP7_75t_L g320 ( .A(n_269), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_269), .B(n_278), .Y(n_470) );
AND2x2_ASAP7_75t_L g495 ( .A(n_270), .B(n_355), .Y(n_495) );
OAI32xp33_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_280), .A3(n_285), .B1(n_287), .B2(n_290), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g368 ( .A(n_275), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g468 ( .A(n_275), .B(n_422), .Y(n_468) );
AND2x4_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
AND2x2_ASAP7_75t_L g364 ( .A(n_276), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g450 ( .A(n_276), .Y(n_450) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_277), .B(n_279), .Y(n_484) );
INVx3_ASAP7_75t_L g301 ( .A(n_278), .Y(n_301) );
NAND2x1p5_ASAP7_75t_L g479 ( .A(n_278), .B(n_406), .Y(n_479) );
INVx3_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_279), .Y(n_338) );
AND2x2_ASAP7_75t_L g357 ( .A(n_279), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g491 ( .A(n_281), .Y(n_491) );
NAND2x1_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx1_ASAP7_75t_L g331 ( .A(n_282), .Y(n_331) );
NOR2x1_ASAP7_75t_L g432 ( .A(n_282), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_285), .B(n_391), .Y(n_390) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g323 ( .A(n_286), .B(n_291), .Y(n_323) );
AND2x4_ASAP7_75t_L g345 ( .A(n_286), .B(n_295), .Y(n_345) );
AND2x4_ASAP7_75t_SL g416 ( .A(n_286), .B(n_417), .Y(n_416) );
NOR2x1_ASAP7_75t_L g442 ( .A(n_286), .B(n_367), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_287), .A2(n_410), .B1(n_413), .B2(n_415), .Y(n_409) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx2_ASAP7_75t_SL g429 ( .A(n_288), .Y(n_429) );
INVx2_ASAP7_75t_L g321 ( .A(n_289), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_294), .Y(n_290) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_292), .B(n_298), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_292), .A2(n_428), .B1(n_431), .B2(n_434), .Y(n_430) );
INVx1_ASAP7_75t_L g352 ( .A(n_293), .Y(n_352) );
AND2x2_ASAP7_75t_L g375 ( .A(n_293), .B(n_334), .Y(n_375) );
INVx2_ASAP7_75t_L g298 ( .A(n_294), .Y(n_298) );
OAI21xp5_ASAP7_75t_SL g296 ( .A1(n_297), .A2(n_299), .B(n_303), .Y(n_296) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_300), .A2(n_372), .B1(n_376), .B2(n_377), .Y(n_371) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_301), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_301), .B(n_369), .Y(n_385) );
INVx1_ASAP7_75t_L g389 ( .A(n_301), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
NOR3xp33_ASAP7_75t_L g306 ( .A(n_307), .B(n_322), .C(n_326), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_311), .B1(n_316), .B2(n_319), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g336 ( .A(n_309), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g376 ( .A(n_309), .B(n_363), .Y(n_376) );
AND2x2_ASAP7_75t_L g428 ( .A(n_309), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g445 ( .A(n_309), .B(n_395), .Y(n_445) );
AND2x2_ASAP7_75t_L g500 ( .A(n_309), .B(n_394), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx4_ASAP7_75t_L g367 ( .A(n_312), .Y(n_367) );
AND2x2_ASAP7_75t_L g377 ( .A(n_312), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx2_ASAP7_75t_L g382 ( .A(n_315), .Y(n_382) );
AND2x2_ASAP7_75t_L g391 ( .A(n_315), .B(n_375), .Y(n_391) );
INVx1_ASAP7_75t_L g426 ( .A(n_317), .Y(n_426) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g347 ( .A(n_318), .Y(n_347) );
INVxp67_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_320), .B(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_321), .B(n_389), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_330), .B(n_335), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_328), .B(n_367), .Y(n_476) );
INVx2_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
AOI21xp33_ASAP7_75t_SL g339 ( .A1(n_331), .A2(n_340), .B(n_342), .Y(n_339) );
AND2x2_ASAP7_75t_L g486 ( .A(n_331), .B(n_345), .Y(n_486) );
AND2x4_ASAP7_75t_L g349 ( .A(n_332), .B(n_350), .Y(n_349) );
INVx2_ASAP7_75t_SL g383 ( .A(n_332), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_332), .B(n_399), .Y(n_465) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AOI21xp33_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_348), .B(n_353), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_345), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_345), .B(n_350), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_346), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g408 ( .A(n_346), .Y(n_408) );
INVx1_ASAP7_75t_L g412 ( .A(n_346), .Y(n_412) );
AND2x2_ASAP7_75t_L g496 ( .A(n_346), .B(n_464), .Y(n_496) );
AND2x2_ASAP7_75t_L g499 ( .A(n_346), .B(n_416), .Y(n_499) );
INVx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x4_ASAP7_75t_SL g350 ( .A(n_351), .B(n_352), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_351), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_355), .B(n_357), .Y(n_354) );
INVx1_ASAP7_75t_L g478 ( .A(n_355), .Y(n_478) );
AND2x2_ASAP7_75t_L g369 ( .A(n_356), .B(n_370), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_359), .B(n_437), .Y(n_527) );
INVxp67_ASAP7_75t_L g529 ( .A(n_359), .Y(n_529) );
NAND4xp75_ASAP7_75t_L g359 ( .A(n_360), .B(n_379), .C(n_400), .D(n_418), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_371), .Y(n_360) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
NAND2x1p5_ASAP7_75t_L g449 ( .A(n_363), .B(n_450), .Y(n_449) );
NAND2x1p5_ASAP7_75t_L g435 ( .A(n_364), .B(n_429), .Y(n_435) );
NAND2xp5_ASAP7_75t_R g451 ( .A(n_367), .B(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g501 ( .A(n_367), .Y(n_501) );
INVx2_ASAP7_75t_L g414 ( .A(n_369), .Y(n_414) );
BUFx3_ASAP7_75t_L g406 ( .A(n_370), .Y(n_406) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g457 ( .A(n_375), .Y(n_457) );
AND2x2_ASAP7_75t_L g411 ( .A(n_377), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g433 ( .A(n_378), .Y(n_433) );
AOI21xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_384), .B(n_386), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_382), .B(n_416), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_383), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_385), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_390), .B1(n_392), .B2(n_396), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
OA21x2_ASAP7_75t_L g401 ( .A1(n_394), .A2(n_402), .B(n_403), .Y(n_401) );
INVx1_ASAP7_75t_L g422 ( .A(n_394), .Y(n_422) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g453 ( .A(n_395), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g461 ( .A(n_395), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_396), .B(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g431 ( .A(n_399), .B(n_432), .Y(n_431) );
AOI21xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_407), .B(n_409), .Y(n_400) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OR2x2_ASAP7_75t_L g448 ( .A(n_405), .B(n_449), .Y(n_448) );
INVx3_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_412), .Y(n_460) );
INVx2_ASAP7_75t_SL g452 ( .A(n_416), .Y(n_452) );
AND2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_430), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_423), .B1(n_425), .B2(n_428), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g481 ( .A(n_425), .Y(n_481) );
NOR2x1_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
INVx3_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_437), .B(n_473), .Y(n_436) );
INVxp67_ASAP7_75t_L g533 ( .A(n_437), .Y(n_533) );
NAND3xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_446), .C(n_458), .Y(n_437) );
NOR2x1_ASAP7_75t_L g438 ( .A(n_439), .B(n_443), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
AOI22xp33_ASAP7_75t_SL g446 ( .A1(n_447), .A2(n_451), .B1(n_453), .B2(n_455), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NOR3xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_462), .C(n_469), .Y(n_458) );
AOI21xp33_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_466), .B(n_467), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVxp67_ASAP7_75t_L g532 ( .A(n_473), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_492), .Y(n_473) );
NOR3xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_482), .C(n_489), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B1(n_480), .B2(n_481), .Y(n_475) );
OR2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
NOR3xp33_ASAP7_75t_L g489 ( .A(n_483), .B(n_488), .C(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVxp67_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AOI222xp33_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_496), .B1(n_497), .B2(n_499), .C1(n_500), .C2(n_501), .Y(n_492) );
INVx1_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NOR2x1_ASAP7_75t_R g507 ( .A(n_508), .B(n_513), .Y(n_507) );
BUFx3_ASAP7_75t_L g835 ( .A(n_508), .Y(n_835) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_510), .Y(n_509) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_513), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_523), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_516), .B(n_518), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_517), .Y(n_516) );
NOR2xp33_ASAP7_75t_SL g518 ( .A(n_519), .B(n_522), .Y(n_518) );
INVx1_ASAP7_75t_SL g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_822), .B1(n_829), .B2(n_830), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_534), .B1(n_538), .B2(n_819), .Y(n_524) );
AO22x2_ASAP7_75t_L g830 ( .A1(n_525), .A2(n_535), .B1(n_538), .B2(n_820), .Y(n_830) );
AOI211x1_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_527), .B(n_528), .C(n_531), .Y(n_525) );
INVx4_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
INVx3_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_537), .Y(n_536) );
INVx3_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_749), .Y(n_539) );
NOR4xp25_ASAP7_75t_SL g540 ( .A(n_541), .B(n_642), .C(n_686), .D(n_713), .Y(n_540) );
OAI221xp5_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_605), .B1(n_615), .B2(n_630), .C(n_632), .Y(n_541) );
AOI32xp33_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_572), .A3(n_579), .B1(n_590), .B2(n_601), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g784 ( .A(n_543), .B(n_785), .Y(n_784) );
AOI22xp5_ASAP7_75t_L g812 ( .A1(n_543), .A2(n_755), .B1(n_813), .B2(n_816), .Y(n_812) );
AND2x4_ASAP7_75t_SL g543 ( .A(n_544), .B(n_554), .Y(n_543) );
INVx5_ASAP7_75t_L g604 ( .A(n_544), .Y(n_604) );
OR2x2_ASAP7_75t_L g631 ( .A(n_544), .B(n_603), .Y(n_631) );
AND2x4_ASAP7_75t_L g633 ( .A(n_544), .B(n_564), .Y(n_633) );
INVx2_ASAP7_75t_L g648 ( .A(n_544), .Y(n_648) );
OR2x2_ASAP7_75t_L g660 ( .A(n_544), .B(n_573), .Y(n_660) );
AND2x2_ASAP7_75t_L g667 ( .A(n_544), .B(n_563), .Y(n_667) );
AND2x2_ASAP7_75t_SL g709 ( .A(n_544), .B(n_592), .Y(n_709) );
HB1xp67_ASAP7_75t_L g766 ( .A(n_544), .Y(n_766) );
OR2x6_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
INVx3_ASAP7_75t_SL g661 ( .A(n_554), .Y(n_661) );
AND2x2_ASAP7_75t_L g680 ( .A(n_554), .B(n_604), .Y(n_680) );
AOI32xp33_ASAP7_75t_L g795 ( .A1(n_554), .A2(n_666), .A3(n_696), .B1(n_726), .B2(n_761), .Y(n_795) );
AND2x4_ASAP7_75t_L g554 ( .A(n_555), .B(n_563), .Y(n_554) );
AND2x2_ASAP7_75t_L g635 ( .A(n_555), .B(n_573), .Y(n_635) );
OR2x2_ASAP7_75t_L g651 ( .A(n_555), .B(n_564), .Y(n_651) );
INVx1_ASAP7_75t_L g674 ( .A(n_555), .Y(n_674) );
INVx2_ASAP7_75t_L g690 ( .A(n_555), .Y(n_690) );
AND2x2_ASAP7_75t_L g727 ( .A(n_555), .B(n_592), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_555), .B(n_564), .Y(n_746) );
HB1xp67_ASAP7_75t_L g815 ( .A(n_555), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_561), .Y(n_556) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g782 ( .A(n_564), .B(n_573), .Y(n_782) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_564), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_570), .Y(n_565) );
OR2x2_ASAP7_75t_L g630 ( .A(n_572), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g636 ( .A(n_572), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g649 ( .A(n_572), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g811 ( .A(n_572), .B(n_680), .Y(n_811) );
BUFx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g740 ( .A(n_573), .B(n_690), .Y(n_740) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
BUFx6f_ASAP7_75t_L g592 ( .A(n_574), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g809 ( .A(n_579), .B(n_707), .Y(n_809) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_580), .B(n_757), .Y(n_756) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g594 ( .A(n_581), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g616 ( .A(n_581), .Y(n_616) );
AND2x2_ASAP7_75t_L g640 ( .A(n_581), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_581), .B(n_618), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_581), .B(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g698 ( .A(n_581), .Y(n_698) );
OR2x2_ASAP7_75t_L g717 ( .A(n_581), .B(n_644), .Y(n_717) );
INVx1_ASAP7_75t_L g724 ( .A(n_581), .Y(n_724) );
NOR2xp33_ASAP7_75t_R g776 ( .A(n_581), .B(n_607), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_581), .B(n_619), .Y(n_780) );
INVx3_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_588), .Y(n_583) );
AOI32xp33_ASAP7_75t_L g803 ( .A1(n_590), .A2(n_639), .A3(n_804), .B1(n_805), .B2(n_806), .Y(n_803) );
INVx3_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVx2_ASAP7_75t_L g670 ( .A(n_592), .Y(n_670) );
AND2x4_ASAP7_75t_L g689 ( .A(n_592), .B(n_690), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_592), .B(n_661), .Y(n_718) );
OR2x2_ASAP7_75t_L g772 ( .A(n_592), .B(n_773), .Y(n_772) );
OR2x2_ASAP7_75t_L g730 ( .A(n_593), .B(n_731), .Y(n_730) );
OR2x2_ASAP7_75t_L g788 ( .A(n_593), .B(n_789), .Y(n_788) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_594), .B(n_607), .Y(n_754) );
AND2x2_ASAP7_75t_L g791 ( .A(n_594), .B(n_757), .Y(n_791) );
INVx2_ASAP7_75t_L g641 ( .A(n_595), .Y(n_641) );
INVx2_ASAP7_75t_L g644 ( .A(n_595), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_595), .B(n_607), .Y(n_664) );
INVx1_ASAP7_75t_L g695 ( .A(n_595), .Y(n_695) );
OR2x2_ASAP7_75t_L g721 ( .A(n_595), .B(n_607), .Y(n_721) );
HB1xp67_ASAP7_75t_L g773 ( .A(n_595), .Y(n_773) );
BUFx3_ASAP7_75t_L g802 ( .A(n_595), .Y(n_802) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g671 ( .A(n_602), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_602), .B(n_689), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_602), .B(n_760), .Y(n_759) );
AND2x4_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_603), .B(n_674), .Y(n_673) );
OAI21xp33_ASAP7_75t_L g703 ( .A1(n_603), .A2(n_670), .B(n_688), .Y(n_703) );
OAI32xp33_ASAP7_75t_L g725 ( .A1(n_604), .A2(n_726), .A3(n_728), .B1(n_730), .B2(n_732), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_604), .B(n_689), .Y(n_798) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g731 ( .A(n_606), .Y(n_731) );
NOR2x1p5_ASAP7_75t_L g801 ( .A(n_606), .B(n_802), .Y(n_801) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x4_ASAP7_75t_L g617 ( .A(n_607), .B(n_618), .Y(n_617) );
AND2x4_ASAP7_75t_SL g639 ( .A(n_607), .B(n_619), .Y(n_639) );
OR2x2_ASAP7_75t_L g643 ( .A(n_607), .B(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g678 ( .A(n_607), .Y(n_678) );
AND2x2_ASAP7_75t_L g696 ( .A(n_607), .B(n_697), .Y(n_696) );
OR2x2_ASAP7_75t_L g707 ( .A(n_607), .B(n_619), .Y(n_707) );
OR2x2_ASAP7_75t_L g769 ( .A(n_607), .B(n_770), .Y(n_769) );
OR2x2_ASAP7_75t_L g786 ( .A(n_607), .B(n_717), .Y(n_786) );
INVx1_ASAP7_75t_L g818 ( .A(n_607), .Y(n_818) );
OR2x6_ASAP7_75t_L g607 ( .A(n_608), .B(n_614), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_616), .B(n_695), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_617), .B(n_729), .Y(n_728) );
AOI222xp33_ASAP7_75t_L g733 ( .A1(n_617), .A2(n_734), .B1(n_739), .B2(n_741), .C1(n_744), .C2(n_747), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_617), .B(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g761 ( .A(n_617), .B(n_640), .Y(n_761) );
AND2x2_ASAP7_75t_L g723 ( .A(n_618), .B(n_724), .Y(n_723) );
OR2x2_ASAP7_75t_L g738 ( .A(n_618), .B(n_643), .Y(n_738) );
INVx3_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_619), .B(n_644), .Y(n_676) );
AND2x4_ASAP7_75t_L g697 ( .A(n_619), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g757 ( .A(n_619), .B(n_678), .Y(n_757) );
AND2x4_ASAP7_75t_L g619 ( .A(n_620), .B(n_625), .Y(n_619) );
INVx1_ASAP7_75t_SL g637 ( .A(n_631), .Y(n_637) );
NAND2xp33_ASAP7_75t_SL g806 ( .A(n_631), .B(n_661), .Y(n_806) );
A2O1A1Ixp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B(n_636), .C(n_638), .Y(n_632) );
INVx2_ASAP7_75t_SL g683 ( .A(n_633), .Y(n_683) );
AND2x2_ASAP7_75t_L g687 ( .A(n_634), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_635), .B(n_683), .Y(n_682) );
O2A1O1Ixp33_ASAP7_75t_L g708 ( .A1(n_635), .A2(n_673), .B(n_709), .C(n_710), .Y(n_708) );
AND2x2_ASAP7_75t_L g785 ( .A(n_635), .B(n_766), .Y(n_785) );
AND2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
AND2x4_ASAP7_75t_L g684 ( .A(n_639), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_SL g789 ( .A(n_639), .Y(n_789) );
OAI211xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_645), .B(n_652), .C(n_679), .Y(n_642) );
INVx2_ASAP7_75t_L g654 ( .A(n_643), .Y(n_654) );
OR2x2_ASAP7_75t_L g701 ( .A(n_643), .B(n_702), .Y(n_701) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_644), .Y(n_685) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_649), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_647), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g739 ( .A(n_647), .B(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_647), .B(n_727), .Y(n_793) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AOI222xp33_ASAP7_75t_L g751 ( .A1(n_649), .A2(n_752), .B1(n_753), .B2(n_755), .C1(n_758), .C2(n_761), .Y(n_751) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_650), .A2(n_715), .B1(n_718), .B2(n_719), .C(n_725), .Y(n_714) );
AND2x2_ASAP7_75t_L g752 ( .A(n_650), .B(n_709), .Y(n_752) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2xp33_ASAP7_75t_SL g665 ( .A(n_651), .B(n_666), .Y(n_665) );
AOI221x1_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_657), .B1(n_662), .B2(n_665), .C(n_668), .Y(n_652) );
AND2x4_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
AND2x2_ASAP7_75t_L g805 ( .A(n_655), .B(n_743), .Y(n_805) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OR2x2_ASAP7_75t_L g663 ( .A(n_656), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_661), .Y(n_658) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
OAI32xp33_ASAP7_75t_L g771 ( .A1(n_661), .A2(n_702), .A3(n_772), .B1(n_774), .B2(n_778), .Y(n_771) );
OAI21xp33_ASAP7_75t_SL g790 ( .A1(n_662), .A2(n_791), .B(n_792), .Y(n_790) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AOI21xp33_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_672), .B(n_675), .Y(n_668) );
OR2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
OR2x2_ASAP7_75t_L g672 ( .A(n_670), .B(n_673), .Y(n_672) );
OR2x2_ASAP7_75t_L g745 ( .A(n_670), .B(n_746), .Y(n_745) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_674), .A2(n_700), .B1(n_703), .B2(n_704), .C(n_708), .Y(n_699) );
INVx1_ASAP7_75t_L g775 ( .A(n_674), .Y(n_775) );
HB1xp67_ASAP7_75t_L g781 ( .A(n_674), .Y(n_781) );
OR2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
OAI21xp33_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_681), .B(n_684), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_683), .B(n_748), .Y(n_747) );
OAI21xp5_ASAP7_75t_SL g686 ( .A1(n_687), .A2(n_691), .B(n_699), .Y(n_686) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_690), .Y(n_760) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_696), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_693), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVxp67_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g712 ( .A(n_695), .Y(n_712) );
INVx1_ASAP7_75t_L g702 ( .A(n_697), .Y(n_702) );
AND2x2_ASAP7_75t_SL g711 ( .A(n_697), .B(n_712), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_697), .B(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_697), .B(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
OR2x2_ASAP7_75t_L g716 ( .A(n_707), .B(n_717), .Y(n_716) );
INVx2_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_712), .Y(n_777) );
NAND2xp5_ASAP7_75t_SL g713 ( .A(n_714), .B(n_733), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g729 ( .A(n_717), .Y(n_729) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
OR2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
INVx1_ASAP7_75t_SL g743 ( .A(n_721), .Y(n_743) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_723), .B(n_801), .Y(n_800) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_724), .Y(n_737) );
BUFx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_SL g734 ( .A(n_735), .B(n_738), .Y(n_734) );
INVxp67_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g748 ( .A(n_740), .Y(n_748) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g767 ( .A(n_746), .Y(n_767) );
NOR4xp25_ASAP7_75t_L g749 ( .A(n_750), .B(n_783), .C(n_794), .D(n_807), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_751), .B(n_762), .Y(n_750) );
O2A1O1Ixp33_ASAP7_75t_L g762 ( .A1(n_752), .A2(n_763), .B(n_768), .C(n_771), .Y(n_762) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
NAND2xp5_ASAP7_75t_SL g764 ( .A(n_765), .B(n_767), .Y(n_764) );
OAI211xp5_ASAP7_75t_L g774 ( .A1(n_765), .A2(n_775), .B(n_776), .C(n_777), .Y(n_774) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
OAI21xp33_ASAP7_75t_SL g778 ( .A1(n_779), .A2(n_781), .B(n_782), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
AND2x2_ASAP7_75t_SL g813 ( .A(n_782), .B(n_814), .Y(n_813) );
OAI221xp5_ASAP7_75t_SL g783 ( .A1(n_784), .A2(n_786), .B1(n_787), .B2(n_788), .C(n_790), .Y(n_783) );
INVx1_ASAP7_75t_SL g787 ( .A(n_785), .Y(n_787) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
NAND3xp33_ASAP7_75t_SL g794 ( .A(n_795), .B(n_796), .C(n_803), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_797), .B(n_799), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
OAI21xp33_ASAP7_75t_L g807 ( .A1(n_808), .A2(n_810), .B(n_812), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVxp33_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_SL g816 ( .A(n_817), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_820), .Y(n_819) );
CKINVDCx11_ASAP7_75t_R g820 ( .A(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g829 ( .A(n_822), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g824 ( .A(n_825), .Y(n_824) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_833), .Y(n_831) );
CKINVDCx11_ASAP7_75t_R g833 ( .A(n_834), .Y(n_833) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_835), .Y(n_834) );
NOR2xp33_ASAP7_75t_L g836 ( .A(n_837), .B(n_838), .Y(n_836) );
endmodule