module fake_aes_10006_n_41 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_41);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
INVx2_ASAP7_75t_L g12 ( .A(n_7), .Y(n_12) );
AND2x4_ASAP7_75t_L g13 ( .A(n_10), .B(n_2), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_1), .Y(n_14) );
BUFx6f_ASAP7_75t_L g15 ( .A(n_4), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_5), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_9), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_1), .Y(n_18) );
NAND2xp5_ASAP7_75t_SL g19 ( .A(n_13), .B(n_0), .Y(n_19) );
NOR3xp33_ASAP7_75t_SL g20 ( .A(n_17), .B(n_0), .C(n_2), .Y(n_20) );
AND3x2_ASAP7_75t_SL g21 ( .A(n_12), .B(n_3), .C(n_4), .Y(n_21) );
INVx3_ASAP7_75t_L g22 ( .A(n_13), .Y(n_22) );
O2A1O1Ixp33_ASAP7_75t_SL g23 ( .A1(n_19), .A2(n_17), .B(n_18), .C(n_16), .Y(n_23) );
CKINVDCx5p33_ASAP7_75t_R g24 ( .A(n_20), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_22), .Y(n_25) );
NOR2xp67_ASAP7_75t_L g26 ( .A(n_24), .B(n_22), .Y(n_26) );
AND2x2_ASAP7_75t_L g27 ( .A(n_25), .B(n_19), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g28 ( .A(n_27), .B(n_25), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_27), .B(n_25), .Y(n_29) );
NOR3xp33_ASAP7_75t_SL g30 ( .A(n_28), .B(n_21), .C(n_26), .Y(n_30) );
AOI32xp33_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_14), .A3(n_21), .B1(n_23), .B2(n_7), .Y(n_31) );
OAI211xp5_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_15), .B(n_5), .C(n_6), .Y(n_32) );
NOR2xp33_ASAP7_75t_R g33 ( .A(n_30), .B(n_3), .Y(n_33) );
NAND2xp5_ASAP7_75t_L g34 ( .A(n_30), .B(n_15), .Y(n_34) );
INVxp67_ASAP7_75t_L g35 ( .A(n_34), .Y(n_35) );
NOR2x1_ASAP7_75t_L g36 ( .A(n_32), .B(n_15), .Y(n_36) );
NAND4xp25_ASAP7_75t_L g37 ( .A(n_33), .B(n_6), .C(n_8), .D(n_9), .Y(n_37) );
AOI31xp33_ASAP7_75t_L g38 ( .A1(n_36), .A2(n_8), .A3(n_10), .B(n_11), .Y(n_38) );
BUFx2_ASAP7_75t_L g39 ( .A(n_35), .Y(n_39) );
INVx1_ASAP7_75t_L g40 ( .A(n_39), .Y(n_40) );
AOI22xp5_ASAP7_75t_SL g41 ( .A1(n_40), .A2(n_39), .B1(n_38), .B2(n_37), .Y(n_41) );
endmodule