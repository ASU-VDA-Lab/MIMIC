module fake_jpeg_5444_n_104 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_104);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_104;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_22),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_39),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_24),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_3),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_17),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_0),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_64),
.A2(n_65),
.B(n_46),
.C(n_43),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_51),
.B(n_0),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_66),
.Y(n_70)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_64),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_69),
.B1(n_53),
.B2(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_58),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_59),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_78),
.Y(n_87)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_2),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_72),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_73),
.A2(n_61),
.B1(n_60),
.B2(n_52),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_79),
.A2(n_69),
.B1(n_68),
.B2(n_61),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_70),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_80),
.B(n_4),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_83),
.B1(n_85),
.B2(n_87),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_79),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_84),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_75),
.A2(n_47),
.B1(n_49),
.B2(n_48),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_1),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_86),
.Y(n_88)
);

OA21x2_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_91),
.B(n_4),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_54),
.C(n_6),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_92),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_95),
.A2(n_92),
.B1(n_94),
.B2(n_88),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_10),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_11),
.Y(n_98)
);

AOI322xp5_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_12),
.A3(n_13),
.B1(n_14),
.B2(n_16),
.C1(n_18),
.C2(n_20),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_99),
.A2(n_23),
.B(n_28),
.Y(n_100)
);

NOR4xp25_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_30),
.C(n_32),
.D(n_33),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_34),
.B(n_35),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_37),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_38),
.Y(n_104)
);


endmodule