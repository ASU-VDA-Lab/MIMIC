module fake_jpeg_26406_n_104 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_7),
.B(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_9),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_26),
.Y(n_30)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_28),
.Y(n_31)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_21),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_27),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_22),
.B1(n_13),
.B2(n_11),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_13),
.B1(n_18),
.B2(n_11),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_22),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_27),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_35),
.A2(n_13),
.B1(n_28),
.B2(n_14),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_39),
.B(n_47),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_40),
.B(n_41),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_36),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_43),
.B(n_46),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_23),
.Y(n_45)
);

AND2x6_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_1),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_17),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_15),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_18),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_50),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_49),
.A2(n_18),
.B1(n_19),
.B2(n_12),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_11),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_51),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_17),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_58),
.B(n_45),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_60),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_64),
.B1(n_60),
.B2(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_12),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_63),
.B(n_19),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_41),
.B(n_42),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_73),
.B(n_74),
.Y(n_77)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_75),
.Y(n_79)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_42),
.B(n_46),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_64),
.B1(n_55),
.B2(n_62),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_75),
.A2(n_58),
.B1(n_56),
.B2(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_78),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_56),
.C(n_59),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_80),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_59),
.C(n_57),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_46),
.B(n_43),
.C(n_16),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_14),
.B(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_69),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_89),
.Y(n_92)
);

AO21x1_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_43),
.B(n_16),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_87),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_71),
.B1(n_53),
.B2(n_21),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_83),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_8),
.Y(n_97)
);

XOR2x2_ASAP7_75t_SL g91 ( 
.A(n_88),
.B(n_78),
.Y(n_91)
);

AOI322xp5_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_93),
.A3(n_34),
.B1(n_8),
.B2(n_17),
.C1(n_5),
.C2(n_1),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_76),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_95),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_92),
.A2(n_86),
.B1(n_81),
.B2(n_21),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_34),
.C(n_2),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_1),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_2),
.C(n_3),
.Y(n_102)
);

AOI322xp5_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_94),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_102),
.C(n_100),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_4),
.Y(n_104)
);


endmodule