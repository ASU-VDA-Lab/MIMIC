module fake_ariane_1766_n_988 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_988);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_988;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_961;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_952;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_214;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_207;
wire n_790;
wire n_898;
wire n_857;
wire n_363;
wire n_720;
wire n_968;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_285;
wire n_473;
wire n_801;
wire n_202;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_903;
wire n_315;
wire n_871;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_485;
wire n_401;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_839;
wire n_928;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_277;
wire n_248;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_920;
wire n_899;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_455;
wire n_365;
wire n_429;
wire n_654;
wire n_588;
wire n_986;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_935;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_772;
wire n_747;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_966;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_213;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_583;
wire n_509;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_963;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_981;
wire n_882;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_289;
wire n_542;
wire n_548;
wire n_815;
wire n_973;
wire n_523;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_976;
wire n_909;
wire n_849;
wire n_353;
wire n_767;
wire n_736;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_80),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_3),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_54),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_45),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_84),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_113),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_70),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_83),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_146),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_127),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_26),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_93),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_86),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_57),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_40),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_134),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_153),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_165),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_52),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_119),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_123),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_105),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_142),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_106),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_49),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_25),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_78),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_91),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_177),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_79),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_174),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_60),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_154),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_46),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_3),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_162),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_32),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_103),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_122),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_115),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_108),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_69),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_120),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_56),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_61),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_64),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_22),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_58),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_110),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_43),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_124),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_19),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_41),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_125),
.Y(n_253)
);

BUFx10_ASAP7_75t_L g254 ( 
.A(n_111),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_143),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_71),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_167),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_0),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_6),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_36),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_173),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_196),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_74),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_160),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_18),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_169),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_89),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_172),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_63),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_95),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_55),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_178),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_112),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_23),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_23),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_101),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_200),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_225),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_204),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_259),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_224),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_224),
.Y(n_282)
);

NOR2xp67_ASAP7_75t_L g283 ( 
.A(n_234),
.B(n_0),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_232),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_232),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_205),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_215),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_217),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_220),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_241),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_207),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_265),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_246),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_254),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_238),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_254),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_259),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_251),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_198),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_199),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_208),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_204),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_258),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_212),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_274),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_275),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_213),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_201),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_213),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_221),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_226),
.B(n_1),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_230),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_239),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_244),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_240),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_253),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_244),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_202),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_216),
.B(n_1),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_256),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_260),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_261),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_262),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_267),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_203),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_206),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_209),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_264),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_210),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_279),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_302),
.B(n_268),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_279),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_299),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_309),
.B(n_229),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_300),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_301),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_304),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_310),
.Y(n_338)
);

BUFx8_ASAP7_75t_L g339 ( 
.A(n_277),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_312),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_313),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_315),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_316),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_320),
.Y(n_344)
);

OR2x6_ASAP7_75t_L g345 ( 
.A(n_296),
.B(n_219),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_321),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_322),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_324),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_292),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_297),
.Y(n_350)
);

NAND3xp33_ASAP7_75t_L g351 ( 
.A(n_311),
.B(n_249),
.C(n_229),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_280),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_328),
.B(n_270),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_323),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_283),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_295),
.Y(n_356)
);

AND2x4_ASAP7_75t_L g357 ( 
.A(n_298),
.B(n_278),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_293),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_308),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_329),
.Y(n_360)
);

AND2x4_ASAP7_75t_L g361 ( 
.A(n_325),
.B(n_249),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_326),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_307),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_303),
.B(n_236),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_305),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_307),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_306),
.B(n_222),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_314),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_314),
.Y(n_369)
);

AND2x4_ASAP7_75t_L g370 ( 
.A(n_317),
.B(n_237),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_317),
.B(n_272),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_319),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_327),
.B(n_271),
.Y(n_373)
);

NAND2xp33_ASAP7_75t_SL g374 ( 
.A(n_318),
.B(n_231),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_318),
.Y(n_375)
);

OA21x2_ASAP7_75t_L g376 ( 
.A1(n_286),
.A2(n_214),
.B(n_211),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_327),
.Y(n_377)
);

OA21x2_ASAP7_75t_L g378 ( 
.A1(n_287),
.A2(n_223),
.B(n_218),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_294),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_291),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_288),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_289),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_290),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_285),
.B(n_227),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_284),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_281),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_330),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_L g388 ( 
.A1(n_351),
.A2(n_231),
.B1(n_247),
.B2(n_263),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_348),
.Y(n_389)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_332),
.B(n_281),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_332),
.B(n_359),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_330),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_348),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_333),
.Y(n_394)
);

INVx5_ASAP7_75t_L g395 ( 
.A(n_348),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_330),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_333),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_330),
.Y(n_398)
);

OR2x2_ASAP7_75t_L g399 ( 
.A(n_352),
.B(n_282),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_332),
.B(n_2),
.Y(n_400)
);

NAND2xp33_ASAP7_75t_L g401 ( 
.A(n_359),
.B(n_231),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_330),
.Y(n_402)
);

INVx5_ASAP7_75t_L g403 ( 
.A(n_348),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_336),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_336),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_335),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_361),
.B(n_228),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_361),
.B(n_233),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_335),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_383),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_357),
.B(n_282),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_340),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_340),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_342),
.Y(n_414)
);

AND2x6_ASAP7_75t_L g415 ( 
.A(n_360),
.B(n_231),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_337),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_336),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_342),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_357),
.B(n_284),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_343),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_354),
.B(n_247),
.Y(n_421)
);

AND2x2_ASAP7_75t_SL g422 ( 
.A(n_370),
.B(n_371),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_343),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_337),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_346),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_338),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_346),
.Y(n_427)
);

AND3x2_ASAP7_75t_L g428 ( 
.A(n_370),
.B(n_2),
.C(n_4),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_357),
.B(n_235),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_361),
.B(n_242),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_357),
.B(n_243),
.Y(n_431)
);

BUFx10_ASAP7_75t_L g432 ( 
.A(n_367),
.Y(n_432)
);

INVx4_ASAP7_75t_L g433 ( 
.A(n_360),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_361),
.B(n_245),
.Y(n_434)
);

INVx5_ASAP7_75t_L g435 ( 
.A(n_350),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_338),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_341),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_334),
.B(n_4),
.Y(n_438)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_364),
.Y(n_439)
);

INVx4_ASAP7_75t_L g440 ( 
.A(n_360),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_354),
.B(n_248),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_364),
.B(n_250),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_383),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_341),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_344),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_344),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_347),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_347),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_349),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_334),
.B(n_252),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_349),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_350),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_373),
.A2(n_276),
.B1(n_273),
.B2(n_269),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_350),
.B(n_255),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_331),
.Y(n_455)
);

AND3x4_ASAP7_75t_L g456 ( 
.A(n_375),
.B(n_5),
.C(n_6),
.Y(n_456)
);

INVx4_ASAP7_75t_L g457 ( 
.A(n_345),
.Y(n_457)
);

OR2x2_ASAP7_75t_L g458 ( 
.A(n_353),
.B(n_5),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_355),
.B(n_257),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_345),
.B(n_355),
.Y(n_460)
);

NOR2xp67_ASAP7_75t_L g461 ( 
.A(n_443),
.B(n_382),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_389),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_445),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_389),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_410),
.B(n_363),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_445),
.Y(n_466)
);

NOR2xp67_ASAP7_75t_L g467 ( 
.A(n_443),
.B(n_382),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_409),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_409),
.Y(n_469)
);

NAND2x1p5_ASAP7_75t_L g470 ( 
.A(n_457),
.B(n_381),
.Y(n_470)
);

AO22x2_ASAP7_75t_L g471 ( 
.A1(n_456),
.A2(n_385),
.B1(n_372),
.B2(n_370),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_393),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_455),
.B(n_362),
.Y(n_473)
);

AO22x2_ASAP7_75t_L g474 ( 
.A1(n_456),
.A2(n_385),
.B1(n_372),
.B2(n_370),
.Y(n_474)
);

AO22x2_ASAP7_75t_L g475 ( 
.A1(n_411),
.A2(n_371),
.B1(n_366),
.B2(n_368),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_393),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_399),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_391),
.B(n_362),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_451),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_451),
.Y(n_480)
);

NAND2xp33_ASAP7_75t_L g481 ( 
.A(n_395),
.B(n_365),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_394),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_391),
.B(n_365),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_439),
.A2(n_374),
.B1(n_345),
.B2(n_351),
.Y(n_484)
);

NAND2x1p5_ASAP7_75t_L g485 ( 
.A(n_457),
.B(n_381),
.Y(n_485)
);

OAI221xp5_ASAP7_75t_L g486 ( 
.A1(n_458),
.A2(n_356),
.B1(n_345),
.B2(n_358),
.C(n_384),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_449),
.B(n_345),
.Y(n_487)
);

NAND2x1p5_ASAP7_75t_L g488 ( 
.A(n_460),
.B(n_381),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_397),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_412),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_449),
.B(n_358),
.Y(n_491)
);

AO22x2_ASAP7_75t_L g492 ( 
.A1(n_419),
.A2(n_371),
.B1(n_368),
.B2(n_366),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_409),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_460),
.B(n_381),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_409),
.Y(n_495)
);

AO22x2_ASAP7_75t_L g496 ( 
.A1(n_390),
.A2(n_371),
.B1(n_363),
.B2(n_375),
.Y(n_496)
);

AO22x2_ASAP7_75t_L g497 ( 
.A1(n_390),
.A2(n_369),
.B1(n_377),
.B2(n_380),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_433),
.B(n_376),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_460),
.A2(n_376),
.B1(n_378),
.B2(n_356),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_424),
.Y(n_500)
);

AO22x2_ASAP7_75t_L g501 ( 
.A1(n_438),
.A2(n_369),
.B1(n_377),
.B2(n_380),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_432),
.Y(n_502)
);

AO22x2_ASAP7_75t_L g503 ( 
.A1(n_438),
.A2(n_379),
.B1(n_386),
.B2(n_339),
.Y(n_503)
);

NAND2x1p5_ASAP7_75t_L g504 ( 
.A(n_422),
.B(n_381),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_413),
.Y(n_505)
);

NAND2x1p5_ASAP7_75t_L g506 ( 
.A(n_422),
.B(n_376),
.Y(n_506)
);

INVxp67_ASAP7_75t_SL g507 ( 
.A(n_400),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_433),
.B(n_440),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_440),
.B(n_376),
.Y(n_509)
);

AO22x2_ASAP7_75t_L g510 ( 
.A1(n_438),
.A2(n_379),
.B1(n_386),
.B2(n_339),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_429),
.B(n_386),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_424),
.Y(n_512)
);

AO22x2_ASAP7_75t_L g513 ( 
.A1(n_431),
.A2(n_386),
.B1(n_339),
.B2(n_378),
.Y(n_513)
);

NOR2xp67_ASAP7_75t_L g514 ( 
.A(n_435),
.B(n_386),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_414),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_418),
.Y(n_516)
);

AO22x2_ASAP7_75t_L g517 ( 
.A1(n_421),
.A2(n_339),
.B1(n_378),
.B2(n_9),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_424),
.Y(n_518)
);

AO22x2_ASAP7_75t_L g519 ( 
.A1(n_421),
.A2(n_378),
.B1(n_8),
.B2(n_9),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_420),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_423),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_452),
.B(n_266),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_425),
.Y(n_523)
);

NAND3xp33_ASAP7_75t_SL g524 ( 
.A(n_453),
.B(n_7),
.C(n_8),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_427),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_406),
.A2(n_247),
.B1(n_263),
.B2(n_11),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_452),
.B(n_247),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_406),
.Y(n_528)
);

AO22x2_ASAP7_75t_L g529 ( 
.A1(n_441),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_432),
.B(n_10),
.Y(n_530)
);

INVx8_ASAP7_75t_L g531 ( 
.A(n_415),
.Y(n_531)
);

NAND2x1p5_ASAP7_75t_L g532 ( 
.A(n_404),
.B(n_263),
.Y(n_532)
);

NAND2x1p5_ASAP7_75t_L g533 ( 
.A(n_404),
.B(n_263),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_405),
.B(n_12),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_400),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_416),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_405),
.B(n_12),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_416),
.Y(n_538)
);

OAI221xp5_ASAP7_75t_L g539 ( 
.A1(n_442),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.C(n_16),
.Y(n_539)
);

BUFx6f_ASAP7_75t_SL g540 ( 
.A(n_400),
.Y(n_540)
);

AO22x2_ASAP7_75t_L g541 ( 
.A1(n_428),
.A2(n_430),
.B1(n_407),
.B2(n_434),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_426),
.Y(n_542)
);

OAI221xp5_ASAP7_75t_L g543 ( 
.A1(n_450),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.C(n_16),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_426),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_494),
.B(n_435),
.Y(n_545)
);

NAND2xp33_ASAP7_75t_SL g546 ( 
.A(n_473),
.B(n_454),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_494),
.B(n_435),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_461),
.B(n_435),
.Y(n_548)
);

NAND2xp33_ASAP7_75t_SL g549 ( 
.A(n_502),
.B(n_408),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_467),
.B(n_417),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_478),
.B(n_417),
.Y(n_551)
);

NAND2xp33_ASAP7_75t_SL g552 ( 
.A(n_540),
.B(n_459),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_483),
.B(n_395),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_535),
.B(n_395),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_491),
.B(n_395),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_504),
.B(n_403),
.Y(n_556)
);

NAND2xp33_ASAP7_75t_SL g557 ( 
.A(n_530),
.B(n_424),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_484),
.B(n_403),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_SL g559 ( 
.A(n_487),
.B(n_437),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_465),
.B(n_436),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_488),
.B(n_403),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_511),
.B(n_403),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_507),
.B(n_437),
.Y(n_563)
);

NAND2xp33_ASAP7_75t_SL g564 ( 
.A(n_482),
.B(n_437),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_499),
.B(n_514),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_509),
.B(n_437),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_477),
.B(n_387),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_471),
.B(n_436),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_470),
.B(n_387),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_489),
.B(n_428),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_485),
.B(n_387),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_490),
.B(n_387),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_505),
.B(n_515),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_516),
.B(n_396),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_520),
.B(n_396),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_521),
.B(n_396),
.Y(n_576)
);

NAND2xp33_ASAP7_75t_SL g577 ( 
.A(n_523),
.B(n_396),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_525),
.B(n_444),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_498),
.B(n_398),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_506),
.B(n_398),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_463),
.B(n_444),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_466),
.B(n_398),
.Y(n_582)
);

NAND2xp33_ASAP7_75t_SL g583 ( 
.A(n_508),
.B(n_398),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_534),
.B(n_402),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_537),
.B(n_402),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_479),
.B(n_402),
.Y(n_586)
);

NAND2xp33_ASAP7_75t_SL g587 ( 
.A(n_522),
.B(n_402),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_468),
.B(n_446),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_480),
.B(n_392),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_462),
.B(n_446),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_464),
.B(n_447),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_469),
.B(n_392),
.Y(n_592)
);

NAND2xp33_ASAP7_75t_SL g593 ( 
.A(n_472),
.B(n_447),
.Y(n_593)
);

NAND2xp33_ASAP7_75t_SL g594 ( 
.A(n_476),
.B(n_448),
.Y(n_594)
);

NAND2xp33_ASAP7_75t_SL g595 ( 
.A(n_493),
.B(n_495),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_471),
.B(n_448),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_474),
.B(n_388),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_SL g598 ( 
.A(n_500),
.B(n_388),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_512),
.B(n_518),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_526),
.B(n_415),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_532),
.B(n_415),
.Y(n_601)
);

NAND2xp33_ASAP7_75t_SL g602 ( 
.A(n_529),
.B(n_415),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_533),
.B(n_415),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_528),
.B(n_401),
.Y(n_604)
);

NAND2xp33_ASAP7_75t_SL g605 ( 
.A(n_529),
.B(n_17),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_541),
.B(n_401),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_536),
.B(n_17),
.Y(n_607)
);

NAND2xp33_ASAP7_75t_SL g608 ( 
.A(n_486),
.B(n_18),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_538),
.B(n_19),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_542),
.B(n_20),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_581),
.Y(n_611)
);

OA21x2_ASAP7_75t_L g612 ( 
.A1(n_579),
.A2(n_527),
.B(n_544),
.Y(n_612)
);

BUFx4f_ASAP7_75t_SL g613 ( 
.A(n_570),
.Y(n_613)
);

NAND3x1_ASAP7_75t_L g614 ( 
.A(n_605),
.B(n_474),
.C(n_597),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_560),
.Y(n_615)
);

OAI21x1_ASAP7_75t_L g616 ( 
.A1(n_580),
.A2(n_524),
.B(n_481),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_573),
.Y(n_617)
);

OAI21x1_ASAP7_75t_L g618 ( 
.A1(n_566),
.A2(n_541),
.B(n_531),
.Y(n_618)
);

BUFx10_ASAP7_75t_L g619 ( 
.A(n_570),
.Y(n_619)
);

AO31x2_ASAP7_75t_L g620 ( 
.A1(n_606),
.A2(n_513),
.A3(n_519),
.B(n_517),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_578),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_588),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_581),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_610),
.A2(n_539),
.B1(n_543),
.B2(n_519),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_549),
.Y(n_625)
);

AO31x2_ASAP7_75t_L g626 ( 
.A1(n_590),
.A2(n_591),
.A3(n_565),
.B(n_598),
.Y(n_626)
);

OA21x2_ASAP7_75t_L g627 ( 
.A1(n_584),
.A2(n_513),
.B(n_517),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_588),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_551),
.A2(n_475),
.B(n_492),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_L g630 ( 
.A1(n_610),
.A2(n_475),
.B(n_492),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_567),
.B(n_531),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_568),
.B(n_503),
.Y(n_632)
);

AO21x1_ASAP7_75t_L g633 ( 
.A1(n_602),
.A2(n_510),
.B(n_503),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_596),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_552),
.Y(n_635)
);

NOR4xp25_ASAP7_75t_L g636 ( 
.A(n_609),
.B(n_501),
.C(n_510),
.D(n_497),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_546),
.A2(n_496),
.B(n_501),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_607),
.Y(n_638)
);

AOI21xp33_ASAP7_75t_L g639 ( 
.A1(n_558),
.A2(n_496),
.B(n_497),
.Y(n_639)
);

OAI21x1_ASAP7_75t_L g640 ( 
.A1(n_585),
.A2(n_118),
.B(n_195),
.Y(n_640)
);

AO31x2_ASAP7_75t_L g641 ( 
.A1(n_587),
.A2(n_117),
.A3(n_194),
.B(n_192),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_550),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_562),
.B(n_21),
.Y(n_643)
);

NAND2x1p5_ASAP7_75t_L g644 ( 
.A(n_545),
.B(n_27),
.Y(n_644)
);

NAND2xp33_ASAP7_75t_R g645 ( 
.A(n_608),
.B(n_28),
.Y(n_645)
);

OA21x2_ASAP7_75t_L g646 ( 
.A1(n_604),
.A2(n_126),
.B(n_191),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_564),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_547),
.B(n_24),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_599),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_556),
.B(n_24),
.Y(n_650)
);

A2O1A1Ixp33_ASAP7_75t_L g651 ( 
.A1(n_593),
.A2(n_25),
.B(n_29),
.C(n_30),
.Y(n_651)
);

OAI21x1_ASAP7_75t_L g652 ( 
.A1(n_553),
.A2(n_31),
.B(n_33),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_572),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_592),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_557),
.B(n_34),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_583),
.A2(n_35),
.B(n_37),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_574),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_594),
.A2(n_38),
.B(n_39),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_595),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_563),
.B(n_42),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_575),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_561),
.B(n_44),
.Y(n_662)
);

OAI22xp5_ASAP7_75t_L g663 ( 
.A1(n_600),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_555),
.A2(n_577),
.B(n_576),
.Y(n_664)
);

NAND2xp33_ASAP7_75t_L g665 ( 
.A(n_548),
.B(n_51),
.Y(n_665)
);

AOI221xp5_ASAP7_75t_L g666 ( 
.A1(n_624),
.A2(n_589),
.B1(n_559),
.B2(n_586),
.C(n_582),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_613),
.Y(n_667)
);

OAI21x1_ASAP7_75t_L g668 ( 
.A1(n_640),
.A2(n_571),
.B(n_569),
.Y(n_668)
);

AOI221xp5_ASAP7_75t_SL g669 ( 
.A1(n_642),
.A2(n_554),
.B1(n_603),
.B2(n_601),
.C(n_65),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_619),
.Y(n_670)
);

OA21x2_ASAP7_75t_L g671 ( 
.A1(n_630),
.A2(n_53),
.B(n_59),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_619),
.B(n_62),
.Y(n_672)
);

OAI21x1_ASAP7_75t_L g673 ( 
.A1(n_652),
.A2(n_66),
.B(n_67),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_626),
.Y(n_674)
);

AOI221x1_ASAP7_75t_L g675 ( 
.A1(n_624),
.A2(n_68),
.B1(n_72),
.B2(n_73),
.C(n_75),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_628),
.B(n_197),
.Y(n_676)
);

OA21x2_ASAP7_75t_L g677 ( 
.A1(n_630),
.A2(n_76),
.B(n_77),
.Y(n_677)
);

OA21x2_ASAP7_75t_L g678 ( 
.A1(n_637),
.A2(n_81),
.B(n_82),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_617),
.Y(n_679)
);

OAI21x1_ASAP7_75t_L g680 ( 
.A1(n_612),
.A2(n_85),
.B(n_87),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_615),
.B(n_88),
.Y(n_681)
);

OAI21x1_ASAP7_75t_L g682 ( 
.A1(n_612),
.A2(n_90),
.B(n_92),
.Y(n_682)
);

AOI221xp5_ASAP7_75t_L g683 ( 
.A1(n_636),
.A2(n_642),
.B1(n_639),
.B2(n_638),
.C(n_650),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_633),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_684)
);

O2A1O1Ixp33_ASAP7_75t_SL g685 ( 
.A1(n_651),
.A2(n_98),
.B(n_99),
.C(n_100),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_622),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_643),
.B(n_190),
.Y(n_687)
);

AOI221xp5_ASAP7_75t_L g688 ( 
.A1(n_636),
.A2(n_102),
.B1(n_104),
.B2(n_107),
.C(n_109),
.Y(n_688)
);

AO21x2_ASAP7_75t_L g689 ( 
.A1(n_629),
.A2(n_114),
.B(n_116),
.Y(n_689)
);

OAI21x1_ASAP7_75t_L g690 ( 
.A1(n_664),
.A2(n_121),
.B(n_128),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_625),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_648),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_639),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_693)
);

BUFx2_ASAP7_75t_L g694 ( 
.A(n_635),
.Y(n_694)
);

OAI21xp33_ASAP7_75t_SL g695 ( 
.A1(n_616),
.A2(n_132),
.B(n_133),
.Y(n_695)
);

O2A1O1Ixp33_ASAP7_75t_SL g696 ( 
.A1(n_655),
.A2(n_135),
.B(n_136),
.C(n_137),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_623),
.Y(n_697)
);

OAI21x1_ASAP7_75t_L g698 ( 
.A1(n_656),
.A2(n_138),
.B(n_139),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_611),
.Y(n_699)
);

AOI22x1_ASAP7_75t_L g700 ( 
.A1(n_647),
.A2(n_140),
.B1(n_141),
.B2(n_144),
.Y(n_700)
);

OAI21x1_ASAP7_75t_L g701 ( 
.A1(n_618),
.A2(n_145),
.B(n_147),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_634),
.Y(n_702)
);

AO31x2_ASAP7_75t_L g703 ( 
.A1(n_663),
.A2(n_632),
.A3(n_621),
.B(n_658),
.Y(n_703)
);

OA21x2_ASAP7_75t_L g704 ( 
.A1(n_629),
.A2(n_148),
.B(n_149),
.Y(n_704)
);

OA21x2_ASAP7_75t_L g705 ( 
.A1(n_653),
.A2(n_150),
.B(n_151),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_649),
.Y(n_706)
);

AOI21x1_ASAP7_75t_L g707 ( 
.A1(n_660),
.A2(n_152),
.B(n_155),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_SL g708 ( 
.A(n_628),
.B(n_156),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_626),
.Y(n_709)
);

INVxp67_ASAP7_75t_L g710 ( 
.A(n_622),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_627),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_711)
);

OAI21x1_ASAP7_75t_L g712 ( 
.A1(n_646),
.A2(n_161),
.B(n_163),
.Y(n_712)
);

OAI21x1_ASAP7_75t_L g713 ( 
.A1(n_646),
.A2(n_164),
.B(n_166),
.Y(n_713)
);

AO21x2_ASAP7_75t_L g714 ( 
.A1(n_657),
.A2(n_661),
.B(n_663),
.Y(n_714)
);

AO31x2_ASAP7_75t_L g715 ( 
.A1(n_626),
.A2(n_168),
.A3(n_171),
.B(n_175),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_650),
.Y(n_716)
);

AO22x2_ASAP7_75t_L g717 ( 
.A1(n_620),
.A2(n_176),
.B1(n_179),
.B2(n_180),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_622),
.B(n_189),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_627),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_647),
.B(n_184),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_674),
.Y(n_721)
);

AOI222xp33_ASAP7_75t_L g722 ( 
.A1(n_683),
.A2(n_662),
.B1(n_614),
.B2(n_645),
.C1(n_659),
.C2(n_665),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_716),
.A2(n_662),
.B1(n_631),
.B2(n_654),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_674),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_679),
.Y(n_725)
);

BUFx2_ASAP7_75t_L g726 ( 
.A(n_714),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_697),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_709),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_SL g729 ( 
.A(n_667),
.B(n_644),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_709),
.Y(n_730)
);

OR2x6_ASAP7_75t_L g731 ( 
.A(n_717),
.B(n_677),
.Y(n_731)
);

AOI21xp33_ASAP7_75t_L g732 ( 
.A1(n_692),
.A2(n_654),
.B(n_620),
.Y(n_732)
);

BUFx2_ASAP7_75t_L g733 ( 
.A(n_714),
.Y(n_733)
);

OAI21x1_ASAP7_75t_L g734 ( 
.A1(n_680),
.A2(n_641),
.B(n_654),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_694),
.A2(n_620),
.B1(n_641),
.B2(n_187),
.Y(n_735)
);

AO21x2_ASAP7_75t_L g736 ( 
.A1(n_689),
.A2(n_641),
.B(n_186),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_715),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_667),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_702),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_715),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_686),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_715),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_706),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_699),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_705),
.Y(n_745)
);

HB1xp67_ASAP7_75t_L g746 ( 
.A(n_686),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_705),
.Y(n_747)
);

INVx1_ASAP7_75t_SL g748 ( 
.A(n_691),
.Y(n_748)
);

HB1xp67_ASAP7_75t_L g749 ( 
.A(n_686),
.Y(n_749)
);

BUFx2_ASAP7_75t_L g750 ( 
.A(n_703),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_705),
.Y(n_751)
);

OA21x2_ASAP7_75t_L g752 ( 
.A1(n_675),
.A2(n_185),
.B(n_188),
.Y(n_752)
);

AO31x2_ASAP7_75t_L g753 ( 
.A1(n_717),
.A2(n_718),
.A3(n_677),
.B(n_671),
.Y(n_753)
);

OAI21xp5_ASAP7_75t_L g754 ( 
.A1(n_666),
.A2(n_669),
.B(n_695),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_710),
.Y(n_755)
);

INVxp67_ASAP7_75t_SL g756 ( 
.A(n_671),
.Y(n_756)
);

OR2x2_ASAP7_75t_L g757 ( 
.A(n_703),
.B(n_710),
.Y(n_757)
);

AOI21x1_ASAP7_75t_L g758 ( 
.A1(n_707),
.A2(n_668),
.B(n_682),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_717),
.B(n_687),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_671),
.Y(n_760)
);

AO21x2_ASAP7_75t_L g761 ( 
.A1(n_689),
.A2(n_713),
.B(n_712),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_686),
.Y(n_762)
);

INVxp67_ASAP7_75t_SL g763 ( 
.A(n_677),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_720),
.B(n_703),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_681),
.Y(n_765)
);

OA21x2_ASAP7_75t_L g766 ( 
.A1(n_701),
.A2(n_719),
.B(n_711),
.Y(n_766)
);

BUFx2_ASAP7_75t_L g767 ( 
.A(n_703),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_678),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_720),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_678),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_720),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_678),
.Y(n_772)
);

AOI222xp33_ASAP7_75t_L g773 ( 
.A1(n_688),
.A2(n_693),
.B1(n_684),
.B2(n_719),
.C1(n_711),
.C2(n_708),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_676),
.B(n_670),
.Y(n_774)
);

CKINVDCx20_ASAP7_75t_R g775 ( 
.A(n_691),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_670),
.Y(n_776)
);

INVx2_ASAP7_75t_SL g777 ( 
.A(n_676),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_704),
.B(n_684),
.Y(n_778)
);

OAI21x1_ASAP7_75t_L g779 ( 
.A1(n_698),
.A2(n_690),
.B(n_673),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_672),
.B(n_693),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_739),
.B(n_704),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_725),
.B(n_704),
.Y(n_782)
);

XNOR2xp5_ASAP7_75t_SL g783 ( 
.A(n_775),
.B(n_696),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_765),
.B(n_700),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_727),
.B(n_755),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_743),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_774),
.B(n_685),
.Y(n_787)
);

INVxp67_ASAP7_75t_L g788 ( 
.A(n_741),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_R g789 ( 
.A(n_775),
.B(n_696),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_746),
.B(n_685),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_744),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_777),
.B(n_774),
.Y(n_792)
);

BUFx10_ASAP7_75t_L g793 ( 
.A(n_774),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_749),
.B(n_762),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_738),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_R g796 ( 
.A(n_738),
.B(n_777),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_769),
.B(n_771),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_776),
.B(n_764),
.Y(n_798)
);

NAND2xp33_ASAP7_75t_R g799 ( 
.A(n_731),
.B(n_759),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_757),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_748),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_R g802 ( 
.A(n_729),
.B(n_750),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_731),
.B(n_723),
.Y(n_803)
);

INVxp67_ASAP7_75t_L g804 ( 
.A(n_722),
.Y(n_804)
);

NAND2xp33_ASAP7_75t_R g805 ( 
.A(n_731),
.B(n_778),
.Y(n_805)
);

NAND2xp33_ASAP7_75t_R g806 ( 
.A(n_731),
.B(n_778),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_780),
.B(n_750),
.Y(n_807)
);

AND2x4_ASAP7_75t_L g808 ( 
.A(n_721),
.B(n_724),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_767),
.B(n_732),
.Y(n_809)
);

NAND2xp33_ASAP7_75t_R g810 ( 
.A(n_752),
.B(n_766),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_721),
.B(n_724),
.Y(n_811)
);

XOR2x2_ASAP7_75t_SL g812 ( 
.A(n_735),
.B(n_773),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_767),
.B(n_726),
.Y(n_813)
);

NAND2xp33_ASAP7_75t_R g814 ( 
.A(n_752),
.B(n_766),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_728),
.B(n_730),
.Y(n_815)
);

NAND2xp33_ASAP7_75t_R g816 ( 
.A(n_752),
.B(n_766),
.Y(n_816)
);

INVxp67_ASAP7_75t_L g817 ( 
.A(n_726),
.Y(n_817)
);

NAND2xp33_ASAP7_75t_R g818 ( 
.A(n_733),
.B(n_754),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_733),
.B(n_734),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_760),
.B(n_751),
.Y(n_820)
);

NAND2xp33_ASAP7_75t_SL g821 ( 
.A(n_736),
.B(n_760),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_R g822 ( 
.A(n_758),
.B(n_742),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_728),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_756),
.B(n_763),
.Y(n_824)
);

NAND2xp33_ASAP7_75t_R g825 ( 
.A(n_737),
.B(n_740),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_745),
.B(n_751),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_730),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_737),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_740),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_798),
.B(n_742),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_813),
.B(n_753),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_828),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_808),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_800),
.B(n_753),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_827),
.Y(n_835)
);

INVx1_ASAP7_75t_SL g836 ( 
.A(n_795),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_785),
.B(n_753),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_808),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_829),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_811),
.Y(n_840)
);

INVxp67_ASAP7_75t_L g841 ( 
.A(n_794),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_787),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_807),
.B(n_753),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_819),
.B(n_753),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_804),
.A2(n_736),
.B1(n_761),
.B2(n_772),
.Y(n_845)
);

BUFx2_ASAP7_75t_L g846 ( 
.A(n_822),
.Y(n_846)
);

INVx4_ASAP7_75t_L g847 ( 
.A(n_787),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_786),
.B(n_745),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_791),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_788),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_811),
.Y(n_851)
);

NAND2x1p5_ASAP7_75t_SL g852 ( 
.A(n_790),
.B(n_747),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_781),
.B(n_747),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_815),
.Y(n_854)
);

INVx4_ASAP7_75t_L g855 ( 
.A(n_795),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_797),
.B(n_768),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_815),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_820),
.Y(n_858)
);

INVxp67_ASAP7_75t_L g859 ( 
.A(n_795),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_782),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_797),
.B(n_768),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_823),
.B(n_736),
.Y(n_862)
);

INVxp67_ASAP7_75t_L g863 ( 
.A(n_801),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_826),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_817),
.B(n_770),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_792),
.B(n_761),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_793),
.B(n_758),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_818),
.A2(n_770),
.B1(n_772),
.B2(n_761),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_842),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_831),
.B(n_824),
.Y(n_870)
);

OAI21xp33_ASAP7_75t_SL g871 ( 
.A1(n_847),
.A2(n_784),
.B(n_783),
.Y(n_871)
);

BUFx2_ASAP7_75t_L g872 ( 
.A(n_846),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_832),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_831),
.B(n_803),
.Y(n_874)
);

OAI21x1_ASAP7_75t_L g875 ( 
.A1(n_845),
.A2(n_734),
.B(n_862),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_837),
.B(n_809),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_850),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_844),
.B(n_803),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_832),
.Y(n_879)
);

INVxp67_ASAP7_75t_L g880 ( 
.A(n_833),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_846),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_860),
.B(n_796),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_835),
.Y(n_883)
);

BUFx2_ASAP7_75t_L g884 ( 
.A(n_852),
.Y(n_884)
);

OAI31xp33_ASAP7_75t_SL g885 ( 
.A1(n_844),
.A2(n_812),
.A3(n_789),
.B(n_816),
.Y(n_885)
);

OAI33xp33_ASAP7_75t_L g886 ( 
.A1(n_858),
.A2(n_814),
.A3(n_810),
.B1(n_799),
.B2(n_825),
.B3(n_805),
.Y(n_886)
);

OAI31xp33_ASAP7_75t_L g887 ( 
.A1(n_843),
.A2(n_821),
.A3(n_806),
.B(n_802),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_839),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_868),
.A2(n_779),
.B1(n_793),
.B2(n_843),
.Y(n_889)
);

BUFx2_ASAP7_75t_L g890 ( 
.A(n_852),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_841),
.B(n_779),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_835),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_855),
.Y(n_893)
);

AND2x2_ASAP7_75t_SL g894 ( 
.A(n_868),
.B(n_847),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_842),
.B(n_847),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_839),
.Y(n_896)
);

INVxp67_ASAP7_75t_SL g897 ( 
.A(n_884),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_883),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_883),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_892),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_872),
.B(n_842),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_873),
.Y(n_902)
);

OR2x2_ASAP7_75t_L g903 ( 
.A(n_876),
.B(n_852),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_870),
.B(n_858),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_873),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_879),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_872),
.B(n_842),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_881),
.B(n_847),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_881),
.B(n_863),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_879),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_870),
.B(n_860),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_888),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_908),
.B(n_881),
.Y(n_913)
);

NAND2xp33_ASAP7_75t_SL g914 ( 
.A(n_909),
.B(n_877),
.Y(n_914)
);

NAND2xp33_ASAP7_75t_SL g915 ( 
.A(n_909),
.B(n_869),
.Y(n_915)
);

NOR2xp67_ASAP7_75t_L g916 ( 
.A(n_903),
.B(n_871),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_904),
.B(n_871),
.Y(n_917)
);

NOR4xp25_ASAP7_75t_SL g918 ( 
.A(n_897),
.B(n_890),
.C(n_884),
.D(n_896),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_908),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_911),
.B(n_891),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_903),
.B(n_891),
.Y(n_921)
);

NOR2x1_ASAP7_75t_L g922 ( 
.A(n_901),
.B(n_890),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_R g923 ( 
.A(n_901),
.B(n_893),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_912),
.B(n_876),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_924),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_917),
.A2(n_894),
.B1(n_889),
.B2(n_895),
.Y(n_926)
);

OR2x2_ASAP7_75t_L g927 ( 
.A(n_920),
.B(n_910),
.Y(n_927)
);

INVx1_ASAP7_75t_SL g928 ( 
.A(n_914),
.Y(n_928)
);

CKINVDCx16_ASAP7_75t_R g929 ( 
.A(n_923),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_913),
.B(n_907),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_919),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_921),
.Y(n_932)
);

OR2x2_ASAP7_75t_L g933 ( 
.A(n_917),
.B(n_906),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_916),
.B(n_907),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_922),
.Y(n_935)
);

OAI21xp33_ASAP7_75t_SL g936 ( 
.A1(n_928),
.A2(n_894),
.B(n_918),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_925),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_927),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_932),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_933),
.B(n_905),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_937),
.Y(n_941)
);

OAI221xp5_ASAP7_75t_L g942 ( 
.A1(n_936),
.A2(n_926),
.B1(n_928),
.B2(n_885),
.C(n_889),
.Y(n_942)
);

NAND2x1p5_ASAP7_75t_L g943 ( 
.A(n_939),
.B(n_931),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_941),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_943),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_942),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_941),
.Y(n_947)
);

AND3x2_ASAP7_75t_L g948 ( 
.A(n_944),
.B(n_935),
.C(n_934),
.Y(n_948)
);

NOR3xp33_ASAP7_75t_L g949 ( 
.A(n_946),
.B(n_929),
.C(n_926),
.Y(n_949)
);

NOR3xp33_ASAP7_75t_L g950 ( 
.A(n_945),
.B(n_938),
.C(n_940),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_947),
.B(n_930),
.Y(n_951)
);

NAND4xp25_ASAP7_75t_L g952 ( 
.A(n_945),
.B(n_915),
.C(n_893),
.D(n_895),
.Y(n_952)
);

INVx1_ASAP7_75t_SL g953 ( 
.A(n_945),
.Y(n_953)
);

NOR3xp33_ASAP7_75t_L g954 ( 
.A(n_946),
.B(n_886),
.C(n_882),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_948),
.Y(n_955)
);

INVx1_ASAP7_75t_SL g956 ( 
.A(n_953),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_949),
.A2(n_875),
.B(n_887),
.C(n_894),
.Y(n_957)
);

OAI311xp33_ASAP7_75t_L g958 ( 
.A1(n_951),
.A2(n_952),
.A3(n_950),
.B1(n_954),
.C1(n_866),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_953),
.A2(n_902),
.B1(n_896),
.B2(n_888),
.Y(n_959)
);

AOI221xp5_ASAP7_75t_L g960 ( 
.A1(n_953),
.A2(n_864),
.B1(n_867),
.B2(n_834),
.C(n_900),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_956),
.B(n_895),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_955),
.B(n_895),
.Y(n_962)
);

AO22x1_ASAP7_75t_L g963 ( 
.A1(n_955),
.A2(n_869),
.B1(n_855),
.B2(n_836),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_957),
.B(n_869),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_959),
.Y(n_965)
);

NOR2xp67_ASAP7_75t_L g966 ( 
.A(n_958),
.B(n_869),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_R g967 ( 
.A(n_965),
.B(n_855),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_961),
.B(n_960),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_962),
.B(n_855),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_964),
.B(n_859),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_R g971 ( 
.A(n_963),
.B(n_851),
.Y(n_971)
);

NAND2xp33_ASAP7_75t_L g972 ( 
.A(n_967),
.B(n_966),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_968),
.B(n_900),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_969),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_970),
.A2(n_971),
.B(n_875),
.Y(n_975)
);

XNOR2xp5_ASAP7_75t_L g976 ( 
.A(n_973),
.B(n_874),
.Y(n_976)
);

OA22x2_ASAP7_75t_L g977 ( 
.A1(n_974),
.A2(n_864),
.B1(n_898),
.B2(n_899),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_972),
.A2(n_899),
.B(n_898),
.Y(n_978)
);

OAI21xp33_ASAP7_75t_SL g979 ( 
.A1(n_977),
.A2(n_975),
.B(n_978),
.Y(n_979)
);

AOI31xp33_ASAP7_75t_L g980 ( 
.A1(n_976),
.A2(n_874),
.A3(n_878),
.B(n_851),
.Y(n_980)
);

AOI31xp33_ASAP7_75t_L g981 ( 
.A1(n_979),
.A2(n_878),
.A3(n_880),
.B(n_833),
.Y(n_981)
);

AOI31xp33_ASAP7_75t_L g982 ( 
.A1(n_980),
.A2(n_838),
.A3(n_840),
.B(n_849),
.Y(n_982)
);

OAI322xp33_ASAP7_75t_L g983 ( 
.A1(n_981),
.A2(n_849),
.A3(n_892),
.B1(n_835),
.B2(n_840),
.C1(n_838),
.C2(n_848),
.Y(n_983)
);

AOI222xp33_ASAP7_75t_SL g984 ( 
.A1(n_983),
.A2(n_982),
.B1(n_854),
.B2(n_857),
.C1(n_865),
.C2(n_834),
.Y(n_984)
);

OAI22xp33_ASAP7_75t_L g985 ( 
.A1(n_983),
.A2(n_853),
.B1(n_857),
.B2(n_854),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_985),
.Y(n_986)
);

OAI221xp5_ASAP7_75t_R g987 ( 
.A1(n_986),
.A2(n_984),
.B1(n_865),
.B2(n_848),
.C(n_853),
.Y(n_987)
);

AOI211xp5_ASAP7_75t_L g988 ( 
.A1(n_987),
.A2(n_856),
.B(n_861),
.C(n_830),
.Y(n_988)
);


endmodule