module fake_jpeg_20961_n_313 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_27),
.Y(n_37)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_38),
.Y(n_48)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_31),
.Y(n_56)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp33_ASAP7_75t_SL g44 ( 
.A(n_17),
.B(n_8),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_44),
.B(n_35),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_39),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_46),
.A2(n_29),
.B(n_30),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_59),
.Y(n_71)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_24),
.B1(n_23),
.B2(n_19),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_50),
.A2(n_55),
.B1(n_37),
.B2(n_41),
.Y(n_76)
);

INVx2_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_51),
.A2(n_43),
.B1(n_33),
.B2(n_28),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_24),
.B1(n_23),
.B2(n_19),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_36),
.A2(n_24),
.B1(n_34),
.B2(n_25),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_60),
.B1(n_35),
.B2(n_16),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_34),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_36),
.A2(n_16),
.B1(n_32),
.B2(n_25),
.Y(n_60)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_65),
.B(n_99),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_41),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_66),
.B(n_74),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_70),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_18),
.B(n_22),
.C(n_20),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_72),
.B(n_79),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_32),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_73),
.B(n_77),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_41),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_76),
.A2(n_83),
.B1(n_94),
.B2(n_100),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_22),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_80),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_60),
.B(n_18),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_53),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_SL g81 ( 
.A1(n_51),
.A2(n_37),
.B(n_39),
.C(n_41),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_81),
.A2(n_103),
.B(n_95),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_20),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_82),
.B(n_85),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_50),
.A2(n_37),
.B1(n_42),
.B2(n_40),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_42),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_87),
.A2(n_104),
.B(n_61),
.Y(n_117)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_31),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_89),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_45),
.B(n_31),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_90),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_20),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_98),
.Y(n_105)
);

BUFx4f_ASAP7_75t_SL g92 ( 
.A(n_48),
.Y(n_92)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_55),
.A2(n_40),
.B1(n_42),
.B2(n_37),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_52),
.A2(n_29),
.B1(n_30),
.B2(n_38),
.Y(n_96)
);

NOR2x1_ASAP7_75t_R g115 ( 
.A(n_96),
.B(n_97),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_31),
.Y(n_98)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_52),
.A2(n_42),
.B1(n_40),
.B2(n_38),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_61),
.A2(n_38),
.B1(n_30),
.B2(n_29),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_101),
.A2(n_102),
.B1(n_61),
.B2(n_62),
.Y(n_112)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_52),
.A2(n_40),
.B1(n_42),
.B2(n_57),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_103),
.A2(n_62),
.B1(n_54),
.B2(n_43),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_112),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_70),
.B(n_86),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_71),
.B(n_43),
.C(n_62),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_119),
.C(n_96),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g159 ( 
.A1(n_117),
.A2(n_105),
.B1(n_134),
.B2(n_120),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_28),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_81),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_66),
.B(n_12),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_120),
.A2(n_121),
.B1(n_128),
.B2(n_83),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_74),
.A2(n_54),
.B1(n_43),
.B2(n_28),
.Y(n_121)
);

OAI32xp33_ASAP7_75t_L g124 ( 
.A1(n_72),
.A2(n_28),
.A3(n_26),
.B1(n_21),
.B2(n_17),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_104),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_65),
.A2(n_43),
.B1(n_26),
.B2(n_21),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_107),
.B(n_87),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_135),
.B(n_161),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_136),
.B(n_165),
.Y(n_186)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_138),
.A2(n_139),
.B1(n_142),
.B2(n_146),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_114),
.A2(n_115),
.B1(n_124),
.B2(n_131),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_140),
.A2(n_143),
.B1(n_150),
.B2(n_157),
.Y(n_169)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_129),
.A2(n_87),
.B1(n_69),
.B2(n_104),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_127),
.A2(n_69),
.B1(n_104),
.B2(n_81),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_128),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_81),
.B1(n_64),
.B2(n_88),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_118),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_153),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_149),
.A2(n_111),
.B1(n_123),
.B2(n_122),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_129),
.A2(n_75),
.B1(n_67),
.B2(n_85),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_113),
.Y(n_152)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_108),
.B(n_78),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_92),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_155),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_67),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_123),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_160),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_127),
.A2(n_99),
.B1(n_92),
.B2(n_26),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_115),
.B(n_133),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_158),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_121),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_105),
.B(n_84),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_26),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_21),
.Y(n_162)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_105),
.A2(n_21),
.B1(n_17),
.B2(n_2),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_163),
.A2(n_164),
.B1(n_0),
.B2(n_2),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_117),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_107),
.B(n_0),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_141),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_168),
.B(n_172),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_132),
.B(n_119),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_170),
.A2(n_182),
.B(n_183),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

AND2x6_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_106),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_179),
.Y(n_207)
);

AND2x6_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_106),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_181),
.B(n_195),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_142),
.Y(n_183)
);

XNOR2x2_ASAP7_75t_L g185 ( 
.A(n_135),
.B(n_130),
.Y(n_185)
);

XNOR2x1_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_15),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_188),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_110),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_190),
.B(n_157),
.Y(n_205)
);

OA21x2_ASAP7_75t_L g191 ( 
.A1(n_138),
.A2(n_147),
.B(n_159),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_182),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_143),
.A2(n_134),
.B1(n_110),
.B2(n_132),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_192),
.A2(n_164),
.B1(n_163),
.B2(n_156),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_194),
.Y(n_197)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_144),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_196),
.B(n_122),
.Y(n_215)
);

O2A1O1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_198),
.A2(n_201),
.B(n_0),
.C(n_3),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_181),
.A2(n_155),
.B(n_150),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_136),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_204),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_145),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_205),
.A2(n_169),
.B1(n_191),
.B2(n_192),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_189),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_206),
.B(n_209),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_208),
.A2(n_169),
.B1(n_205),
.B2(n_172),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_153),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_166),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_211),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_193),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_137),
.C(n_139),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_214),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_173),
.B(n_152),
.C(n_111),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_215),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_167),
.B(n_165),
.Y(n_216)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

NAND3xp33_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_185),
.C(n_179),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_175),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_218),
.B(n_178),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_177),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_220),
.Y(n_227)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_180),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_222),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_174),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_194),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_191),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_229),
.Y(n_257)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_219),
.Y(n_231)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_231),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_234),
.A2(n_243),
.B1(n_217),
.B2(n_201),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_197),
.A2(n_183),
.B1(n_223),
.B2(n_206),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_238),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_190),
.Y(n_240)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_213),
.A2(n_176),
.B1(n_170),
.B2(n_4),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_212),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_176),
.Y(n_242)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_208),
.Y(n_254)
);

FAx1_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_212),
.CI(n_236),
.CON(n_246),
.SN(n_246)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_246),
.A2(n_250),
.B1(n_243),
.B2(n_231),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_226),
.B(n_207),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_248),
.Y(n_275)
);

NAND2x1_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_244),
.Y(n_250)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_254),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_256),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_204),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_202),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_263),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_199),
.C(n_209),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_233),
.C(n_237),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_199),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_227),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_198),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_272),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_247),
.A2(n_225),
.B1(n_240),
.B2(n_232),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_267),
.A2(n_253),
.B1(n_246),
.B2(n_249),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_257),
.A2(n_232),
.B1(n_227),
.B2(n_240),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_245),
.B(n_261),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_269),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_271),
.A2(n_246),
.B(n_262),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_220),
.C(n_222),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_272),
.C(n_270),
.Y(n_279)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_258),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_254),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_250),
.A2(n_10),
.B1(n_3),
.B2(n_5),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_281),
.C(n_285),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_280),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_259),
.C(n_263),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_288),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_271),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_10),
.C(n_5),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_266),
.A2(n_11),
.B(n_6),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_274),
.A2(n_6),
.B(n_9),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_275),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_298),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_264),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_294),
.Y(n_303)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_292),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_267),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_270),
.C(n_264),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_284),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_6),
.Y(n_298)
);

AOI21x1_ASAP7_75t_SL g299 ( 
.A1(n_295),
.A2(n_282),
.B(n_287),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_301),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_296),
.A2(n_287),
.B1(n_281),
.B2(n_285),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_293),
.C(n_298),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_305),
.A2(n_306),
.B(n_302),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_293),
.Y(n_306)
);

AOI321xp33_ASAP7_75t_L g310 ( 
.A1(n_308),
.A2(n_309),
.A3(n_301),
.B1(n_299),
.B2(n_290),
.C(n_14),
.Y(n_310)
);

NOR2x1_ASAP7_75t_L g309 ( 
.A(n_307),
.B(n_300),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_310),
.A2(n_10),
.B(n_13),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_15),
.B(n_14),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_312),
.B(n_0),
.Y(n_313)
);


endmodule