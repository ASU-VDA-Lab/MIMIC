module real_aes_7593_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_725;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g179 ( .A1(n_0), .A2(n_180), .B(n_181), .C(n_185), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_1), .B(n_174), .Y(n_187) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_2), .B(n_92), .C(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g126 ( .A(n_2), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_3), .B(n_159), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_4), .A2(n_168), .B(n_480), .Y(n_479) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_5), .A2(n_148), .B(n_165), .C(n_524), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_6), .A2(n_168), .B(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_7), .B(n_174), .Y(n_486) );
AO21x2_ASAP7_75t_L g261 ( .A1(n_8), .A2(n_140), .B(n_262), .Y(n_261) );
AND2x6_ASAP7_75t_L g165 ( .A(n_9), .B(n_166), .Y(n_165) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_10), .A2(n_148), .B(n_165), .C(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g577 ( .A(n_11), .Y(n_577) );
INVx1_ASAP7_75t_L g110 ( .A(n_12), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_12), .B(n_39), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_13), .B(n_184), .Y(n_526) );
INVx1_ASAP7_75t_L g145 ( .A(n_14), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_15), .B(n_159), .Y(n_268) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_16), .A2(n_160), .B(n_535), .C(n_537), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_17), .B(n_174), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_18), .B(n_202), .Y(n_500) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_19), .A2(n_148), .B(n_194), .C(n_201), .Y(n_193) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_20), .A2(n_183), .B(n_236), .C(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_21), .B(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_22), .B(n_184), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_23), .B(n_184), .Y(n_475) );
CKINVDCx16_ASAP7_75t_R g504 ( .A(n_24), .Y(n_504) );
INVx1_ASAP7_75t_L g474 ( .A(n_25), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_26), .A2(n_148), .B(n_201), .C(n_265), .Y(n_264) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_27), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_28), .Y(n_522) );
INVx1_ASAP7_75t_L g498 ( .A(n_29), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_30), .A2(n_168), .B(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g150 ( .A(n_31), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_32), .A2(n_163), .B(n_217), .C(n_218), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_33), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_34), .A2(n_183), .B(n_483), .C(n_485), .Y(n_482) );
INVxp67_ASAP7_75t_L g499 ( .A(n_35), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_36), .B(n_267), .Y(n_266) );
CKINVDCx14_ASAP7_75t_R g481 ( .A(n_37), .Y(n_481) );
A2O1A1Ixp33_ASAP7_75t_L g472 ( .A1(n_38), .A2(n_148), .B(n_201), .C(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_39), .B(n_110), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g574 ( .A1(n_40), .A2(n_185), .B(n_575), .C(n_576), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_41), .B(n_192), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_42), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_43), .B(n_159), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_44), .B(n_168), .Y(n_263) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_45), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_46), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_47), .A2(n_163), .B(n_217), .C(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g182 ( .A(n_48), .Y(n_182) );
AOI22xp33_ASAP7_75t_L g128 ( .A1(n_49), .A2(n_129), .B1(n_443), .B2(n_444), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_49), .Y(n_443) );
INVx1_ASAP7_75t_L g246 ( .A(n_50), .Y(n_246) );
INVx1_ASAP7_75t_L g542 ( .A(n_51), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_52), .B(n_168), .Y(n_243) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_53), .A2(n_72), .B1(n_131), .B2(n_132), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_53), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g206 ( .A(n_54), .Y(n_206) );
AOI222xp33_ASAP7_75t_SL g449 ( .A1(n_55), .A2(n_450), .B1(n_456), .B2(n_726), .C1(n_727), .C2(n_728), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_56), .A2(n_104), .B1(n_115), .B2(n_732), .Y(n_103) );
CKINVDCx14_ASAP7_75t_R g573 ( .A(n_57), .Y(n_573) );
INVx1_ASAP7_75t_L g166 ( .A(n_58), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_59), .B(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_60), .B(n_174), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_61), .A2(n_155), .B(n_200), .C(n_257), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g453 ( .A1(n_62), .A2(n_71), .B1(n_454), .B2(n_455), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_62), .Y(n_454) );
INVx1_ASAP7_75t_L g144 ( .A(n_63), .Y(n_144) );
INVx1_ASAP7_75t_SL g484 ( .A(n_64), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_65), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_66), .B(n_159), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_67), .B(n_174), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_68), .B(n_160), .Y(n_233) );
INVx1_ASAP7_75t_L g507 ( .A(n_69), .Y(n_507) );
CKINVDCx16_ASAP7_75t_R g177 ( .A(n_70), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_71), .Y(n_455) );
INVx1_ASAP7_75t_L g132 ( .A(n_72), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_73), .B(n_196), .Y(n_195) );
A2O1A1Ixp33_ASAP7_75t_L g147 ( .A1(n_74), .A2(n_148), .B(n_153), .C(n_163), .Y(n_147) );
CKINVDCx16_ASAP7_75t_R g255 ( .A(n_75), .Y(n_255) );
INVx1_ASAP7_75t_L g114 ( .A(n_76), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_77), .A2(n_168), .B(n_572), .Y(n_571) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_78), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_79), .A2(n_168), .B(n_532), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_80), .A2(n_192), .B(n_494), .Y(n_493) );
CKINVDCx16_ASAP7_75t_R g471 ( .A(n_81), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_82), .A2(n_451), .B1(n_452), .B2(n_453), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_82), .Y(n_451) );
INVx1_ASAP7_75t_L g533 ( .A(n_83), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_84), .B(n_198), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_85), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_86), .A2(n_168), .B(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g536 ( .A(n_87), .Y(n_536) );
INVx2_ASAP7_75t_L g142 ( .A(n_88), .Y(n_142) );
INVx1_ASAP7_75t_L g525 ( .A(n_89), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_90), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_91), .B(n_184), .Y(n_234) );
OR2x2_ASAP7_75t_L g123 ( .A(n_92), .B(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g460 ( .A(n_92), .B(n_125), .Y(n_460) );
INVx2_ASAP7_75t_L g725 ( .A(n_92), .Y(n_725) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_93), .A2(n_148), .B(n_163), .C(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_94), .B(n_168), .Y(n_215) );
INVx1_ASAP7_75t_L g219 ( .A(n_95), .Y(n_219) );
INVxp67_ASAP7_75t_L g258 ( .A(n_96), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_97), .B(n_140), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_98), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g154 ( .A(n_99), .Y(n_154) );
INVx1_ASAP7_75t_L g229 ( .A(n_100), .Y(n_229) );
INVx2_ASAP7_75t_L g545 ( .A(n_101), .Y(n_545) );
AND2x2_ASAP7_75t_L g248 ( .A(n_102), .B(n_204), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
CKINVDCx6p67_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_107), .Y(n_733) );
CKINVDCx9p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_448), .Y(n_115) );
BUFx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
NAND3xp33_ASAP7_75t_L g448 ( .A(n_117), .B(n_445), .C(n_449), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_128), .B(n_445), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_123), .Y(n_447) );
NOR2x2_ASAP7_75t_L g726 ( .A(n_124), .B(n_725), .Y(n_726) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g724 ( .A(n_125), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
INVx1_ASAP7_75t_L g444 ( .A(n_129), .Y(n_444) );
XNOR2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_133), .Y(n_129) );
INVx1_ASAP7_75t_L g457 ( .A(n_133), .Y(n_457) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_133), .A2(n_462), .B1(n_729), .B2(n_730), .Y(n_728) );
OR3x1_ASAP7_75t_L g133 ( .A(n_134), .B(n_351), .C(n_400), .Y(n_133) );
NAND5xp2_ASAP7_75t_L g134 ( .A(n_135), .B(n_285), .C(n_314), .D(n_322), .E(n_337), .Y(n_134) );
O2A1O1Ixp33_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_208), .B(n_224), .C(n_269), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_137), .B(n_188), .Y(n_136) );
AND2x2_ASAP7_75t_L g280 ( .A(n_137), .B(n_277), .Y(n_280) );
AND2x2_ASAP7_75t_L g313 ( .A(n_137), .B(n_189), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_137), .B(n_212), .Y(n_406) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_173), .Y(n_137) );
INVx2_ASAP7_75t_L g211 ( .A(n_138), .Y(n_211) );
BUFx2_ASAP7_75t_L g380 ( .A(n_138), .Y(n_380) );
AO21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_146), .B(n_171), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_139), .B(n_172), .Y(n_171) );
INVx3_ASAP7_75t_L g174 ( .A(n_139), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_139), .B(n_223), .Y(n_222) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_139), .A2(n_228), .B(n_238), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_139), .B(n_477), .Y(n_476) );
AO21x2_ASAP7_75t_L g502 ( .A1(n_139), .A2(n_503), .B(n_510), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_139), .B(n_528), .Y(n_527) );
INVx4_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_140), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_140), .A2(n_263), .B(n_264), .Y(n_262) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g240 ( .A(n_141), .Y(n_240) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
AND2x2_ASAP7_75t_SL g204 ( .A(n_142), .B(n_143), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_167), .Y(n_146) );
INVx5_ASAP7_75t_L g178 ( .A(n_148), .Y(n_178) );
AND2x6_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_149), .Y(n_162) );
BUFx3_ASAP7_75t_L g186 ( .A(n_149), .Y(n_186) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g170 ( .A(n_150), .Y(n_170) );
INVx1_ASAP7_75t_L g237 ( .A(n_150), .Y(n_237) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_152), .Y(n_157) );
INVx3_ASAP7_75t_L g160 ( .A(n_152), .Y(n_160) );
AND2x2_ASAP7_75t_L g169 ( .A(n_152), .B(n_170), .Y(n_169) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_152), .Y(n_184) );
INVx1_ASAP7_75t_L g267 ( .A(n_152), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .B(n_158), .C(n_161), .Y(n_153) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
OAI22xp33_ASAP7_75t_L g497 ( .A1(n_156), .A2(n_159), .B1(n_498), .B2(n_499), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_156), .B(n_536), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_156), .B(n_545), .Y(n_544) );
INVx4_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g196 ( .A(n_157), .Y(n_196) );
INVx2_ASAP7_75t_L g180 ( .A(n_159), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_159), .B(n_258), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_159), .A2(n_199), .B(n_474), .C(n_475), .Y(n_473) );
INVx5_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_160), .B(n_577), .Y(n_576) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx3_ASAP7_75t_L g485 ( .A(n_162), .Y(n_485) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
O2A1O1Ixp33_ASAP7_75t_SL g176 ( .A1(n_164), .A2(n_177), .B(n_178), .C(n_179), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_L g254 ( .A1(n_164), .A2(n_178), .B(n_255), .C(n_256), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_L g480 ( .A1(n_164), .A2(n_178), .B(n_481), .C(n_482), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_SL g494 ( .A1(n_164), .A2(n_178), .B(n_495), .C(n_496), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_SL g532 ( .A1(n_164), .A2(n_178), .B(n_533), .C(n_534), .Y(n_532) );
O2A1O1Ixp33_ASAP7_75t_SL g541 ( .A1(n_164), .A2(n_178), .B(n_542), .C(n_543), .Y(n_541) );
O2A1O1Ixp33_ASAP7_75t_SL g572 ( .A1(n_164), .A2(n_178), .B(n_573), .C(n_574), .Y(n_572) );
INVx4_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
AND2x4_ASAP7_75t_L g168 ( .A(n_165), .B(n_169), .Y(n_168) );
BUFx3_ASAP7_75t_L g201 ( .A(n_165), .Y(n_201) );
NAND2x1p5_ASAP7_75t_L g230 ( .A(n_165), .B(n_169), .Y(n_230) );
BUFx2_ASAP7_75t_L g192 ( .A(n_168), .Y(n_192) );
INVx1_ASAP7_75t_L g200 ( .A(n_170), .Y(n_200) );
AND2x2_ASAP7_75t_L g188 ( .A(n_173), .B(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g278 ( .A(n_173), .Y(n_278) );
AND2x2_ASAP7_75t_L g364 ( .A(n_173), .B(n_277), .Y(n_364) );
AND2x2_ASAP7_75t_L g419 ( .A(n_173), .B(n_211), .Y(n_419) );
OA21x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_187), .Y(n_173) );
INVx2_ASAP7_75t_L g217 ( .A(n_178), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_183), .B(n_484), .Y(n_483) );
INVx4_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g575 ( .A(n_184), .Y(n_575) );
INVx2_ASAP7_75t_L g509 ( .A(n_185), .Y(n_509) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_186), .Y(n_221) );
INVx1_ASAP7_75t_L g537 ( .A(n_186), .Y(n_537) );
INVx1_ASAP7_75t_L g336 ( .A(n_188), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_188), .B(n_212), .Y(n_383) );
INVx5_ASAP7_75t_L g277 ( .A(n_189), .Y(n_277) );
AND2x4_ASAP7_75t_L g298 ( .A(n_189), .B(n_278), .Y(n_298) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_189), .Y(n_320) );
AND2x2_ASAP7_75t_L g395 ( .A(n_189), .B(n_380), .Y(n_395) );
AND2x2_ASAP7_75t_L g398 ( .A(n_189), .B(n_213), .Y(n_398) );
OR2x6_ASAP7_75t_L g189 ( .A(n_190), .B(n_205), .Y(n_189) );
AOI21xp5_ASAP7_75t_SL g190 ( .A1(n_191), .A2(n_193), .B(n_202), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_197), .B(n_199), .Y(n_194) );
INVx2_ASAP7_75t_L g198 ( .A(n_196), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_L g218 ( .A1(n_198), .A2(n_219), .B(n_220), .C(n_221), .Y(n_218) );
O2A1O1Ixp33_ASAP7_75t_L g245 ( .A1(n_198), .A2(n_221), .B(n_246), .C(n_247), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g506 ( .A1(n_198), .A2(n_507), .B(n_508), .C(n_509), .Y(n_506) );
O2A1O1Ixp5_ASAP7_75t_L g524 ( .A1(n_198), .A2(n_509), .B(n_525), .C(n_526), .Y(n_524) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_200), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_203), .B(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g207 ( .A(n_204), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_204), .A2(n_215), .B(n_216), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_204), .A2(n_243), .B(n_244), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_204), .A2(n_230), .B(n_471), .C(n_472), .Y(n_470) );
OA21x2_ASAP7_75t_L g570 ( .A1(n_204), .A2(n_571), .B(n_578), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_207), .A2(n_521), .B(n_527), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_208), .B(n_278), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_208), .B(n_409), .Y(n_408) );
INVx2_ASAP7_75t_SL g208 ( .A(n_209), .Y(n_208) );
OR2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_212), .Y(n_209) );
AND2x2_ASAP7_75t_L g303 ( .A(n_210), .B(n_278), .Y(n_303) );
AND2x2_ASAP7_75t_L g321 ( .A(n_210), .B(n_213), .Y(n_321) );
INVx1_ASAP7_75t_L g341 ( .A(n_210), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_210), .B(n_277), .Y(n_386) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_210), .Y(n_428) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_211), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_212), .B(n_276), .Y(n_275) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_212), .Y(n_330) );
O2A1O1Ixp33_ASAP7_75t_L g333 ( .A1(n_212), .A2(n_273), .B(n_334), .C(n_336), .Y(n_333) );
AND2x2_ASAP7_75t_L g340 ( .A(n_212), .B(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g349 ( .A(n_212), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g353 ( .A(n_212), .B(n_277), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_212), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g368 ( .A(n_212), .B(n_278), .Y(n_368) );
AND2x2_ASAP7_75t_L g418 ( .A(n_212), .B(n_419), .Y(n_418) );
INVx5_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
BUFx2_ASAP7_75t_L g282 ( .A(n_213), .Y(n_282) );
AND2x2_ASAP7_75t_L g323 ( .A(n_213), .B(n_276), .Y(n_323) );
AND2x2_ASAP7_75t_L g335 ( .A(n_213), .B(n_310), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_213), .B(n_364), .Y(n_382) );
OR2x6_ASAP7_75t_L g213 ( .A(n_214), .B(n_222), .Y(n_213) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_249), .Y(n_224) );
INVx1_ASAP7_75t_L g271 ( .A(n_225), .Y(n_271) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_241), .Y(n_225) );
OR2x2_ASAP7_75t_L g273 ( .A(n_226), .B(n_241), .Y(n_273) );
NAND3xp33_ASAP7_75t_L g279 ( .A(n_226), .B(n_280), .C(n_281), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_226), .B(n_251), .Y(n_290) );
OR2x2_ASAP7_75t_L g305 ( .A(n_226), .B(n_293), .Y(n_305) );
AND2x2_ASAP7_75t_L g311 ( .A(n_226), .B(n_260), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_226), .B(n_442), .Y(n_441) );
INVx5_ASAP7_75t_SL g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_227), .B(n_251), .Y(n_308) );
AND2x2_ASAP7_75t_L g347 ( .A(n_227), .B(n_261), .Y(n_347) );
NAND2xp5_ASAP7_75t_SL g375 ( .A(n_227), .B(n_260), .Y(n_375) );
OR2x2_ASAP7_75t_L g378 ( .A(n_227), .B(n_260), .Y(n_378) );
OAI21xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_231), .Y(n_228) );
OAI21xp5_ASAP7_75t_L g503 ( .A1(n_230), .A2(n_504), .B(n_505), .Y(n_503) );
OAI21xp5_ASAP7_75t_L g521 ( .A1(n_230), .A2(n_522), .B(n_523), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_235), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_235), .A2(n_266), .B(n_268), .Y(n_265) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
INVx2_ASAP7_75t_L g492 ( .A(n_240), .Y(n_492) );
INVx5_ASAP7_75t_SL g293 ( .A(n_241), .Y(n_293) );
OR2x2_ASAP7_75t_L g299 ( .A(n_241), .B(n_250), .Y(n_299) );
AND2x2_ASAP7_75t_L g315 ( .A(n_241), .B(n_316), .Y(n_315) );
AOI321xp33_ASAP7_75t_L g322 ( .A1(n_241), .A2(n_323), .A3(n_324), .B1(n_325), .B2(n_331), .C(n_333), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_241), .B(n_249), .Y(n_332) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_241), .Y(n_345) );
OR2x2_ASAP7_75t_L g392 ( .A(n_241), .B(n_290), .Y(n_392) );
AND2x2_ASAP7_75t_L g414 ( .A(n_241), .B(n_311), .Y(n_414) );
AND2x2_ASAP7_75t_L g433 ( .A(n_241), .B(n_251), .Y(n_433) );
OR2x6_ASAP7_75t_L g241 ( .A(n_242), .B(n_248), .Y(n_241) );
INVx1_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_260), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_251), .B(n_260), .Y(n_274) );
AND2x2_ASAP7_75t_L g283 ( .A(n_251), .B(n_284), .Y(n_283) );
INVx3_ASAP7_75t_L g310 ( .A(n_251), .Y(n_310) );
AND2x2_ASAP7_75t_L g316 ( .A(n_251), .B(n_311), .Y(n_316) );
INVxp67_ASAP7_75t_L g346 ( .A(n_251), .Y(n_346) );
OR2x2_ASAP7_75t_L g388 ( .A(n_251), .B(n_293), .Y(n_388) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_253), .B(n_259), .Y(n_251) );
OA21x2_ASAP7_75t_L g478 ( .A1(n_252), .A2(n_479), .B(n_486), .Y(n_478) );
OA21x2_ASAP7_75t_L g530 ( .A1(n_252), .A2(n_531), .B(n_538), .Y(n_530) );
OA21x2_ASAP7_75t_L g539 ( .A1(n_252), .A2(n_540), .B(n_546), .Y(n_539) );
OR2x2_ASAP7_75t_L g270 ( .A(n_260), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_SL g284 ( .A(n_260), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_260), .B(n_273), .Y(n_317) );
AND2x2_ASAP7_75t_L g366 ( .A(n_260), .B(n_310), .Y(n_366) );
AND2x2_ASAP7_75t_L g404 ( .A(n_260), .B(n_293), .Y(n_404) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_261), .B(n_293), .Y(n_292) );
A2O1A1Ixp33_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_272), .B(n_275), .C(n_279), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_270), .A2(n_272), .B1(n_397), .B2(n_399), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_272), .A2(n_295), .B1(n_350), .B2(n_436), .Y(n_435) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVx1_ASAP7_75t_SL g424 ( .A(n_273), .Y(n_424) );
INVx1_ASAP7_75t_SL g324 ( .A(n_274), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_276), .B(n_296), .Y(n_326) );
AOI222xp33_ASAP7_75t_L g337 ( .A1(n_276), .A2(n_317), .B1(n_324), .B2(n_338), .C1(n_342), .C2(n_348), .Y(n_337) );
AND2x2_ASAP7_75t_L g427 ( .A(n_276), .B(n_428), .Y(n_427) );
AND2x4_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx2_ASAP7_75t_L g302 ( .A(n_277), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_277), .B(n_297), .Y(n_372) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_277), .Y(n_409) );
AND2x2_ASAP7_75t_L g412 ( .A(n_277), .B(n_321), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_277), .B(n_428), .Y(n_438) );
INVx1_ASAP7_75t_L g329 ( .A(n_278), .Y(n_329) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_278), .Y(n_357) );
O2A1O1Ixp33_ASAP7_75t_L g420 ( .A1(n_280), .A2(n_421), .B(n_422), .C(n_425), .Y(n_420) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
NAND3xp33_ASAP7_75t_L g343 ( .A(n_282), .B(n_344), .C(n_347), .Y(n_343) );
OR2x2_ASAP7_75t_L g371 ( .A(n_282), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_282), .B(n_298), .Y(n_399) );
OR2x2_ASAP7_75t_L g304 ( .A(n_284), .B(n_305), .Y(n_304) );
AOI211xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_288), .B(n_294), .C(n_306), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_287), .B(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g393 ( .A(n_288), .B(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_289), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g307 ( .A(n_292), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_293), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g361 ( .A(n_293), .B(n_311), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_293), .B(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_293), .B(n_310), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_299), .B1(n_300), .B2(n_304), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_296), .B(n_368), .Y(n_367) );
BUFx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_298), .B(n_340), .Y(n_339) );
OAI221xp5_ASAP7_75t_SL g362 ( .A1(n_299), .A2(n_363), .B1(n_365), .B2(n_367), .C(n_369), .Y(n_362) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
AND2x2_ASAP7_75t_L g417 ( .A(n_302), .B(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g430 ( .A(n_302), .B(n_419), .Y(n_430) );
INVx1_ASAP7_75t_L g350 ( .A(n_303), .Y(n_350) );
INVx1_ASAP7_75t_L g421 ( .A(n_304), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g410 ( .A1(n_305), .A2(n_388), .B(n_411), .Y(n_410) );
AOI21xp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_309), .B(n_312), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OAI21xp5_ASAP7_75t_SL g314 ( .A1(n_315), .A2(n_317), .B(n_318), .Y(n_314) );
INVx1_ASAP7_75t_L g354 ( .A(n_315), .Y(n_354) );
AOI221xp5_ASAP7_75t_L g401 ( .A1(n_316), .A2(n_402), .B1(n_405), .B2(n_407), .C(n_410), .Y(n_401) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g413 ( .A1(n_324), .A2(n_414), .B1(n_415), .B2(n_417), .Y(n_413) );
NAND2xp5_ASAP7_75t_SL g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVx1_ASAP7_75t_L g390 ( .A(n_326), .Y(n_390) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NOR2xp67_ASAP7_75t_SL g328 ( .A(n_329), .B(n_330), .Y(n_328) );
AND2x2_ASAP7_75t_L g394 ( .A(n_330), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g359 ( .A(n_335), .Y(n_359) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_340), .B(n_364), .Y(n_416) );
INVxp67_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_346), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g432 ( .A(n_347), .B(n_433), .Y(n_432) );
AND2x4_ASAP7_75t_L g439 ( .A(n_347), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OAI211xp5_ASAP7_75t_SL g351 ( .A1(n_352), .A2(n_354), .B(n_355), .C(n_389), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AOI211xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_358), .B(n_362), .C(n_381), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_SL g442 ( .A(n_366), .Y(n_442) );
AND2x2_ASAP7_75t_L g379 ( .A(n_368), .B(n_380), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_373), .B1(n_377), .B2(n_379), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
OR2x2_ASAP7_75t_L g387 ( .A(n_375), .B(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g440 ( .A(n_376), .Y(n_440) );
INVxp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AOI31xp33_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_383), .A3(n_384), .B(n_387), .Y(n_381) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AOI211xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B(n_393), .C(n_396), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
CKINVDCx16_ASAP7_75t_R g397 ( .A(n_398), .Y(n_397) );
NAND5xp2_ASAP7_75t_L g400 ( .A(n_401), .B(n_413), .C(n_420), .D(n_434), .E(n_437), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_412), .A2(n_438), .B1(n_439), .B2(n_441), .Y(n_437) );
INVx1_ASAP7_75t_SL g436 ( .A(n_414), .Y(n_436) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AOI21xp33_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_429), .B(n_431), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVxp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
CKINVDCx16_ASAP7_75t_R g727 ( .A(n_450), .Y(n_727) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OAI22xp5_ASAP7_75t_SL g456 ( .A1(n_457), .A2(n_458), .B1(n_461), .B2(n_724), .Y(n_456) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g729 ( .A(n_459), .Y(n_729) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OR3x1_ASAP7_75t_L g462 ( .A(n_463), .B(n_635), .C(n_682), .Y(n_462) );
NAND3xp33_ASAP7_75t_SL g463 ( .A(n_464), .B(n_581), .C(n_606), .Y(n_463) );
AOI221xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_519), .B1(n_547), .B2(n_550), .C(n_558), .Y(n_464) );
OAI21xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_487), .B(n_512), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_467), .B(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_467), .B(n_563), .Y(n_679) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_478), .Y(n_467) );
AND2x2_ASAP7_75t_L g549 ( .A(n_468), .B(n_518), .Y(n_549) );
AND2x2_ASAP7_75t_L g599 ( .A(n_468), .B(n_517), .Y(n_599) );
AND2x2_ASAP7_75t_L g620 ( .A(n_468), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g625 ( .A(n_468), .B(n_592), .Y(n_625) );
OR2x2_ASAP7_75t_L g633 ( .A(n_468), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g705 ( .A(n_468), .B(n_501), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_468), .B(n_654), .Y(n_719) );
INVx3_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g564 ( .A(n_469), .B(n_478), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_469), .B(n_501), .Y(n_565) );
AND2x4_ASAP7_75t_L g587 ( .A(n_469), .B(n_518), .Y(n_587) );
AND2x2_ASAP7_75t_L g617 ( .A(n_469), .B(n_489), .Y(n_617) );
AND2x2_ASAP7_75t_L g626 ( .A(n_469), .B(n_616), .Y(n_626) );
AND2x2_ASAP7_75t_L g642 ( .A(n_469), .B(n_502), .Y(n_642) );
OR2x2_ASAP7_75t_L g651 ( .A(n_469), .B(n_634), .Y(n_651) );
AND2x2_ASAP7_75t_L g657 ( .A(n_469), .B(n_592), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_469), .B(n_663), .Y(n_662) );
OR2x2_ASAP7_75t_L g671 ( .A(n_469), .B(n_514), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_469), .B(n_560), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g710 ( .A(n_469), .B(n_621), .Y(n_710) );
OR2x6_ASAP7_75t_L g469 ( .A(n_470), .B(n_476), .Y(n_469) );
INVx2_ASAP7_75t_L g518 ( .A(n_478), .Y(n_518) );
AND2x2_ASAP7_75t_L g616 ( .A(n_478), .B(n_501), .Y(n_616) );
AND2x2_ASAP7_75t_L g621 ( .A(n_478), .B(n_502), .Y(n_621) );
INVx1_ASAP7_75t_L g677 ( .A(n_478), .Y(n_677) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g586 ( .A(n_488), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_501), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_489), .B(n_549), .Y(n_548) );
BUFx3_ASAP7_75t_L g563 ( .A(n_489), .Y(n_563) );
OR2x2_ASAP7_75t_L g634 ( .A(n_489), .B(n_501), .Y(n_634) );
OR2x2_ASAP7_75t_L g695 ( .A(n_489), .B(n_602), .Y(n_695) );
OA21x2_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_493), .B(n_500), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AO21x2_ASAP7_75t_L g514 ( .A1(n_491), .A2(n_515), .B(n_516), .Y(n_514) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g515 ( .A(n_493), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_500), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_501), .B(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g654 ( .A(n_501), .B(n_514), .Y(n_654) );
INVx2_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
BUFx2_ASAP7_75t_L g593 ( .A(n_502), .Y(n_593) );
INVx1_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_513), .A2(n_699), .B1(n_703), .B2(n_706), .C(n_707), .Y(n_698) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_517), .Y(n_513) );
INVx1_ASAP7_75t_SL g561 ( .A(n_514), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_514), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g693 ( .A(n_514), .B(n_549), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_517), .B(n_563), .Y(n_685) );
AND2x2_ASAP7_75t_L g592 ( .A(n_518), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_SL g596 ( .A(n_519), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_519), .B(n_602), .Y(n_632) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_529), .Y(n_519) );
AND2x2_ASAP7_75t_L g557 ( .A(n_520), .B(n_530), .Y(n_557) );
INVx4_ASAP7_75t_L g569 ( .A(n_520), .Y(n_569) );
BUFx3_ASAP7_75t_L g612 ( .A(n_520), .Y(n_612) );
AND3x2_ASAP7_75t_L g627 ( .A(n_520), .B(n_628), .C(n_629), .Y(n_627) );
AND2x2_ASAP7_75t_L g709 ( .A(n_529), .B(n_623), .Y(n_709) );
AND2x2_ASAP7_75t_L g717 ( .A(n_529), .B(n_602), .Y(n_717) );
INVx1_ASAP7_75t_SL g722 ( .A(n_529), .Y(n_722) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_539), .Y(n_529) );
INVx1_ASAP7_75t_SL g580 ( .A(n_530), .Y(n_580) );
AND2x2_ASAP7_75t_L g603 ( .A(n_530), .B(n_569), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_530), .B(n_553), .Y(n_605) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_530), .Y(n_645) );
OR2x2_ASAP7_75t_L g650 ( .A(n_530), .B(n_569), .Y(n_650) );
INVx2_ASAP7_75t_L g555 ( .A(n_539), .Y(n_555) );
AND2x2_ASAP7_75t_L g590 ( .A(n_539), .B(n_570), .Y(n_590) );
OR2x2_ASAP7_75t_L g610 ( .A(n_539), .B(n_570), .Y(n_610) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_539), .Y(n_630) );
INVx1_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
AOI21xp33_ASAP7_75t_L g680 ( .A1(n_548), .A2(n_589), .B(n_681), .Y(n_680) );
AOI322xp5_ASAP7_75t_L g716 ( .A1(n_550), .A2(n_560), .A3(n_587), .B1(n_717), .B2(n_718), .C1(n_720), .C2(n_723), .Y(n_716) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_556), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_552), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_553), .B(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g579 ( .A(n_554), .B(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g647 ( .A(n_555), .B(n_569), .Y(n_647) );
AND2x2_ASAP7_75t_L g714 ( .A(n_555), .B(n_570), .Y(n_714) );
INVx1_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g655 ( .A(n_557), .B(n_609), .Y(n_655) );
AOI31xp33_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_562), .A3(n_565), .B(n_566), .Y(n_558) );
AND2x2_ASAP7_75t_L g614 ( .A(n_560), .B(n_592), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_560), .B(n_584), .Y(n_696) );
AND2x2_ASAP7_75t_L g715 ( .A(n_560), .B(n_620), .Y(n_715) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_563), .B(n_592), .Y(n_604) );
NAND2x1p5_ASAP7_75t_L g638 ( .A(n_563), .B(n_621), .Y(n_638) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_563), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_563), .B(n_705), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_564), .B(n_621), .Y(n_653) );
INVx1_ASAP7_75t_L g697 ( .A(n_564), .Y(n_697) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_579), .Y(n_567) );
INVxp67_ASAP7_75t_L g649 ( .A(n_568), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_569), .B(n_580), .Y(n_585) );
INVx1_ASAP7_75t_L g691 ( .A(n_569), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_569), .B(n_668), .Y(n_702) );
BUFx3_ASAP7_75t_L g602 ( .A(n_570), .Y(n_602) );
AND2x2_ASAP7_75t_L g628 ( .A(n_570), .B(n_580), .Y(n_628) );
INVx2_ASAP7_75t_L g668 ( .A(n_570), .Y(n_668) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_579), .B(n_701), .Y(n_700) );
AOI211xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_586), .B(n_588), .C(n_597), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AOI21xp33_ASAP7_75t_L g631 ( .A1(n_583), .A2(n_632), .B(n_633), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_584), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_584), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g664 ( .A(n_585), .B(n_610), .Y(n_664) );
INVx3_ASAP7_75t_L g595 ( .A(n_587), .Y(n_595) );
OAI22xp5_ASAP7_75t_SL g588 ( .A1(n_589), .A2(n_591), .B1(n_594), .B2(n_596), .Y(n_588) );
OAI21xp5_ASAP7_75t_SL g613 ( .A1(n_590), .A2(n_614), .B(n_615), .Y(n_613) );
AND2x2_ASAP7_75t_L g639 ( .A(n_590), .B(n_603), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_590), .B(n_691), .Y(n_690) );
INVxp67_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OR2x2_ASAP7_75t_L g594 ( .A(n_593), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g663 ( .A(n_593), .Y(n_663) );
OAI21xp5_ASAP7_75t_SL g607 ( .A1(n_594), .A2(n_608), .B(n_613), .Y(n_607) );
OAI22xp33_ASAP7_75t_SL g597 ( .A1(n_598), .A2(n_600), .B1(n_604), .B2(n_605), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_599), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
INVx1_ASAP7_75t_L g623 ( .A(n_602), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_602), .B(n_645), .Y(n_644) );
NOR3xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_618), .C(n_631), .Y(n_606) );
OAI22xp5_ASAP7_75t_SL g673 ( .A1(n_608), .A2(n_674), .B1(n_678), .B2(n_679), .Y(n_673) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_609), .B(n_611), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OR2x2_ASAP7_75t_L g678 ( .A(n_610), .B(n_611), .Y(n_678) );
AND2x2_ASAP7_75t_L g686 ( .A(n_611), .B(n_667), .Y(n_686) );
CKINVDCx16_ASAP7_75t_R g611 ( .A(n_612), .Y(n_611) );
O2A1O1Ixp33_ASAP7_75t_SL g694 ( .A1(n_612), .A2(n_695), .B(n_696), .C(n_697), .Y(n_694) );
OR2x2_ASAP7_75t_L g721 ( .A(n_612), .B(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
OAI21xp33_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_622), .B(n_624), .Y(n_618) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
O2A1O1Ixp33_ASAP7_75t_L g656 ( .A1(n_620), .A2(n_657), .B(n_658), .C(n_661), .Y(n_656) );
OAI21xp33_ASAP7_75t_SL g624 ( .A1(n_625), .A2(n_626), .B(n_627), .Y(n_624) );
AND2x2_ASAP7_75t_L g689 ( .A(n_628), .B(n_647), .Y(n_689) );
INVxp67_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g667 ( .A(n_630), .B(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g672 ( .A(n_632), .Y(n_672) );
NAND3xp33_ASAP7_75t_SL g635 ( .A(n_636), .B(n_656), .C(n_669), .Y(n_635) );
AOI211xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_639), .B(n_640), .C(n_648), .Y(n_636) );
INVx1_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
INVx1_ASAP7_75t_L g706 ( .A(n_643), .Y(n_706) );
OR2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_646), .Y(n_643) );
INVx1_ASAP7_75t_L g666 ( .A(n_645), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_645), .B(n_714), .Y(n_713) );
INVxp67_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
A2O1A1Ixp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_650), .B(n_651), .C(n_652), .Y(n_648) );
INVx2_ASAP7_75t_SL g660 ( .A(n_650), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_651), .A2(n_662), .B1(n_664), .B2(n_665), .Y(n_661) );
OAI21xp33_ASAP7_75t_SL g652 ( .A1(n_653), .A2(n_654), .B(n_655), .Y(n_652) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
AOI211xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_672), .B(n_673), .C(n_680), .Y(n_669) );
INVx1_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
INVxp33_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g723 ( .A(n_677), .Y(n_723) );
NAND4xp25_ASAP7_75t_L g682 ( .A(n_683), .B(n_698), .C(n_711), .D(n_716), .Y(n_682) );
AOI211xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_686), .B(n_687), .C(n_694), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_690), .B(n_692), .Y(n_687) );
AOI21xp33_ASAP7_75t_L g707 ( .A1(n_688), .A2(n_708), .B(n_710), .Y(n_707) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_695), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_715), .Y(n_711) );
INVxp67_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g731 ( .A(n_724), .Y(n_731) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_733), .Y(n_732) );
endmodule