module fake_jpeg_6984_n_96 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_96);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_96;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_62;
wire n_43;
wire n_82;

BUFx3_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_25),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

INVx8_ASAP7_75t_SL g44 ( 
.A(n_36),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_59),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_0),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_54),
.Y(n_65)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_61),
.Y(n_68)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_45),
.B1(n_47),
.B2(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_55),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_66),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_0),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_59),
.A2(n_43),
.B1(n_48),
.B2(n_51),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_64),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_71),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_75),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g76 ( 
.A(n_72),
.B(n_68),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_76),
.A2(n_46),
.B(n_39),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_67),
.Y(n_77)
);

AO22x1_ASAP7_75t_L g82 ( 
.A1(n_77),
.A2(n_79),
.B1(n_80),
.B2(n_2),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_72),
.A2(n_53),
.B1(n_52),
.B2(n_50),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_4),
.C(n_11),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_82),
.A2(n_74),
.B1(n_6),
.B2(n_8),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_85),
.B(n_86),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_87),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_84),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_83),
.C(n_15),
.Y(n_90)
);

AOI322xp5_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_13),
.A3(n_17),
.B1(n_18),
.B2(n_19),
.C1(n_21),
.C2(n_22),
.Y(n_91)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_23),
.B(n_24),
.Y(n_92)
);

MAJx2_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_26),
.C(n_28),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_29),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_31),
.Y(n_96)
);


endmodule