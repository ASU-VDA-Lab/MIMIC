module fake_jpeg_24803_n_283 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_283);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_283;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_181;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_31),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_19),
.Y(n_44)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_40),
.A2(n_19),
.B1(n_29),
.B2(n_31),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_45),
.B1(n_50),
.B2(n_51),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_29),
.B(n_22),
.C(n_17),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_36),
.B(n_35),
.C(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_33),
.A2(n_19),
.B1(n_29),
.B2(n_17),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_54),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_49),
.B(n_57),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_19),
.B1(n_31),
.B2(n_18),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_33),
.A2(n_18),
.B1(n_22),
.B2(n_24),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_33),
.A2(n_18),
.B1(n_24),
.B2(n_23),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_52),
.A2(n_28),
.B1(n_21),
.B2(n_25),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_20),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_37),
.B(n_18),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_35),
.C(n_36),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_16),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_36),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_32),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_60),
.A2(n_59),
.B(n_84),
.Y(n_112)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_62),
.Y(n_94)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_65),
.Y(n_101)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_66),
.B(n_68),
.Y(n_111)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVxp33_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_16),
.Y(n_73)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_16),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_75),
.Y(n_105)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_43),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_77),
.Y(n_90)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_78),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_79),
.A2(n_41),
.B1(n_42),
.B2(n_21),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_16),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_84),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_55),
.C(n_47),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_35),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_54),
.B(n_38),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_86),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_47),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_96),
.C(n_97),
.Y(n_135)
);

AND2x6_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_55),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_67),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_55),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_104),
.B1(n_107),
.B2(n_77),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_85),
.A2(n_65),
.B1(n_60),
.B2(n_63),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_99),
.A2(n_108),
.B1(n_68),
.B2(n_78),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_45),
.B1(n_51),
.B2(n_52),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_61),
.A2(n_35),
.B1(n_50),
.B2(n_55),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g108 ( 
.A1(n_77),
.A2(n_76),
.B1(n_72),
.B2(n_69),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_113),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_20),
.B(n_32),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_39),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_107),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_115),
.A2(n_116),
.B1(n_132),
.B2(n_90),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_99),
.A2(n_59),
.B1(n_86),
.B2(n_39),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_100),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_117),
.B(n_119),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g118 ( 
.A(n_91),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_125),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_86),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_100),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_120),
.B(n_124),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_64),
.Y(n_121)
);

BUFx24_ASAP7_75t_SL g156 ( 
.A(n_121),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_122),
.B(n_131),
.Y(n_148)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_129),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_113),
.Y(n_127)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_88),
.B(n_82),
.Y(n_128)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_105),
.B(n_82),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_134),
.Y(n_166)
);

XNOR2x1_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_34),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_89),
.A2(n_39),
.B1(n_70),
.B2(n_62),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_66),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_133),
.Y(n_155)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_136),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_16),
.Y(n_137)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_108),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_138),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_112),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_139),
.A2(n_140),
.B(n_87),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_141),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_171),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_145),
.A2(n_161),
.B(n_169),
.Y(n_187)
);

OAI32xp33_ASAP7_75t_L g147 ( 
.A1(n_116),
.A2(n_93),
.A3(n_98),
.B1(n_89),
.B2(n_104),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_164),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_107),
.B1(n_95),
.B2(n_71),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_150),
.A2(n_163),
.B1(n_30),
.B2(n_28),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_106),
.C(n_87),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_151),
.B(n_167),
.C(n_25),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_131),
.Y(n_174)
);

OA21x2_ASAP7_75t_L g157 ( 
.A1(n_115),
.A2(n_107),
.B(n_90),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_157),
.A2(n_140),
.B(n_126),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_159),
.A2(n_162),
.B(n_168),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_139),
.A2(n_106),
.B(n_20),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_123),
.A2(n_14),
.B(n_15),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_114),
.A2(n_103),
.B1(n_34),
.B2(n_90),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_27),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_34),
.C(n_32),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_123),
.A2(n_30),
.B(n_28),
.Y(n_168)
);

AND2x2_ASAP7_75t_SL g169 ( 
.A(n_127),
.B(n_27),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_173),
.A2(n_178),
.B(n_184),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_182),
.Y(n_216)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_181),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_171),
.A2(n_125),
.B1(n_128),
.B2(n_124),
.Y(n_178)
);

INVxp67_ASAP7_75t_SL g179 ( 
.A(n_153),
.Y(n_179)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_179),
.Y(n_198)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_170),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_180),
.B(n_183),
.Y(n_218)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_129),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_164),
.B(n_134),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_157),
.A2(n_136),
.B(n_118),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_164),
.B(n_27),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_185),
.B(n_197),
.Y(n_214)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_193),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_190),
.C(n_167),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_141),
.Y(n_189)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_11),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_149),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_192),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_158),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_163),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_143),
.Y(n_194)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_195),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_196),
.A2(n_146),
.B1(n_153),
.B2(n_30),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_23),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_200),
.Y(n_224)
);

OA21x2_ASAP7_75t_SL g200 ( 
.A1(n_187),
.A2(n_156),
.B(n_145),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_151),
.C(n_144),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_209),
.C(n_193),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_148),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_206),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_190),
.B(n_154),
.Y(n_206)
);

OAI322xp33_ASAP7_75t_L g208 ( 
.A1(n_187),
.A2(n_169),
.A3(n_154),
.B1(n_144),
.B2(n_161),
.C1(n_160),
.C2(n_147),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_210),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_160),
.C(n_150),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_159),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_213),
.A2(n_189),
.B1(n_176),
.B2(n_178),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_177),
.A2(n_146),
.B1(n_25),
.B2(n_21),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_215),
.A2(n_196),
.B1(n_195),
.B2(n_181),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_212),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_218),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_223),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_173),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_230),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

NOR3xp33_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_186),
.C(n_175),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_226),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_203),
.A2(n_176),
.B(n_172),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_231),
.C(n_235),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_203),
.A2(n_184),
.B(n_194),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_233),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_204),
.B(n_194),
.Y(n_230)
);

A2O1A1O1Ixp25_ASAP7_75t_L g231 ( 
.A1(n_210),
.A2(n_8),
.B(n_15),
.C(n_2),
.D(n_3),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_211),
.A2(n_26),
.B1(n_24),
.B2(n_0),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_207),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_234),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_206),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_209),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_8),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_205),
.C(n_216),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_248),
.C(n_227),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_244),
.B(n_245),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_207),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_231),
.A2(n_202),
.B1(n_211),
.B2(n_213),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_246),
.A2(n_26),
.B1(n_7),
.B2(n_3),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_199),
.C(n_215),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_SL g249 ( 
.A(n_237),
.B(n_224),
.C(n_221),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_249),
.A2(n_248),
.B(n_241),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_240),
.A2(n_232),
.B1(n_227),
.B2(n_214),
.Y(n_250)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_247),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_252),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_257),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_242),
.B(n_8),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_256),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_7),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_26),
.C(n_1),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_259),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_0),
.C(n_1),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_263),
.A2(n_11),
.B(n_4),
.Y(n_273)
);

NOR2xp67_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_243),
.Y(n_265)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_265),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_9),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_267),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_9),
.Y(n_267)
);

AOI21x1_ASAP7_75t_L g269 ( 
.A1(n_268),
.A2(n_263),
.B(n_260),
.Y(n_269)
);

AOI322xp5_ASAP7_75t_L g277 ( 
.A1(n_269),
.A2(n_1),
.A3(n_5),
.B1(n_12),
.B2(n_13),
.C1(n_15),
.C2(n_271),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_264),
.A2(n_252),
.B(n_262),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_4),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_0),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_5),
.C(n_13),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_273),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_275),
.Y(n_280)
);

O2A1O1Ixp33_ASAP7_75t_SL g279 ( 
.A1(n_276),
.A2(n_277),
.B(n_278),
.C(n_274),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_279),
.B(n_272),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_280),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_278),
.Y(n_283)
);


endmodule