module real_jpeg_4773_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_173;
wire n_105;
wire n_40;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_244;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_2),
.A2(n_172),
.B1(n_173),
.B2(n_176),
.Y(n_171)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_2),
.Y(n_176)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_4),
.Y(n_178)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_4),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_4),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_5),
.A2(n_96),
.B1(n_99),
.B2(n_100),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_5),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_5),
.A2(n_99),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_5),
.A2(n_25),
.B1(n_99),
.B2(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_6),
.B(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_6),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_6),
.A2(n_129),
.B1(n_188),
.B2(n_191),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_6),
.B(n_86),
.C(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_6),
.B(n_120),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_6),
.B(n_34),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_6),
.B(n_145),
.Y(n_232)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_8),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_9),
.A2(n_55),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_9),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_9),
.A2(n_105),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_10),
.Y(n_163)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_10),
.Y(n_169)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_11),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_11),
.Y(n_86)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_11),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_12),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_12),
.A2(n_43),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_12),
.A2(n_43),
.B1(n_122),
.B2(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_182),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_180),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_136),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_16),
.B(n_136),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_74),
.C(n_106),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_17),
.B(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_49),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_18),
.B(n_49),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_30),
.B(n_32),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_20),
.A2(n_33),
.B1(n_171),
.B2(n_177),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_21),
.Y(n_202)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

BUFx8_ASAP7_75t_L g175 ( 
.A(n_23),
.Y(n_175)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_23),
.Y(n_206)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_30),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_32),
.A2(n_226),
.B(n_229),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_38),
.Y(n_32)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_33),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_33),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_38),
.B(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_40),
.Y(n_172)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_42),
.Y(n_228)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_48),
.Y(n_198)
);

AOI32xp33_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_55),
.A3(n_59),
.B1(n_64),
.B2(n_66),
.Y(n_49)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_50),
.Y(n_133)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_53),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_54),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_54),
.Y(n_155)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_58),
.Y(n_144)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_58),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

INVxp33_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

NAND2xp33_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_74),
.A2(n_106),
.B1(n_107),
.B2(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_74),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_88),
.B1(n_95),
.B2(n_103),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_75),
.A2(n_103),
.B(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_75),
.A2(n_140),
.B(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_76),
.B(n_141),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_88),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_82),
.B1(n_85),
.B2(n_87),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_81),
.Y(n_190)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22x1_ASAP7_75t_L g88 ( 
.A1(n_85),
.A2(n_89),
.B1(n_92),
.B2(n_94),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_88),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_88),
.A2(n_95),
.B(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AO22x2_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_120)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_98),
.Y(n_195)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_125),
.B(n_131),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_108),
.B(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_109),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_120),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_113),
.B1(n_116),
.B2(n_118),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_115),
.Y(n_166)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_120),
.Y(n_135)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_129),
.B(n_130),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_160),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_129),
.A2(n_207),
.B(n_208),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.Y(n_131)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_135),
.A2(n_149),
.B(n_156),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_147),
.B2(n_179),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_146),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_145),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_158),
.Y(n_147)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_170),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.Y(n_162)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_173),
.B(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_244),
.B(n_249),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_218),
.B(n_243),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_199),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_185),
.B(n_199),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_193),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_186),
.A2(n_193),
.B1(n_194),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_186),
.Y(n_241)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_212),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_200),
.B(n_213),
.C(n_217),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_207),
.B(n_208),
.Y(n_200)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_201),
.Y(n_237)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_216),
.B2(n_217),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_234),
.B(n_242),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_224),
.B(n_233),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_232),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_232),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_240),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_240),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_246),
.Y(n_249)
);


endmodule