module fake_jpeg_1126_n_116 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_116);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_116;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_0),
.Y(n_41)
);

XNOR2x1_ASAP7_75t_SL g49 ( 
.A(n_41),
.B(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_35),
.B1(n_31),
.B2(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_31),
.Y(n_54)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

BUFx4f_ASAP7_75t_SL g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_30),
.Y(n_66)
);

OR2x2_ASAP7_75t_SL g58 ( 
.A(n_49),
.B(n_39),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_32),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_44),
.B1(n_46),
.B2(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_57),
.B(n_60),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_58),
.B(n_59),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_40),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_39),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_54),
.A2(n_43),
.B1(n_42),
.B2(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_55),
.Y(n_73)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_48),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_30),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_65),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_73),
.B1(n_74),
.B2(n_4),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_72),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_0),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_1),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_1),
.Y(n_88)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

XNOR2x2_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_53),
.Y(n_79)
);

OA21x2_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_87),
.B(n_6),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_13),
.C(n_27),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_85),
.C(n_16),
.Y(n_96)
);

NOR3xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_36),
.C(n_2),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_88),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_12),
.C(n_24),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_2),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_68),
.B(n_10),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_36),
.B(n_3),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_89),
.A2(n_6),
.B(n_8),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_90),
.Y(n_95)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_83),
.B(n_5),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_94),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_5),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_100),
.C(n_87),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_99),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_8),
.B1(n_9),
.B2(n_14),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_91),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_104),
.Y(n_108)
);

BUFx12_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_105),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_102),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_105),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_111),
.B(n_94),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_112),
.A2(n_95),
.B1(n_92),
.B2(n_103),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_101),
.Y(n_114)
);

OAI221xp5_ASAP7_75t_SL g115 ( 
.A1(n_114),
.A2(n_107),
.B1(n_18),
.B2(n_21),
.C(n_22),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_17),
.Y(n_116)
);


endmodule