module fake_netlist_6_3551_n_1800 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1800);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1800;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g175 ( 
.A(n_118),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_49),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_100),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_165),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_135),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_46),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_79),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_98),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_37),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_54),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_78),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_8),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_80),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_73),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_15),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_107),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_71),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_113),
.Y(n_192)
);

BUFx8_ASAP7_75t_SL g193 ( 
.A(n_126),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_88),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_138),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_152),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_61),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_128),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_38),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_0),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_54),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_38),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_57),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_106),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_45),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_154),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_83),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_133),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_2),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_87),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_119),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_155),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_21),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_36),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_10),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_123),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_41),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_72),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_27),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_170),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_150),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_140),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_142),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_168),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_17),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_15),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_51),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_21),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_85),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_51),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_163),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_162),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_112),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_37),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_33),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_147),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_90),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_49),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_82),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_164),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_36),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_45),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_159),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_50),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_5),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_47),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_13),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_161),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_59),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_25),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_109),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_114),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_120),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_13),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_158),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_144),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_75),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_166),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_69),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_39),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_34),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_17),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_2),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_104),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_93),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_137),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_34),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_4),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_141),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_130),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_22),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_44),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_103),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_84),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_116),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_148),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_139),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_32),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_121),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_67),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_127),
.Y(n_282)
);

BUFx8_ASAP7_75t_SL g283 ( 
.A(n_43),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_89),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_95),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_172),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_97),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_33),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_20),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_3),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_23),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_50),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_102),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_25),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_92),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_3),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_8),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_96),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_160),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_65),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_76),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_134),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_31),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_18),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_117),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_157),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_47),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_20),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_64),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_31),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_77),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_108),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_115),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_48),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_173),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_145),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_146),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_16),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_129),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_23),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_6),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_125),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_111),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_63),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_74),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_153),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_156),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_16),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_171),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_27),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_4),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_52),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_99),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_110),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_58),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_28),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_62),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_18),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_131),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_122),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_70),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_132),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_5),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_1),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_101),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_53),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_7),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_66),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_0),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_22),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_52),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_86),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_193),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_283),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_178),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_179),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_242),
.Y(n_357)
);

INVxp33_ASAP7_75t_L g358 ( 
.A(n_176),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_305),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_213),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_352),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_221),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_239),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_239),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_230),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_352),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_239),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_180),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_239),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_184),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_181),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_239),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_182),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_257),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_289),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_316),
.Y(n_376)
);

NOR2xp67_ASAP7_75t_L g377 ( 
.A(n_207),
.B(n_1),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_188),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_317),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_319),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_327),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_289),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_191),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_186),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_209),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_289),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_289),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_211),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_176),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_333),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_289),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_211),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_183),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_183),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_189),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_192),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_209),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_229),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_249),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_196),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_198),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_341),
.Y(n_402)
);

INVxp67_ASAP7_75t_SL g403 ( 
.A(n_329),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_211),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_229),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_345),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_292),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_292),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_216),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_201),
.Y(n_410)
);

CKINVDCx14_ASAP7_75t_R g411 ( 
.A(n_185),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_249),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_200),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_204),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_201),
.Y(n_415)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_329),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_203),
.Y(n_417)
);

INVxp33_ASAP7_75t_SL g418 ( 
.A(n_215),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_203),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_175),
.B(n_6),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_207),
.B(n_7),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_206),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_206),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_205),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_208),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_210),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_211),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_210),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_212),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_214),
.B(n_9),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_214),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_231),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_334),
.Y(n_433)
);

INVxp67_ASAP7_75t_SL g434 ( 
.A(n_194),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_216),
.B(n_9),
.Y(n_435)
);

INVxp67_ASAP7_75t_SL g436 ( 
.A(n_194),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_219),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_334),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_175),
.B(n_10),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_231),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_262),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_363),
.Y(n_442)
);

INVx2_ASAP7_75t_SL g443 ( 
.A(n_409),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_409),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_363),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_364),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_355),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_364),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_388),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_388),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_367),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_367),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_369),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_360),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_435),
.B(n_207),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_357),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_356),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_362),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_388),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_392),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_369),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_377),
.B(n_197),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_368),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_392),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_392),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_365),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_371),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_404),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_372),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_404),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_404),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_434),
.B(n_223),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_373),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_427),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_427),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_372),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_370),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_427),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_374),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_375),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_375),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_382),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_382),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_386),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_378),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_383),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_421),
.B(n_195),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_386),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_384),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_387),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_436),
.B(n_225),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_396),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_387),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_391),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_400),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_391),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_410),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_401),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_393),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_414),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_377),
.B(n_232),
.Y(n_501)
);

CKINVDCx8_ASAP7_75t_R g502 ( 
.A(n_361),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_376),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_393),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_394),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_394),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_410),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_420),
.B(n_237),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_439),
.B(n_244),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_435),
.B(n_197),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_424),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_415),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_425),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_415),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_398),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_429),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_437),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_353),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_385),
.B(n_293),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_487),
.B(n_501),
.Y(n_520)
);

NAND2xp33_ASAP7_75t_L g521 ( 
.A(n_508),
.B(n_211),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_487),
.B(n_411),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_447),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_501),
.B(n_418),
.Y(n_524)
);

BUFx4f_ASAP7_75t_L g525 ( 
.A(n_443),
.Y(n_525)
);

INVx1_ASAP7_75t_SL g526 ( 
.A(n_456),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_476),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_476),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_455),
.A2(n_430),
.B1(n_226),
.B2(n_350),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_455),
.A2(n_430),
.B1(n_226),
.B2(n_272),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_490),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_497),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_456),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_462),
.B(n_361),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_444),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_490),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_497),
.Y(n_537)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_462),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_490),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_484),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_443),
.B(n_366),
.Y(n_541)
);

AND2x6_ASAP7_75t_L g542 ( 
.A(n_455),
.B(n_177),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_462),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_508),
.B(n_397),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_462),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_507),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_507),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_490),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_484),
.Y(n_549)
);

OR2x2_ASAP7_75t_L g550 ( 
.A(n_443),
.B(n_366),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_512),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_509),
.B(n_403),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_512),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_484),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_514),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_462),
.B(n_399),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_444),
.Y(n_557)
);

AND2x6_ASAP7_75t_L g558 ( 
.A(n_510),
.B(n_177),
.Y(n_558)
);

BUFx4f_ASAP7_75t_L g559 ( 
.A(n_514),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_519),
.B(n_399),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_510),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_494),
.Y(n_562)
);

INVx4_ASAP7_75t_L g563 ( 
.A(n_480),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_480),
.Y(n_564)
);

AND2x2_ASAP7_75t_SL g565 ( 
.A(n_509),
.B(n_433),
.Y(n_565)
);

OAI22xp33_ASAP7_75t_L g566 ( 
.A1(n_519),
.A2(n_433),
.B1(n_416),
.B2(n_359),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_472),
.B(n_491),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_442),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_472),
.B(n_395),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_449),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_494),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_491),
.B(n_413),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_463),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_463),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_494),
.Y(n_575)
);

NAND2xp33_ASAP7_75t_L g576 ( 
.A(n_510),
.B(n_306),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_477),
.B(n_358),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_442),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_477),
.B(n_389),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_490),
.B(n_224),
.Y(n_580)
);

INVx1_ASAP7_75t_SL g581 ( 
.A(n_454),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_445),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_499),
.A2(n_349),
.B1(n_288),
.B2(n_330),
.Y(n_583)
);

INVx5_ASAP7_75t_L g584 ( 
.A(n_480),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_489),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_445),
.B(n_224),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_449),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_496),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_496),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_489),
.Y(n_590)
);

OR2x2_ASAP7_75t_L g591 ( 
.A(n_457),
.B(n_432),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_458),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_467),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_449),
.Y(n_594)
);

INVxp67_ASAP7_75t_SL g595 ( 
.A(n_449),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_480),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_473),
.B(n_217),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_L g598 ( 
.A(n_485),
.B(n_306),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_486),
.B(n_311),
.Y(n_599)
);

INVx1_ASAP7_75t_SL g600 ( 
.A(n_466),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_492),
.B(n_217),
.Y(n_601)
);

INVx5_ASAP7_75t_L g602 ( 
.A(n_480),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_446),
.B(n_233),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_446),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_448),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_495),
.B(n_340),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_498),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_500),
.B(n_266),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_511),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_513),
.B(n_266),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_516),
.B(n_417),
.Y(n_611)
);

BUFx8_ASAP7_75t_SL g612 ( 
.A(n_479),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_517),
.B(n_282),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_448),
.B(n_233),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_499),
.A2(n_308),
.B1(n_279),
.B2(n_288),
.Y(n_615)
);

AND2x6_ASAP7_75t_L g616 ( 
.A(n_451),
.B(n_187),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_499),
.B(n_315),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_451),
.Y(n_618)
);

AND2x6_ASAP7_75t_L g619 ( 
.A(n_452),
.B(n_187),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_499),
.B(n_315),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_502),
.B(n_354),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_502),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_502),
.B(n_412),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_452),
.B(n_417),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_453),
.B(n_419),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_449),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_505),
.B(n_348),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_453),
.Y(n_628)
);

AND2x2_ASAP7_75t_SL g629 ( 
.A(n_506),
.B(n_282),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_461),
.B(n_419),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_461),
.Y(n_631)
);

OAI22xp33_ASAP7_75t_L g632 ( 
.A1(n_518),
.A2(n_303),
.B1(n_202),
.B2(n_235),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_469),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_469),
.B(n_348),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_505),
.B(n_306),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_481),
.B(n_422),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_505),
.B(n_306),
.Y(n_637)
);

INVx4_ASAP7_75t_L g638 ( 
.A(n_480),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_482),
.B(n_422),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_496),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_482),
.B(n_252),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_488),
.B(n_254),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_449),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_488),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_505),
.B(n_423),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_503),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_480),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_483),
.B(n_258),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_515),
.B(n_306),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_483),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_459),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_483),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_515),
.B(n_438),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_506),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_459),
.Y(n_655)
);

INVx5_ASAP7_75t_L g656 ( 
.A(n_483),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_515),
.B(n_423),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_515),
.A2(n_272),
.B1(n_351),
.B2(n_350),
.Y(n_658)
);

INVx6_ASAP7_75t_L g659 ( 
.A(n_483),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_504),
.B(n_190),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_504),
.B(n_190),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_504),
.A2(n_308),
.B1(n_296),
.B2(n_279),
.Y(n_662)
);

BUFx2_ASAP7_75t_L g663 ( 
.A(n_504),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_504),
.B(n_426),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_483),
.Y(n_665)
);

NAND2xp33_ASAP7_75t_L g666 ( 
.A(n_449),
.B(n_259),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_506),
.A2(n_406),
.B1(n_402),
.B2(n_390),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_474),
.B(n_441),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_459),
.A2(n_296),
.B1(n_262),
.B2(n_351),
.Y(n_669)
);

BUFx10_ASAP7_75t_L g670 ( 
.A(n_483),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_520),
.B(n_269),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_567),
.B(n_493),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_529),
.A2(n_330),
.B1(n_331),
.B2(n_344),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_525),
.B(n_379),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_525),
.B(n_380),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_544),
.B(n_552),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_544),
.B(n_493),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_545),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_552),
.B(n_218),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_612),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_561),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_545),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_654),
.B(n_493),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_565),
.A2(n_381),
.B1(n_275),
.B2(n_281),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_651),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_533),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_527),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_663),
.Y(n_688)
);

INVx4_ASAP7_75t_L g689 ( 
.A(n_528),
.Y(n_689)
);

AO221x1_ASAP7_75t_L g690 ( 
.A1(n_566),
.A2(n_331),
.B1(n_344),
.B2(n_349),
.C(n_222),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_540),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_528),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_531),
.B(n_493),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_531),
.B(n_493),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_532),
.B(n_426),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_569),
.B(n_220),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_565),
.A2(n_560),
.B1(n_524),
.B2(n_556),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_537),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_611),
.B(n_526),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_577),
.B(n_263),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_529),
.A2(n_530),
.B1(n_662),
.B2(n_542),
.Y(n_701)
);

A2O1A1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_559),
.A2(n_302),
.B(n_287),
.C(n_285),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_534),
.A2(n_271),
.B1(n_276),
.B2(n_274),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_530),
.A2(n_240),
.B1(n_277),
.B2(n_278),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_611),
.B(n_265),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_536),
.B(n_493),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_539),
.B(n_199),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_572),
.B(n_267),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_539),
.B(n_199),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_549),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_546),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_559),
.B(n_284),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_528),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_548),
.B(n_222),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_599),
.B(n_227),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_548),
.B(n_234),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_662),
.A2(n_238),
.B1(n_287),
.B2(n_285),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_528),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_547),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_534),
.A2(n_309),
.B1(n_300),
.B2(n_299),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_629),
.B(n_234),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_629),
.B(n_238),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_551),
.Y(n_723)
);

BUFx5_ASAP7_75t_L g724 ( 
.A(n_670),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_549),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_542),
.A2(n_302),
.B1(n_256),
.B2(n_253),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_553),
.B(n_240),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_599),
.B(n_228),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_555),
.B(n_568),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_606),
.B(n_286),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_535),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_554),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_554),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_556),
.A2(n_295),
.B1(n_325),
.B2(n_335),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_606),
.B(n_236),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_592),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_578),
.B(n_241),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_523),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_558),
.A2(n_326),
.B1(n_322),
.B2(n_313),
.Y(n_739)
);

NOR2xp67_ASAP7_75t_L g740 ( 
.A(n_593),
.B(n_298),
.Y(n_740)
);

NAND2x1_ASAP7_75t_L g741 ( 
.A(n_538),
.B(n_474),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_579),
.B(n_243),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_582),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_562),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_604),
.B(n_241),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_605),
.B(n_250),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_562),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_571),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_618),
.B(n_250),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_651),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_628),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_541),
.B(n_550),
.Y(n_752)
);

NAND3xp33_ASAP7_75t_L g753 ( 
.A(n_597),
.B(n_264),
.C(n_268),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_522),
.B(n_597),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_538),
.A2(n_260),
.B1(n_256),
.B2(n_253),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_543),
.A2(n_280),
.B1(n_278),
.B2(n_277),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_571),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_575),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_601),
.B(n_608),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_573),
.Y(n_760)
);

INVxp67_ASAP7_75t_L g761 ( 
.A(n_574),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_591),
.B(n_301),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_631),
.B(n_260),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_575),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_542),
.A2(n_583),
.B1(n_658),
.B2(n_615),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_633),
.B(n_280),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_655),
.Y(n_767)
);

A2O1A1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_664),
.A2(n_323),
.B(n_342),
.C(n_324),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_644),
.B(n_323),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_542),
.B(n_342),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_653),
.Y(n_771)
);

INVxp67_ASAP7_75t_SL g772 ( 
.A(n_570),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_543),
.B(n_474),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_558),
.B(n_474),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_588),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_588),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_589),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_601),
.B(n_312),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_583),
.A2(n_263),
.B1(n_346),
.B2(n_291),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_589),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_655),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_558),
.B(n_450),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_558),
.B(n_450),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_585),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_558),
.B(n_450),
.Y(n_785)
);

NAND2xp33_ASAP7_75t_L g786 ( 
.A(n_616),
.B(n_337),
.Y(n_786)
);

AOI221xp5_ASAP7_75t_L g787 ( 
.A1(n_632),
.A2(n_307),
.B1(n_336),
.B2(n_321),
.C(n_320),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_570),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_668),
.Y(n_789)
);

OAI22xp33_ASAP7_75t_L g790 ( 
.A1(n_557),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_617),
.B(n_450),
.Y(n_791)
);

CKINVDCx20_ASAP7_75t_R g792 ( 
.A(n_607),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_640),
.Y(n_793)
);

AND2x4_ASAP7_75t_L g794 ( 
.A(n_627),
.B(n_428),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_627),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_615),
.A2(n_428),
.B1(n_431),
.B2(n_440),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_648),
.A2(n_478),
.B(n_475),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_640),
.Y(n_798)
);

OAI221xp5_ASAP7_75t_L g799 ( 
.A1(n_658),
.A2(n_431),
.B1(n_440),
.B2(n_441),
.C(n_261),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_617),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_617),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_608),
.B(n_339),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_610),
.B(n_270),
.Y(n_803)
);

OAI22xp5_ASAP7_75t_SL g804 ( 
.A1(n_581),
.A2(n_314),
.B1(n_255),
.B2(n_251),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_620),
.B(n_450),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_610),
.B(n_270),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_616),
.A2(n_270),
.B1(n_248),
.B2(n_338),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_620),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_616),
.A2(n_619),
.B1(n_669),
.B2(n_664),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_620),
.B(n_460),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_590),
.B(n_398),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_645),
.B(n_460),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_613),
.B(n_270),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_645),
.B(n_460),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_600),
.Y(n_815)
);

AO221x1_ASAP7_75t_L g816 ( 
.A1(n_570),
.A2(n_405),
.B1(n_407),
.B2(n_408),
.C(n_468),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_667),
.B(n_646),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_657),
.B(n_460),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_659),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_SL g820 ( 
.A(n_609),
.B(n_343),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_586),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_641),
.B(n_464),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_595),
.A2(n_465),
.B(n_475),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_642),
.B(n_464),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_613),
.B(n_347),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_598),
.B(n_273),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_622),
.B(n_290),
.Y(n_827)
);

NOR3xp33_ASAP7_75t_L g828 ( 
.A(n_623),
.B(n_294),
.C(n_297),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_603),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_580),
.B(n_464),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_521),
.B(n_464),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_614),
.B(n_304),
.Y(n_832)
);

AO22x1_ASAP7_75t_L g833 ( 
.A1(n_616),
.A2(n_310),
.B1(n_318),
.B2(n_328),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_576),
.B(n_468),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_616),
.B(n_468),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_634),
.B(n_332),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_676),
.B(n_621),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_682),
.Y(n_838)
);

O2A1O1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_676),
.A2(n_660),
.B(n_661),
.C(n_649),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_672),
.A2(n_635),
.B(n_637),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_679),
.B(n_624),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_754),
.A2(n_679),
.B1(n_759),
.B2(n_728),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_681),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_701),
.A2(n_669),
.B1(n_661),
.B2(n_660),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_701),
.A2(n_635),
.B1(n_637),
.B2(n_649),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_691),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_682),
.Y(n_847)
);

NAND2x1p5_ASAP7_75t_L g848 ( 
.A(n_678),
.B(n_563),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_715),
.B(n_624),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_677),
.A2(n_666),
.B(n_647),
.Y(n_850)
);

OAI21xp5_ASAP7_75t_L g851 ( 
.A1(n_721),
.A2(n_652),
.B(n_665),
.Y(n_851)
);

AO22x1_ASAP7_75t_L g852 ( 
.A1(n_728),
.A2(n_619),
.B1(n_625),
.B2(n_630),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_722),
.A2(n_650),
.B(n_619),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_671),
.B(n_630),
.Y(n_854)
);

BUFx8_ASAP7_75t_L g855 ( 
.A(n_686),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_688),
.B(n_405),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_671),
.B(n_636),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_742),
.B(n_811),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_800),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_735),
.B(n_636),
.Y(n_860)
);

CKINVDCx10_ASAP7_75t_R g861 ( 
.A(n_680),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_735),
.B(n_639),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_754),
.B(n_639),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_L g864 ( 
.A1(n_812),
.A2(n_619),
.B(n_564),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_742),
.B(n_407),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_682),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_821),
.B(n_594),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_682),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_759),
.A2(n_659),
.B1(n_596),
.B2(n_563),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_808),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_765),
.A2(n_659),
.B1(n_594),
.B2(n_643),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_829),
.B(n_594),
.Y(n_872)
);

AOI21x1_ASAP7_75t_L g873 ( 
.A1(n_741),
.A2(n_773),
.B(n_709),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_696),
.B(n_594),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_791),
.A2(n_564),
.B(n_638),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_814),
.A2(n_638),
.B(n_596),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_696),
.B(n_570),
.Y(n_877)
);

AOI21x1_ASAP7_75t_L g878 ( 
.A1(n_707),
.A2(n_478),
.B(n_465),
.Y(n_878)
);

A2O1A1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_765),
.A2(n_408),
.B(n_465),
.C(n_478),
.Y(n_879)
);

OAI21xp33_ASAP7_75t_L g880 ( 
.A1(n_779),
.A2(n_470),
.B(n_471),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_789),
.B(n_587),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_738),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_697),
.B(n_587),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_805),
.A2(n_587),
.B(n_626),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_698),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_801),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_690),
.A2(n_587),
.B1(n_643),
.B2(n_626),
.Y(n_887)
);

CKINVDCx14_ASAP7_75t_R g888 ( 
.A(n_792),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_832),
.B(n_836),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_711),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_832),
.B(n_643),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_810),
.A2(n_626),
.B(n_656),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_836),
.B(n_626),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_699),
.B(n_11),
.Y(n_894)
);

OAI321xp33_ASAP7_75t_L g895 ( 
.A1(n_807),
.A2(n_11),
.A3(n_12),
.B1(n_14),
.B2(n_19),
.C(n_24),
.Y(n_895)
);

NAND2x1p5_ASAP7_75t_L g896 ( 
.A(n_801),
.B(n_689),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_719),
.B(n_475),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_723),
.B(n_471),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_830),
.A2(n_656),
.B(n_602),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_743),
.B(n_471),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_731),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_710),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_693),
.A2(n_656),
.B(n_602),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_752),
.B(n_14),
.Y(n_904)
);

OAI22xp5_ASAP7_75t_L g905 ( 
.A1(n_809),
.A2(n_470),
.B1(n_468),
.B2(n_602),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_752),
.B(n_19),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_809),
.A2(n_470),
.B1(n_468),
.B2(n_602),
.Y(n_907)
);

O2A1O1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_768),
.A2(n_24),
.B(n_26),
.C(n_28),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_751),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_694),
.A2(n_656),
.B(n_584),
.Y(n_910)
);

NOR3xp33_ASAP7_75t_L g911 ( 
.A(n_787),
.B(n_26),
.C(n_29),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_706),
.A2(n_584),
.B(n_468),
.Y(n_912)
);

OAI22xp33_ASAP7_75t_L g913 ( 
.A1(n_729),
.A2(n_468),
.B1(n_584),
.B2(n_32),
.Y(n_913)
);

INVx2_ASAP7_75t_SL g914 ( 
.A(n_700),
.Y(n_914)
);

BUFx12f_ASAP7_75t_L g915 ( 
.A(n_736),
.Y(n_915)
);

NAND3xp33_ASAP7_75t_L g916 ( 
.A(n_779),
.B(n_29),
.C(n_30),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_794),
.B(n_30),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_771),
.A2(n_68),
.B1(n_169),
.B2(n_167),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_822),
.A2(n_824),
.B(n_683),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_826),
.A2(n_35),
.B(n_39),
.C(n_40),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_687),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_760),
.B(n_35),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_794),
.B(n_40),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_818),
.A2(n_772),
.B(n_714),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_704),
.B(n_41),
.Y(n_925)
);

INVx8_ASAP7_75t_L g926 ( 
.A(n_695),
.Y(n_926)
);

NOR3xp33_ASAP7_75t_L g927 ( 
.A(n_804),
.B(n_42),
.C(n_44),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_716),
.A2(n_91),
.B(n_149),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_770),
.A2(n_81),
.B(n_143),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_704),
.B(n_46),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_774),
.A2(n_94),
.B(n_136),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_695),
.B(n_48),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_726),
.A2(n_60),
.B1(n_105),
.B2(n_124),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_SL g934 ( 
.A(n_815),
.B(n_174),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_788),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_820),
.B(n_53),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_782),
.A2(n_55),
.B(n_56),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_725),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_732),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_736),
.Y(n_940)
);

NAND3xp33_ASAP7_75t_L g941 ( 
.A(n_807),
.B(n_55),
.C(n_56),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_795),
.A2(n_828),
.B1(n_826),
.B2(n_730),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_761),
.B(n_724),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_783),
.A2(n_785),
.B(n_835),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_784),
.B(n_705),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_817),
.B(n_708),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_726),
.B(n_724),
.Y(n_947)
);

CKINVDCx20_ASAP7_75t_R g948 ( 
.A(n_674),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_753),
.A2(n_673),
.B(n_684),
.C(n_717),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_724),
.B(n_763),
.Y(n_950)
);

NOR2x1_ASAP7_75t_L g951 ( 
.A(n_740),
.B(n_675),
.Y(n_951)
);

AOI21x1_ASAP7_75t_L g952 ( 
.A1(n_834),
.A2(n_823),
.B(n_797),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_831),
.A2(n_758),
.B(n_798),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_827),
.B(n_762),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_724),
.B(n_766),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_673),
.B(n_825),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_724),
.B(n_769),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_732),
.A2(n_780),
.B(n_764),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_717),
.A2(n_737),
.B(n_727),
.C(n_745),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_733),
.A2(n_764),
.B(n_798),
.Y(n_960)
);

INVx2_ASAP7_75t_SL g961 ( 
.A(n_746),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_733),
.A2(n_758),
.B(n_793),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_744),
.A2(n_793),
.B(n_780),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_755),
.A2(n_756),
.B(n_749),
.C(n_702),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_724),
.B(n_713),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_803),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_744),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_747),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_747),
.A2(n_776),
.B(n_777),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_806),
.B(n_813),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_748),
.A2(n_775),
.B(n_777),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_718),
.A2(n_689),
.B1(n_739),
.B2(n_692),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_778),
.B(n_802),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_748),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_692),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_692),
.B(n_713),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_757),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_713),
.B(n_776),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_757),
.B(n_775),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_685),
.B(n_750),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_767),
.A2(n_781),
.B(n_786),
.Y(n_981)
);

O2A1O1Ixp5_ASAP7_75t_L g982 ( 
.A1(n_712),
.A2(n_819),
.B(n_833),
.C(n_790),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_788),
.A2(n_819),
.B(n_816),
.Y(n_983)
);

AOI22xp5_ASAP7_75t_L g984 ( 
.A1(n_703),
.A2(n_720),
.B1(n_734),
.B2(n_788),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_796),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_799),
.A2(n_676),
.B(n_679),
.C(n_715),
.Y(n_986)
);

AOI21x1_ASAP7_75t_L g987 ( 
.A1(n_796),
.A2(n_741),
.B(n_773),
.Y(n_987)
);

BUFx12f_ASAP7_75t_L g988 ( 
.A(n_738),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_691),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_676),
.B(n_567),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_681),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_676),
.B(n_526),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_676),
.B(n_526),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_676),
.B(n_526),
.Y(n_994)
);

INVx1_ASAP7_75t_SL g995 ( 
.A(n_686),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_672),
.A2(n_677),
.B(n_791),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_738),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_SL g998 ( 
.A1(n_792),
.A2(n_362),
.B1(n_365),
.B2(n_360),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_681),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_676),
.B(n_526),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_676),
.B(n_567),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_672),
.A2(n_677),
.B(n_791),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_672),
.A2(n_677),
.B(n_791),
.Y(n_1003)
);

AOI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_676),
.A2(n_754),
.B1(n_679),
.B2(n_759),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_676),
.B(n_526),
.Y(n_1005)
);

NOR2x1_ASAP7_75t_L g1006 ( 
.A(n_699),
.B(n_526),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_672),
.A2(n_677),
.B(n_791),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_676),
.B(n_567),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_676),
.B(n_567),
.Y(n_1009)
);

BUFx2_ASAP7_75t_L g1010 ( 
.A(n_686),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_672),
.A2(n_677),
.B(n_791),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_676),
.A2(n_701),
.B1(n_765),
.B2(n_679),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_672),
.A2(n_677),
.B(n_791),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_950),
.A2(n_957),
.B(n_955),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_L g1015 ( 
.A1(n_952),
.A2(n_884),
.B(n_981),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_842),
.A2(n_849),
.B(n_1004),
.C(n_986),
.Y(n_1016)
);

AO22x2_ASAP7_75t_L g1017 ( 
.A1(n_1012),
.A2(n_916),
.B1(n_941),
.B2(n_911),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_992),
.B(n_858),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_885),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_919),
.A2(n_1002),
.B(n_996),
.Y(n_1020)
);

OAI22x1_ASAP7_75t_L g1021 ( 
.A1(n_837),
.A2(n_894),
.B1(n_906),
.B2(n_946),
.Y(n_1021)
);

OR2x6_ASAP7_75t_L g1022 ( 
.A(n_915),
.B(n_926),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_990),
.A2(n_1009),
.B1(n_1001),
.B2(n_1008),
.Y(n_1023)
);

AOI21x1_ASAP7_75t_L g1024 ( 
.A1(n_874),
.A2(n_877),
.B(n_883),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_884),
.A2(n_981),
.B(n_878),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_953),
.A2(n_944),
.B(n_958),
.Y(n_1026)
);

INVxp67_ASAP7_75t_L g1027 ( 
.A(n_1010),
.Y(n_1027)
);

AOI221xp5_ASAP7_75t_SL g1028 ( 
.A1(n_949),
.A2(n_841),
.B1(n_860),
.B2(n_862),
.C(n_857),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_953),
.A2(n_944),
.B(n_958),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_993),
.B(n_994),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_863),
.B(n_854),
.Y(n_1031)
);

HB1xp67_ASAP7_75t_L g1032 ( 
.A(n_901),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_889),
.B(n_865),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_996),
.A2(n_1003),
.B(n_1002),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_1003),
.A2(n_1011),
.B(n_1007),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_1007),
.A2(n_1013),
.B(n_1011),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1000),
.B(n_1005),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_960),
.A2(n_963),
.B(n_962),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_985),
.A2(n_844),
.B1(n_925),
.B2(n_930),
.Y(n_1039)
);

XNOR2xp5_ASAP7_75t_SL g1040 ( 
.A(n_998),
.B(n_882),
.Y(n_1040)
);

INVxp67_ASAP7_75t_SL g1041 ( 
.A(n_838),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_1013),
.A2(n_924),
.B(n_893),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_985),
.B(n_956),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_891),
.A2(n_965),
.B(n_876),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_856),
.B(n_940),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_961),
.B(n_904),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_969),
.A2(n_971),
.B(n_875),
.Y(n_1047)
);

AO21x2_ASAP7_75t_L g1048 ( 
.A1(n_851),
.A2(n_983),
.B(n_864),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_947),
.A2(n_972),
.B(n_853),
.Y(n_1049)
);

AOI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_954),
.A2(n_945),
.B1(n_970),
.B2(n_948),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_984),
.A2(n_845),
.B1(n_959),
.B2(n_890),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_909),
.B(n_921),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_976),
.A2(n_871),
.B(n_839),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_995),
.B(n_914),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_859),
.A2(n_870),
.B1(n_936),
.B2(n_932),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_838),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_840),
.A2(n_850),
.B(n_978),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_L g1058 ( 
.A1(n_892),
.A2(n_873),
.B(n_912),
.Y(n_1058)
);

AOI21x1_ASAP7_75t_L g1059 ( 
.A1(n_983),
.A2(n_850),
.B(n_852),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_942),
.B(n_843),
.Y(n_1060)
);

OA22x2_ASAP7_75t_L g1061 ( 
.A1(n_966),
.A2(n_856),
.B1(n_991),
.B2(n_999),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_892),
.A2(n_899),
.B(n_840),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_867),
.A2(n_872),
.B(n_848),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_879),
.A2(n_982),
.B(n_979),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_855),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_964),
.A2(n_973),
.B(n_929),
.C(n_917),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_899),
.A2(n_987),
.B(n_903),
.Y(n_1067)
);

OAI21xp5_ASAP7_75t_SL g1068 ( 
.A1(n_927),
.A2(n_1006),
.B(n_922),
.Y(n_1068)
);

OAI21xp33_ASAP7_75t_L g1069 ( 
.A1(n_923),
.A2(n_997),
.B(n_934),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_905),
.A2(n_907),
.B(n_939),
.Y(n_1070)
);

OAI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_938),
.A2(n_880),
.B(n_846),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_848),
.A2(n_881),
.B(n_943),
.Y(n_1072)
);

INVx2_ASAP7_75t_SL g1073 ( 
.A(n_855),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_847),
.B(n_868),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_847),
.B(n_868),
.Y(n_1075)
);

NAND2x1_ASAP7_75t_L g1076 ( 
.A(n_886),
.B(n_935),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_951),
.A2(n_895),
.B(n_920),
.C(n_886),
.Y(n_1077)
);

BUFx4_ASAP7_75t_SL g1078 ( 
.A(n_861),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_910),
.A2(n_896),
.B(n_989),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_869),
.A2(n_980),
.B(n_896),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_888),
.B(n_926),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_838),
.B(n_866),
.Y(n_1082)
);

AO31x2_ASAP7_75t_L g1083 ( 
.A1(n_937),
.A2(n_931),
.A3(n_928),
.B(n_933),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_902),
.A2(n_967),
.B(n_974),
.Y(n_1084)
);

NOR2xp67_ASAP7_75t_L g1085 ( 
.A(n_988),
.B(n_937),
.Y(n_1085)
);

OAI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_968),
.A2(n_977),
.B(n_887),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_866),
.B(n_975),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_SL g1088 ( 
.A1(n_931),
.A2(n_908),
.B(n_928),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_926),
.A2(n_918),
.B(n_897),
.C(n_898),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_866),
.Y(n_1090)
);

AO21x1_ASAP7_75t_L g1091 ( 
.A1(n_913),
.A2(n_900),
.B(n_975),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_935),
.A2(n_543),
.B(n_538),
.Y(n_1092)
);

BUFx4f_ASAP7_75t_L g1093 ( 
.A(n_935),
.Y(n_1093)
);

AOI21x1_ASAP7_75t_L g1094 ( 
.A1(n_874),
.A2(n_877),
.B(n_883),
.Y(n_1094)
);

AO21x1_ASAP7_75t_L g1095 ( 
.A1(n_1012),
.A2(n_676),
.B(n_842),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_990),
.B(n_1001),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_950),
.A2(n_543),
.B(n_538),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_950),
.A2(n_543),
.B(n_538),
.Y(n_1098)
);

INVx1_ASAP7_75t_SL g1099 ( 
.A(n_995),
.Y(n_1099)
);

OR2x2_ASAP7_75t_L g1100 ( 
.A(n_992),
.B(n_526),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_856),
.B(n_688),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_990),
.B(n_1001),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_992),
.B(n_526),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_882),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_950),
.A2(n_543),
.B(n_538),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_990),
.B(n_1001),
.Y(n_1106)
);

INVx2_ASAP7_75t_SL g1107 ( 
.A(n_1010),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_838),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_990),
.B(n_1001),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_950),
.A2(n_543),
.B(n_538),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_950),
.A2(n_543),
.B(n_538),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_935),
.Y(n_1112)
);

AO31x2_ASAP7_75t_L g1113 ( 
.A1(n_1012),
.A2(n_986),
.A3(n_1011),
.B(n_1007),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_992),
.B(n_676),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_838),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_950),
.A2(n_543),
.B(n_538),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_990),
.B(n_1001),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_915),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_950),
.A2(n_543),
.B(n_538),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_990),
.B(n_1001),
.Y(n_1120)
);

OAI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1012),
.A2(n_986),
.B(n_676),
.Y(n_1121)
);

O2A1O1Ixp5_ASAP7_75t_L g1122 ( 
.A1(n_849),
.A2(n_676),
.B(n_889),
.C(n_986),
.Y(n_1122)
);

INVx4_ASAP7_75t_L g1123 ( 
.A(n_838),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_952),
.A2(n_884),
.B(n_981),
.Y(n_1124)
);

OAI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1012),
.A2(n_986),
.B(n_676),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_952),
.A2(n_884),
.B(n_981),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_842),
.A2(n_676),
.B(n_849),
.C(n_1004),
.Y(n_1127)
);

AO31x2_ASAP7_75t_L g1128 ( 
.A1(n_1012),
.A2(n_986),
.A3(n_1011),
.B(n_1007),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_SL g1129 ( 
.A1(n_842),
.A2(n_676),
.B(n_715),
.Y(n_1129)
);

OAI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1012),
.A2(n_986),
.B(n_676),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_885),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_992),
.B(n_526),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_990),
.B(n_1001),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_935),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1012),
.A2(n_986),
.B(n_676),
.Y(n_1135)
);

OAI22x1_ASAP7_75t_L g1136 ( 
.A1(n_992),
.A2(n_842),
.B1(n_916),
.B2(n_676),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_990),
.B(n_1001),
.Y(n_1137)
);

HB1xp67_ASAP7_75t_L g1138 ( 
.A(n_1010),
.Y(n_1138)
);

OR2x2_ASAP7_75t_L g1139 ( 
.A(n_992),
.B(n_526),
.Y(n_1139)
);

INVx6_ASAP7_75t_L g1140 ( 
.A(n_915),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_952),
.A2(n_884),
.B(n_981),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_952),
.A2(n_884),
.B(n_981),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_885),
.Y(n_1143)
);

AO31x2_ASAP7_75t_L g1144 ( 
.A1(n_1012),
.A2(n_986),
.A3(n_1011),
.B(n_1007),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_990),
.B(n_1001),
.Y(n_1145)
);

AOI21x1_ASAP7_75t_L g1146 ( 
.A1(n_874),
.A2(n_877),
.B(n_883),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_952),
.A2(n_884),
.B(n_981),
.Y(n_1147)
);

INVx5_ASAP7_75t_L g1148 ( 
.A(n_935),
.Y(n_1148)
);

AOI21x1_ASAP7_75t_SL g1149 ( 
.A1(n_889),
.A2(n_947),
.B(n_930),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1012),
.A2(n_986),
.B(n_676),
.Y(n_1150)
);

OR2x2_ASAP7_75t_L g1151 ( 
.A(n_992),
.B(n_526),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_952),
.A2(n_884),
.B(n_981),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_950),
.A2(n_543),
.B(n_538),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1012),
.A2(n_986),
.B(n_676),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_990),
.B(n_1001),
.Y(n_1155)
);

AOI21xp33_ASAP7_75t_L g1156 ( 
.A1(n_849),
.A2(n_676),
.B(n_842),
.Y(n_1156)
);

AOI21xp33_ASAP7_75t_L g1157 ( 
.A1(n_849),
.A2(n_676),
.B(n_842),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_952),
.A2(n_884),
.B(n_981),
.Y(n_1158)
);

AO31x2_ASAP7_75t_L g1159 ( 
.A1(n_1012),
.A2(n_986),
.A3(n_1011),
.B(n_1007),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_990),
.B(n_1001),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1096),
.B(n_1102),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1099),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1019),
.Y(n_1163)
);

NOR2xp67_ASAP7_75t_L g1164 ( 
.A(n_1104),
.B(n_1050),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1131),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1114),
.A2(n_1129),
.B(n_1127),
.C(n_1016),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1018),
.B(n_1103),
.Y(n_1167)
);

A2O1A1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_1156),
.A2(n_1157),
.B(n_1121),
.C(n_1154),
.Y(n_1168)
);

CKINVDCx8_ASAP7_75t_R g1169 ( 
.A(n_1065),
.Y(n_1169)
);

CKINVDCx20_ASAP7_75t_R g1170 ( 
.A(n_1040),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1101),
.B(n_1045),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_1112),
.Y(n_1172)
);

CKINVDCx20_ASAP7_75t_R g1173 ( 
.A(n_1118),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1020),
.A2(n_1044),
.B(n_1042),
.Y(n_1174)
);

BUFx12f_ASAP7_75t_L g1175 ( 
.A(n_1140),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1034),
.A2(n_1036),
.B(n_1121),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1143),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1052),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1096),
.B(n_1102),
.Y(n_1179)
);

BUFx8_ASAP7_75t_SL g1180 ( 
.A(n_1022),
.Y(n_1180)
);

NAND3xp33_ASAP7_75t_L g1181 ( 
.A(n_1156),
.B(n_1157),
.C(n_1122),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_1100),
.B(n_1139),
.Y(n_1182)
);

HB1xp67_ASAP7_75t_L g1183 ( 
.A(n_1099),
.Y(n_1183)
);

INVx4_ASAP7_75t_L g1184 ( 
.A(n_1148),
.Y(n_1184)
);

INVx5_ASAP7_75t_L g1185 ( 
.A(n_1112),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1125),
.A2(n_1135),
.B(n_1130),
.C(n_1154),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_1138),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1125),
.A2(n_1135),
.B(n_1130),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1106),
.B(n_1109),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1150),
.A2(n_1053),
.B(n_1049),
.Y(n_1190)
);

NAND2x1p5_ASAP7_75t_L g1191 ( 
.A(n_1148),
.B(n_1093),
.Y(n_1191)
);

INVx5_ASAP7_75t_L g1192 ( 
.A(n_1112),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_1140),
.Y(n_1193)
);

OAI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1150),
.A2(n_1066),
.B(n_1051),
.Y(n_1194)
);

INVx1_ASAP7_75t_SL g1195 ( 
.A(n_1151),
.Y(n_1195)
);

AND2x2_ASAP7_75t_SL g1196 ( 
.A(n_1132),
.B(n_1033),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1033),
.B(n_1101),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_1045),
.B(n_1085),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1106),
.B(n_1109),
.Y(n_1199)
);

OAI22x1_ASAP7_75t_L g1200 ( 
.A1(n_1030),
.A2(n_1037),
.B1(n_1060),
.B2(n_1155),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1117),
.B(n_1120),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1021),
.B(n_1046),
.Y(n_1202)
);

NOR2xp67_ASAP7_75t_SL g1203 ( 
.A(n_1148),
.B(n_1107),
.Y(n_1203)
);

OAI21xp33_ASAP7_75t_L g1204 ( 
.A1(n_1117),
.A2(n_1160),
.B(n_1155),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1120),
.B(n_1133),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_1022),
.Y(n_1206)
);

NAND2x1p5_ASAP7_75t_L g1207 ( 
.A(n_1148),
.B(n_1093),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1133),
.A2(n_1160),
.B1(n_1145),
.B2(n_1137),
.Y(n_1208)
);

NAND3xp33_ASAP7_75t_SL g1209 ( 
.A(n_1068),
.B(n_1095),
.C(n_1069),
.Y(n_1209)
);

CKINVDCx20_ASAP7_75t_R g1210 ( 
.A(n_1081),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_1134),
.Y(n_1211)
);

INVxp67_ASAP7_75t_L g1212 ( 
.A(n_1054),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1022),
.B(n_1027),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1014),
.A2(n_1035),
.B(n_1051),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1136),
.A2(n_1017),
.B1(n_1023),
.B2(n_1137),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1035),
.A2(n_1057),
.B(n_1145),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1032),
.B(n_1031),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_1090),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1055),
.B(n_1061),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1061),
.B(n_1017),
.Y(n_1220)
);

A2O1A1Ixp33_ASAP7_75t_SL g1221 ( 
.A1(n_1064),
.A2(n_1070),
.B(n_1086),
.C(n_1080),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1028),
.B(n_1043),
.Y(n_1222)
);

NOR2x1p5_ASAP7_75t_L g1223 ( 
.A(n_1076),
.B(n_1078),
.Y(n_1223)
);

AOI21xp33_ASAP7_75t_L g1224 ( 
.A1(n_1039),
.A2(n_1088),
.B(n_1048),
.Y(n_1224)
);

NAND2xp33_ASAP7_75t_SL g1225 ( 
.A(n_1134),
.B(n_1123),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1070),
.A2(n_1077),
.B1(n_1064),
.B2(n_1089),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1087),
.B(n_1074),
.Y(n_1227)
);

AOI222xp33_ASAP7_75t_L g1228 ( 
.A1(n_1073),
.A2(n_1071),
.B1(n_1086),
.B2(n_1075),
.C1(n_1041),
.C2(n_1082),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1056),
.B(n_1108),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1113),
.B(n_1159),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1071),
.A2(n_1059),
.B1(n_1108),
.B2(n_1115),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1097),
.A2(n_1098),
.B(n_1153),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1105),
.A2(n_1119),
.B(n_1116),
.Y(n_1233)
);

INVxp67_ASAP7_75t_SL g1234 ( 
.A(n_1084),
.Y(n_1234)
);

AND2x2_ASAP7_75t_SL g1235 ( 
.A(n_1091),
.B(n_1149),
.Y(n_1235)
);

NOR2x1p5_ASAP7_75t_SL g1236 ( 
.A(n_1024),
.B(n_1146),
.Y(n_1236)
);

INVx5_ASAP7_75t_L g1237 ( 
.A(n_1083),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1048),
.A2(n_1063),
.B1(n_1072),
.B2(n_1062),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1113),
.Y(n_1239)
);

NAND2x1p5_ASAP7_75t_L g1240 ( 
.A(n_1079),
.B(n_1026),
.Y(n_1240)
);

O2A1O1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1110),
.A2(n_1111),
.B(n_1092),
.C(n_1083),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1094),
.A2(n_1159),
.B1(n_1144),
.B2(n_1128),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1029),
.A2(n_1038),
.B(n_1047),
.Y(n_1243)
);

INVx5_ASAP7_75t_L g1244 ( 
.A(n_1083),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_1128),
.Y(n_1245)
);

A2O1A1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1015),
.A2(n_1141),
.B(n_1158),
.C(n_1142),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1124),
.A2(n_1126),
.B(n_1152),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1128),
.A2(n_1144),
.B1(n_1159),
.B2(n_1147),
.Y(n_1248)
);

INVxp67_ASAP7_75t_L g1249 ( 
.A(n_1025),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1144),
.Y(n_1250)
);

OR2x2_ASAP7_75t_L g1251 ( 
.A(n_1067),
.B(n_1058),
.Y(n_1251)
);

BUFx2_ASAP7_75t_L g1252 ( 
.A(n_1138),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1096),
.B(n_990),
.Y(n_1253)
);

AO21x1_ASAP7_75t_L g1254 ( 
.A1(n_1129),
.A2(n_1157),
.B(n_1156),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1096),
.B(n_990),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1018),
.B(n_1103),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1096),
.B(n_990),
.Y(n_1257)
);

AND2x4_ASAP7_75t_SL g1258 ( 
.A(n_1138),
.B(n_792),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1096),
.B(n_990),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1018),
.B(n_1103),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1018),
.B(n_1103),
.Y(n_1261)
);

INVx5_ASAP7_75t_L g1262 ( 
.A(n_1112),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1020),
.A2(n_1044),
.B(n_1042),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1018),
.B(n_1103),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1101),
.B(n_1045),
.Y(n_1265)
);

OR2x2_ASAP7_75t_SL g1266 ( 
.A(n_1100),
.B(n_916),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1114),
.B(n_992),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1114),
.B(n_990),
.Y(n_1268)
);

A2O1A1Ixp33_ASAP7_75t_SL g1269 ( 
.A1(n_1121),
.A2(n_676),
.B(n_849),
.C(n_679),
.Y(n_1269)
);

A2O1A1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1114),
.A2(n_676),
.B(n_842),
.C(n_1004),
.Y(n_1270)
);

OR2x6_ASAP7_75t_L g1271 ( 
.A(n_1022),
.B(n_926),
.Y(n_1271)
);

NAND2x1p5_ASAP7_75t_L g1272 ( 
.A(n_1148),
.B(n_1093),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1018),
.B(n_1103),
.Y(n_1273)
);

BUFx12f_ASAP7_75t_L g1274 ( 
.A(n_1104),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1018),
.B(n_1103),
.Y(n_1275)
);

INVx3_ASAP7_75t_SL g1276 ( 
.A(n_1104),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1114),
.B(n_990),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_SL g1278 ( 
.A(n_1127),
.B(n_1012),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1114),
.B(n_992),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_SL g1280 ( 
.A1(n_1114),
.A2(n_676),
.B1(n_992),
.B2(n_360),
.Y(n_1280)
);

OR2x2_ASAP7_75t_L g1281 ( 
.A(n_1100),
.B(n_526),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_1101),
.B(n_1045),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1018),
.B(n_1103),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1114),
.B(n_990),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1114),
.B(n_990),
.Y(n_1285)
);

INVx2_ASAP7_75t_SL g1286 ( 
.A(n_1099),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1101),
.B(n_1045),
.Y(n_1287)
);

AND2x6_ASAP7_75t_L g1288 ( 
.A(n_1043),
.B(n_985),
.Y(n_1288)
);

INVx1_ASAP7_75t_SL g1289 ( 
.A(n_1099),
.Y(n_1289)
);

AO22x2_ASAP7_75t_L g1290 ( 
.A1(n_1129),
.A2(n_1012),
.B1(n_1135),
.B2(n_1150),
.Y(n_1290)
);

NAND2x1p5_ASAP7_75t_L g1291 ( 
.A(n_1148),
.B(n_1093),
.Y(n_1291)
);

INVxp67_ASAP7_75t_L g1292 ( 
.A(n_1138),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_1101),
.B(n_1045),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1099),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1165),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1177),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1270),
.A2(n_1279),
.B(n_1267),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1280),
.B(n_1268),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1278),
.A2(n_1209),
.B1(n_1290),
.B2(n_1254),
.Y(n_1299)
);

AO21x2_ASAP7_75t_L g1300 ( 
.A1(n_1243),
.A2(n_1247),
.B(n_1174),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1239),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_L g1302 ( 
.A(n_1162),
.Y(n_1302)
);

OR2x2_ASAP7_75t_L g1303 ( 
.A(n_1168),
.B(n_1230),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1166),
.B(n_1215),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_L g1305 ( 
.A(n_1185),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1278),
.A2(n_1290),
.B1(n_1188),
.B2(n_1194),
.Y(n_1306)
);

OAI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1269),
.A2(n_1186),
.B(n_1181),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1194),
.A2(n_1196),
.B1(n_1226),
.B2(n_1202),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1243),
.A2(n_1233),
.B(n_1232),
.Y(n_1309)
);

BUFx2_ASAP7_75t_R g1310 ( 
.A(n_1180),
.Y(n_1310)
);

CKINVDCx6p67_ASAP7_75t_R g1311 ( 
.A(n_1276),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1252),
.Y(n_1312)
);

BUFx3_ASAP7_75t_L g1313 ( 
.A(n_1171),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1277),
.B(n_1284),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1250),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1230),
.Y(n_1316)
);

AOI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1164),
.A2(n_1285),
.B1(n_1199),
.B2(n_1201),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1245),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1198),
.B(n_1271),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1220),
.B(n_1161),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1191),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_SL g1322 ( 
.A1(n_1195),
.A2(n_1182),
.B1(n_1212),
.B2(n_1170),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1178),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1226),
.A2(n_1261),
.B1(n_1167),
.B2(n_1260),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1171),
.Y(n_1325)
);

INVxp67_ASAP7_75t_SL g1326 ( 
.A(n_1183),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1161),
.B(n_1205),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1256),
.A2(n_1264),
.B1(n_1283),
.B2(n_1275),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1205),
.B(n_1179),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1217),
.Y(n_1330)
);

INVx6_ASAP7_75t_L g1331 ( 
.A(n_1185),
.Y(n_1331)
);

BUFx2_ASAP7_75t_R g1332 ( 
.A(n_1169),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1197),
.Y(n_1333)
);

INVx2_ASAP7_75t_SL g1334 ( 
.A(n_1185),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_SL g1335 ( 
.A1(n_1181),
.A2(n_1208),
.B1(n_1195),
.B2(n_1273),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1227),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1198),
.B(n_1271),
.Y(n_1337)
);

BUFx2_ASAP7_75t_L g1338 ( 
.A(n_1294),
.Y(n_1338)
);

NAND2x1p5_ASAP7_75t_L g1339 ( 
.A(n_1237),
.B(n_1244),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1218),
.Y(n_1340)
);

AOI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1214),
.A2(n_1176),
.B(n_1216),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1189),
.B(n_1208),
.Y(n_1342)
);

CKINVDCx11_ASAP7_75t_R g1343 ( 
.A(n_1175),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_SL g1344 ( 
.A1(n_1190),
.A2(n_1255),
.B1(n_1253),
.B2(n_1257),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1237),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1229),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1219),
.Y(n_1347)
);

INVx4_ASAP7_75t_L g1348 ( 
.A(n_1192),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1274),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1200),
.A2(n_1204),
.B1(n_1253),
.B2(n_1255),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_L g1351 ( 
.A(n_1192),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1289),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1204),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1281),
.B(n_1292),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1289),
.B(n_1258),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1191),
.Y(n_1356)
);

OAI21xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1257),
.A2(n_1259),
.B(n_1228),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_SL g1358 ( 
.A1(n_1259),
.A2(n_1210),
.B1(n_1206),
.B2(n_1288),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1244),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1266),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1244),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1286),
.A2(n_1187),
.B1(n_1213),
.B2(n_1271),
.Y(n_1362)
);

NAND2x1_ASAP7_75t_L g1363 ( 
.A(n_1288),
.B(n_1238),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1288),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1203),
.Y(n_1365)
);

NAND2x1p5_ASAP7_75t_L g1366 ( 
.A(n_1235),
.B(n_1251),
.Y(n_1366)
);

AOI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1213),
.A2(n_1193),
.B1(n_1287),
.B2(n_1293),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1222),
.B(n_1228),
.Y(n_1368)
);

INVxp67_ASAP7_75t_L g1369 ( 
.A(n_1265),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1222),
.B(n_1242),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1231),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1172),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1249),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1293),
.B(n_1282),
.Y(n_1374)
);

NAND2x1p5_ASAP7_75t_L g1375 ( 
.A(n_1263),
.B(n_1262),
.Y(n_1375)
);

BUFx3_ASAP7_75t_L g1376 ( 
.A(n_1265),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1240),
.A2(n_1241),
.B(n_1248),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1172),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1224),
.B(n_1248),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1282),
.A2(n_1287),
.B1(n_1207),
.B2(n_1272),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1211),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1224),
.B(n_1288),
.Y(n_1382)
);

OR2x6_ASAP7_75t_L g1383 ( 
.A(n_1236),
.B(n_1246),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_SL g1384 ( 
.A1(n_1173),
.A2(n_1207),
.B1(n_1272),
.B2(n_1291),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1234),
.Y(n_1385)
);

OA21x2_ASAP7_75t_L g1386 ( 
.A1(n_1221),
.A2(n_1225),
.B(n_1291),
.Y(n_1386)
);

BUFx2_ASAP7_75t_L g1387 ( 
.A(n_1262),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1262),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1223),
.Y(n_1389)
);

CKINVDCx11_ASAP7_75t_R g1390 ( 
.A(n_1169),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1267),
.A2(n_676),
.B1(n_1279),
.B2(n_1114),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_1274),
.Y(n_1392)
);

INVx3_ASAP7_75t_L g1393 ( 
.A(n_1184),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1280),
.A2(n_1114),
.B1(n_676),
.B2(n_1267),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1163),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1267),
.A2(n_676),
.B1(n_1279),
.B2(n_1114),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1303),
.B(n_1316),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1320),
.B(n_1307),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1377),
.A2(n_1309),
.B(n_1341),
.Y(n_1399)
);

AOI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1341),
.A2(n_1363),
.B(n_1383),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1301),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1315),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1303),
.B(n_1316),
.Y(n_1403)
);

CKINVDCx20_ASAP7_75t_R g1404 ( 
.A(n_1390),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1320),
.B(n_1306),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_1363),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_1338),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_1338),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1383),
.Y(n_1409)
);

INVxp67_ASAP7_75t_L g1410 ( 
.A(n_1352),
.Y(n_1410)
);

BUFx6f_ASAP7_75t_L g1411 ( 
.A(n_1383),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1370),
.B(n_1379),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1347),
.B(n_1342),
.Y(n_1413)
);

BUFx6f_ASAP7_75t_L g1414 ( 
.A(n_1383),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1394),
.A2(n_1298),
.B1(n_1297),
.B2(n_1304),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1375),
.A2(n_1339),
.B(n_1371),
.Y(n_1416)
);

OA21x2_ASAP7_75t_L g1417 ( 
.A1(n_1379),
.A2(n_1299),
.B(n_1370),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1373),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1385),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1318),
.Y(n_1420)
);

AO21x2_ASAP7_75t_L g1421 ( 
.A1(n_1300),
.A2(n_1382),
.B(n_1368),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1353),
.Y(n_1422)
);

OR2x6_ASAP7_75t_L g1423 ( 
.A(n_1364),
.B(n_1366),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1342),
.B(n_1327),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1327),
.B(n_1344),
.Y(n_1425)
);

INVxp67_ASAP7_75t_L g1426 ( 
.A(n_1326),
.Y(n_1426)
);

INVx1_ASAP7_75t_SL g1427 ( 
.A(n_1302),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1300),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1329),
.B(n_1304),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1329),
.B(n_1368),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_SL g1431 ( 
.A(n_1332),
.Y(n_1431)
);

OA21x2_ASAP7_75t_L g1432 ( 
.A1(n_1382),
.A2(n_1308),
.B(n_1350),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1323),
.B(n_1360),
.Y(n_1433)
);

AO31x2_ASAP7_75t_L g1434 ( 
.A1(n_1364),
.A2(n_1345),
.A3(n_1361),
.B(n_1359),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1357),
.B(n_1336),
.Y(n_1435)
);

INVx2_ASAP7_75t_SL g1436 ( 
.A(n_1331),
.Y(n_1436)
);

AOI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1386),
.A2(n_1362),
.B(n_1365),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1333),
.Y(n_1438)
);

CKINVDCx6p67_ASAP7_75t_R g1439 ( 
.A(n_1343),
.Y(n_1439)
);

AO21x2_ASAP7_75t_L g1440 ( 
.A1(n_1317),
.A2(n_1295),
.B(n_1296),
.Y(n_1440)
);

INVxp33_ASAP7_75t_L g1441 ( 
.A(n_1355),
.Y(n_1441)
);

AO21x1_ASAP7_75t_SL g1442 ( 
.A1(n_1324),
.A2(n_1330),
.B(n_1346),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1314),
.B(n_1369),
.Y(n_1443)
);

OAI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1391),
.A2(n_1396),
.B(n_1335),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1328),
.B(n_1395),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_SL g1446 ( 
.A1(n_1305),
.A2(n_1351),
.B(n_1348),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1358),
.B(n_1337),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1312),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1319),
.B(n_1337),
.Y(n_1449)
);

INVx2_ASAP7_75t_SL g1450 ( 
.A(n_1331),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1401),
.Y(n_1451)
);

INVx4_ASAP7_75t_L g1452 ( 
.A(n_1440),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1419),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1412),
.B(n_1322),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1412),
.B(n_1340),
.Y(n_1455)
);

INVxp67_ASAP7_75t_L g1456 ( 
.A(n_1440),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1424),
.B(n_1354),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1412),
.B(n_1337),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1421),
.B(n_1312),
.Y(n_1459)
);

BUFx2_ASAP7_75t_L g1460 ( 
.A(n_1434),
.Y(n_1460)
);

INVx5_ASAP7_75t_L g1461 ( 
.A(n_1409),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1415),
.A2(n_1376),
.B1(n_1325),
.B2(n_1313),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1421),
.B(n_1397),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1409),
.B(n_1356),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1424),
.B(n_1384),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1435),
.B(n_1367),
.Y(n_1466)
);

OAI211xp5_ASAP7_75t_L g1467 ( 
.A1(n_1444),
.A2(n_1390),
.B(n_1343),
.C(n_1389),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1444),
.A2(n_1376),
.B1(n_1325),
.B2(n_1313),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1435),
.B(n_1356),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1434),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1421),
.B(n_1372),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1421),
.B(n_1417),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1422),
.B(n_1321),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1398),
.B(n_1381),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1398),
.A2(n_1389),
.B1(n_1374),
.B2(n_1311),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1402),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1417),
.B(n_1378),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_1409),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1399),
.A2(n_1393),
.B(n_1380),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1417),
.B(n_1374),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1422),
.B(n_1387),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1417),
.B(n_1374),
.Y(n_1482)
);

INVx1_ASAP7_75t_SL g1483 ( 
.A(n_1427),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1417),
.B(n_1388),
.Y(n_1484)
);

INVx4_ASAP7_75t_L g1485 ( 
.A(n_1440),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1434),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1403),
.B(n_1311),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1430),
.B(n_1305),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_1404),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1430),
.B(n_1305),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1483),
.B(n_1427),
.Y(n_1491)
);

AOI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1467),
.A2(n_1447),
.B1(n_1432),
.B2(n_1406),
.Y(n_1492)
);

NAND3xp33_ASAP7_75t_L g1493 ( 
.A(n_1467),
.B(n_1425),
.C(n_1445),
.Y(n_1493)
);

OA21x2_ASAP7_75t_L g1494 ( 
.A1(n_1456),
.A2(n_1399),
.B(n_1428),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1466),
.A2(n_1406),
.B1(n_1447),
.B2(n_1432),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1483),
.B(n_1410),
.Y(n_1496)
);

NAND3xp33_ASAP7_75t_L g1497 ( 
.A(n_1466),
.B(n_1425),
.C(n_1445),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_SL g1498 ( 
.A1(n_1472),
.A2(n_1406),
.B1(n_1432),
.B2(n_1405),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1480),
.B(n_1423),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1469),
.B(n_1474),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1469),
.B(n_1474),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1455),
.B(n_1410),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_SL g1503 ( 
.A(n_1487),
.B(n_1406),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1480),
.B(n_1423),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_R g1505 ( 
.A(n_1489),
.B(n_1431),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1455),
.B(n_1426),
.Y(n_1506)
);

NAND3xp33_ASAP7_75t_L g1507 ( 
.A(n_1468),
.B(n_1438),
.C(n_1443),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1455),
.B(n_1426),
.Y(n_1508)
);

OAI21xp5_ASAP7_75t_SL g1509 ( 
.A1(n_1475),
.A2(n_1472),
.B(n_1462),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1482),
.B(n_1423),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1482),
.B(n_1423),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1487),
.A2(n_1431),
.B1(n_1439),
.B2(n_1441),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_SL g1513 ( 
.A(n_1461),
.B(n_1406),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1484),
.B(n_1423),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1451),
.Y(n_1515)
);

NAND3xp33_ASAP7_75t_L g1516 ( 
.A(n_1459),
.B(n_1438),
.C(n_1406),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1484),
.B(n_1423),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1477),
.B(n_1413),
.Y(n_1518)
);

OAI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1479),
.A2(n_1437),
.B(n_1416),
.Y(n_1519)
);

NAND4xp25_ASAP7_75t_L g1520 ( 
.A(n_1459),
.B(n_1457),
.C(n_1471),
.D(n_1481),
.Y(n_1520)
);

OAI21xp5_ASAP7_75t_SL g1521 ( 
.A1(n_1472),
.A2(n_1405),
.B(n_1406),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1458),
.B(n_1407),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1476),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1477),
.B(n_1413),
.Y(n_1524)
);

OAI21xp5_ASAP7_75t_SL g1525 ( 
.A1(n_1454),
.A2(n_1449),
.B(n_1429),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1477),
.B(n_1432),
.Y(n_1526)
);

OAI221xp5_ASAP7_75t_L g1527 ( 
.A1(n_1457),
.A2(n_1448),
.B1(n_1432),
.B2(n_1450),
.C(n_1436),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1458),
.B(n_1407),
.Y(n_1528)
);

OAI21xp5_ASAP7_75t_SL g1529 ( 
.A1(n_1454),
.A2(n_1449),
.B(n_1429),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1471),
.B(n_1434),
.Y(n_1530)
);

OAI21xp33_ASAP7_75t_L g1531 ( 
.A1(n_1465),
.A2(n_1433),
.B(n_1437),
.Y(n_1531)
);

NAND3xp33_ASAP7_75t_L g1532 ( 
.A(n_1481),
.B(n_1433),
.C(n_1420),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_L g1533 ( 
.A(n_1454),
.B(n_1439),
.Y(n_1533)
);

NAND3xp33_ASAP7_75t_SL g1534 ( 
.A(n_1465),
.B(n_1448),
.C(n_1392),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1458),
.B(n_1407),
.Y(n_1535)
);

NOR3xp33_ASAP7_75t_L g1536 ( 
.A(n_1452),
.B(n_1450),
.C(n_1436),
.Y(n_1536)
);

OAI21xp5_ASAP7_75t_SL g1537 ( 
.A1(n_1464),
.A2(n_1449),
.B(n_1411),
.Y(n_1537)
);

OAI21xp5_ASAP7_75t_SL g1538 ( 
.A1(n_1464),
.A2(n_1411),
.B(n_1414),
.Y(n_1538)
);

OA21x2_ASAP7_75t_L g1539 ( 
.A1(n_1456),
.A2(n_1428),
.B(n_1416),
.Y(n_1539)
);

AOI21xp33_ASAP7_75t_L g1540 ( 
.A1(n_1471),
.A2(n_1440),
.B(n_1450),
.Y(n_1540)
);

NAND3xp33_ASAP7_75t_L g1541 ( 
.A(n_1452),
.B(n_1420),
.C(n_1418),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1451),
.B(n_1434),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1451),
.B(n_1434),
.Y(n_1543)
);

NOR3xp33_ASAP7_75t_L g1544 ( 
.A(n_1452),
.B(n_1436),
.C(n_1400),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1488),
.B(n_1490),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1488),
.B(n_1408),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1490),
.B(n_1408),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1523),
.B(n_1500),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1542),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1513),
.B(n_1461),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1526),
.B(n_1460),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1526),
.B(n_1460),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1530),
.B(n_1470),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1530),
.B(n_1470),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1515),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1501),
.B(n_1463),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1518),
.B(n_1463),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1543),
.Y(n_1558)
);

INVxp67_ASAP7_75t_SL g1559 ( 
.A(n_1541),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1520),
.B(n_1524),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1524),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1514),
.Y(n_1562)
);

INVxp67_ASAP7_75t_L g1563 ( 
.A(n_1527),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1532),
.B(n_1486),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1521),
.B(n_1476),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1517),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1539),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1531),
.B(n_1453),
.Y(n_1568)
);

INVx4_ASAP7_75t_L g1569 ( 
.A(n_1494),
.Y(n_1569)
);

INVx3_ASAP7_75t_L g1570 ( 
.A(n_1494),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1506),
.B(n_1453),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1499),
.B(n_1452),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1508),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1499),
.Y(n_1574)
);

NAND2x1_ASAP7_75t_L g1575 ( 
.A(n_1516),
.B(n_1478),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1504),
.B(n_1485),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1504),
.Y(n_1577)
);

INVx4_ASAP7_75t_L g1578 ( 
.A(n_1510),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1491),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1510),
.B(n_1485),
.Y(n_1580)
);

AND2x4_ASAP7_75t_SL g1581 ( 
.A(n_1511),
.B(n_1411),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1502),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1513),
.B(n_1461),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1511),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1545),
.Y(n_1585)
);

OAI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1563),
.A2(n_1497),
.B(n_1493),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1561),
.Y(n_1587)
);

OAI21xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1559),
.A2(n_1503),
.B(n_1492),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1560),
.B(n_1496),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1560),
.B(n_1546),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1560),
.B(n_1547),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1578),
.B(n_1498),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1555),
.Y(n_1593)
);

INVx1_ASAP7_75t_SL g1594 ( 
.A(n_1579),
.Y(n_1594)
);

INVx2_ASAP7_75t_SL g1595 ( 
.A(n_1581),
.Y(n_1595)
);

NOR3xp33_ASAP7_75t_L g1596 ( 
.A(n_1563),
.B(n_1534),
.C(n_1512),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1578),
.B(n_1538),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1561),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1557),
.B(n_1522),
.Y(n_1599)
);

OAI21xp33_ASAP7_75t_L g1600 ( 
.A1(n_1559),
.A2(n_1509),
.B(n_1495),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1578),
.B(n_1537),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1557),
.B(n_1528),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1561),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1578),
.B(n_1461),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1578),
.B(n_1574),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1564),
.B(n_1535),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1564),
.B(n_1503),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1574),
.B(n_1461),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1579),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1574),
.B(n_1461),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1574),
.B(n_1461),
.Y(n_1611)
);

NOR2xp67_ASAP7_75t_L g1612 ( 
.A(n_1550),
.B(n_1485),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1585),
.B(n_1573),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1585),
.B(n_1525),
.Y(n_1614)
);

INVx4_ASAP7_75t_L g1615 ( 
.A(n_1550),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1584),
.B(n_1478),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1555),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1555),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1555),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1584),
.B(n_1553),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1568),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1584),
.B(n_1478),
.Y(n_1622)
);

OR2x6_ASAP7_75t_L g1623 ( 
.A(n_1575),
.B(n_1550),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1589),
.B(n_1556),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1601),
.B(n_1577),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1601),
.B(n_1577),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1609),
.Y(n_1627)
);

OAI31xp33_ASAP7_75t_L g1628 ( 
.A1(n_1600),
.A2(n_1565),
.A3(n_1507),
.B(n_1583),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1586),
.B(n_1585),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1589),
.B(n_1556),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1590),
.B(n_1568),
.Y(n_1631)
);

O2A1O1Ixp33_ASAP7_75t_L g1632 ( 
.A1(n_1588),
.A2(n_1575),
.B(n_1564),
.C(n_1565),
.Y(n_1632)
);

NAND4xp25_ASAP7_75t_L g1633 ( 
.A(n_1600),
.B(n_1533),
.C(n_1565),
.D(n_1544),
.Y(n_1633)
);

NOR2x2_ASAP7_75t_L g1634 ( 
.A(n_1623),
.B(n_1584),
.Y(n_1634)
);

INVx2_ASAP7_75t_SL g1635 ( 
.A(n_1595),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1590),
.B(n_1582),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1594),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1597),
.B(n_1577),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1597),
.B(n_1550),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1587),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1587),
.Y(n_1641)
);

OAI33xp33_ASAP7_75t_L g1642 ( 
.A1(n_1613),
.A2(n_1573),
.A3(n_1571),
.B1(n_1582),
.B2(n_1548),
.B3(n_1473),
.Y(n_1642)
);

BUFx2_ASAP7_75t_SL g1643 ( 
.A(n_1595),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1598),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1592),
.B(n_1562),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1615),
.B(n_1550),
.Y(n_1646)
);

AOI222xp33_ASAP7_75t_L g1647 ( 
.A1(n_1588),
.A2(n_1573),
.B1(n_1529),
.B2(n_1553),
.C1(n_1554),
.C2(n_1548),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1592),
.B(n_1562),
.Y(n_1648)
);

NAND2xp33_ASAP7_75t_L g1649 ( 
.A(n_1596),
.B(n_1505),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1614),
.B(n_1562),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1621),
.B(n_1566),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1591),
.B(n_1566),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1591),
.B(n_1606),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1599),
.B(n_1439),
.Y(n_1654)
);

AOI21xp33_ASAP7_75t_L g1655 ( 
.A1(n_1607),
.A2(n_1575),
.B(n_1623),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1606),
.B(n_1566),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1604),
.B(n_1572),
.Y(n_1657)
);

OAI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1623),
.A2(n_1581),
.B1(n_1583),
.B2(n_1550),
.Y(n_1658)
);

NAND5xp2_ASAP7_75t_L g1659 ( 
.A(n_1604),
.B(n_1536),
.C(n_1519),
.D(n_1540),
.E(n_1572),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1605),
.B(n_1572),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1598),
.Y(n_1661)
);

INVx2_ASAP7_75t_SL g1662 ( 
.A(n_1615),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1603),
.Y(n_1663)
);

OAI21xp33_ASAP7_75t_L g1664 ( 
.A1(n_1607),
.A2(n_1571),
.B(n_1576),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1599),
.A2(n_1442),
.B1(n_1485),
.B2(n_1414),
.Y(n_1665)
);

AND2x4_ASAP7_75t_L g1666 ( 
.A(n_1615),
.B(n_1583),
.Y(n_1666)
);

NAND3x1_ASAP7_75t_SL g1667 ( 
.A(n_1628),
.B(n_1310),
.C(n_1505),
.Y(n_1667)
);

INVx1_ASAP7_75t_SL g1668 ( 
.A(n_1637),
.Y(n_1668)
);

INVx1_ASAP7_75t_SL g1669 ( 
.A(n_1637),
.Y(n_1669)
);

NOR2x1_ASAP7_75t_L g1670 ( 
.A(n_1649),
.B(n_1623),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1643),
.B(n_1615),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1654),
.B(n_1349),
.Y(n_1672)
);

INVx1_ASAP7_75t_SL g1673 ( 
.A(n_1634),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1640),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1645),
.B(n_1648),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1641),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1629),
.B(n_1602),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1644),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1638),
.B(n_1623),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1654),
.B(n_1602),
.Y(n_1680)
);

OAI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1633),
.A2(n_1650),
.B1(n_1658),
.B2(n_1631),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1649),
.B(n_1659),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1661),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1639),
.B(n_1605),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1639),
.B(n_1620),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1627),
.B(n_1620),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1647),
.B(n_1583),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1639),
.A2(n_1583),
.B1(n_1411),
.B2(n_1414),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1625),
.B(n_1616),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1653),
.B(n_1603),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1626),
.B(n_1608),
.Y(n_1691)
);

INVx1_ASAP7_75t_SL g1692 ( 
.A(n_1634),
.Y(n_1692)
);

AO21x2_ASAP7_75t_L g1693 ( 
.A1(n_1632),
.A2(n_1655),
.B(n_1612),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1665),
.A2(n_1583),
.B1(n_1612),
.B2(n_1581),
.Y(n_1694)
);

CKINVDCx16_ASAP7_75t_R g1695 ( 
.A(n_1646),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1646),
.B(n_1608),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1663),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1656),
.Y(n_1698)
);

AOI22x1_ASAP7_75t_L g1699 ( 
.A1(n_1662),
.A2(n_1392),
.B1(n_1349),
.B2(n_1610),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1636),
.Y(n_1700)
);

CKINVDCx16_ASAP7_75t_R g1701 ( 
.A(n_1646),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1635),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1668),
.B(n_1664),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1669),
.B(n_1624),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1670),
.B(n_1635),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1677),
.B(n_1630),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1686),
.B(n_1652),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1674),
.Y(n_1708)
);

AOI21xp33_ASAP7_75t_L g1709 ( 
.A1(n_1682),
.A2(n_1662),
.B(n_1666),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1674),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1675),
.B(n_1660),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1676),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1680),
.B(n_1651),
.Y(n_1713)
);

OAI21xp33_ASAP7_75t_L g1714 ( 
.A1(n_1687),
.A2(n_1665),
.B(n_1666),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1676),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_SL g1716 ( 
.A(n_1681),
.B(n_1666),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1678),
.Y(n_1717)
);

NOR2x1_ASAP7_75t_L g1718 ( 
.A(n_1693),
.B(n_1610),
.Y(n_1718)
);

OAI21xp5_ASAP7_75t_L g1719 ( 
.A1(n_1673),
.A2(n_1692),
.B(n_1694),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1678),
.Y(n_1720)
);

OAI32xp33_ASAP7_75t_L g1721 ( 
.A1(n_1695),
.A2(n_1567),
.A3(n_1569),
.B1(n_1570),
.B2(n_1642),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1675),
.B(n_1657),
.Y(n_1722)
);

CKINVDCx14_ASAP7_75t_R g1723 ( 
.A(n_1672),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1683),
.Y(n_1724)
);

AOI322xp5_ASAP7_75t_L g1725 ( 
.A1(n_1685),
.A2(n_1554),
.A3(n_1553),
.B1(n_1552),
.B2(n_1551),
.C1(n_1558),
.C2(n_1549),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1700),
.B(n_1616),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1683),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1693),
.A2(n_1642),
.B1(n_1442),
.B2(n_1414),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1723),
.B(n_1702),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1705),
.B(n_1695),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1704),
.B(n_1706),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1723),
.B(n_1701),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1705),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1708),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1718),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1716),
.A2(n_1693),
.B1(n_1679),
.B2(n_1684),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1713),
.B(n_1698),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1719),
.B(n_1684),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1709),
.B(n_1700),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1710),
.Y(n_1740)
);

NAND2x1_ASAP7_75t_L g1741 ( 
.A(n_1712),
.B(n_1671),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1715),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1717),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1703),
.B(n_1702),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1716),
.B(n_1698),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1722),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1720),
.Y(n_1747)
);

INVx1_ASAP7_75t_SL g1748 ( 
.A(n_1707),
.Y(n_1748)
);

OAI21xp5_ASAP7_75t_SL g1749 ( 
.A1(n_1736),
.A2(n_1714),
.B(n_1728),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1733),
.B(n_1724),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1733),
.B(n_1727),
.Y(n_1751)
);

AOI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1732),
.A2(n_1721),
.B(n_1728),
.Y(n_1752)
);

AOI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1730),
.A2(n_1726),
.B(n_1711),
.Y(n_1753)
);

AOI221xp5_ASAP7_75t_L g1754 ( 
.A1(n_1745),
.A2(n_1697),
.B1(n_1671),
.B2(n_1679),
.C(n_1685),
.Y(n_1754)
);

OAI211xp5_ASAP7_75t_SL g1755 ( 
.A1(n_1729),
.A2(n_1730),
.B(n_1744),
.C(n_1748),
.Y(n_1755)
);

AOI221xp5_ASAP7_75t_L g1756 ( 
.A1(n_1739),
.A2(n_1697),
.B1(n_1688),
.B2(n_1696),
.C(n_1690),
.Y(n_1756)
);

NAND4xp25_ASAP7_75t_L g1757 ( 
.A(n_1738),
.B(n_1725),
.C(n_1696),
.D(n_1667),
.Y(n_1757)
);

O2A1O1Ixp33_ASAP7_75t_L g1758 ( 
.A1(n_1735),
.A2(n_1741),
.B(n_1738),
.C(n_1743),
.Y(n_1758)
);

OAI21xp33_ASAP7_75t_SL g1759 ( 
.A1(n_1735),
.A2(n_1691),
.B(n_1690),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1743),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1760),
.Y(n_1761)
);

NAND4xp75_ASAP7_75t_L g1762 ( 
.A(n_1752),
.B(n_1734),
.C(n_1740),
.D(n_1742),
.Y(n_1762)
);

NAND3xp33_ASAP7_75t_L g1763 ( 
.A(n_1755),
.B(n_1731),
.C(n_1746),
.Y(n_1763)
);

NOR2x1_ASAP7_75t_L g1764 ( 
.A(n_1758),
.B(n_1747),
.Y(n_1764)
);

NOR2x1p5_ASAP7_75t_SL g1765 ( 
.A(n_1749),
.B(n_1747),
.Y(n_1765)
);

INVxp33_ASAP7_75t_L g1766 ( 
.A(n_1757),
.Y(n_1766)
);

INVxp67_ASAP7_75t_L g1767 ( 
.A(n_1753),
.Y(n_1767)
);

NAND4xp25_ASAP7_75t_SL g1768 ( 
.A(n_1754),
.B(n_1731),
.C(n_1737),
.D(n_1667),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1756),
.B(n_1737),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1750),
.B(n_1689),
.Y(n_1770)
);

AOI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1763),
.A2(n_1759),
.B(n_1751),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1770),
.B(n_1691),
.Y(n_1772)
);

NOR2x1_ASAP7_75t_L g1773 ( 
.A(n_1764),
.B(n_1762),
.Y(n_1773)
);

NAND3xp33_ASAP7_75t_L g1774 ( 
.A(n_1767),
.B(n_1699),
.C(n_1569),
.Y(n_1774)
);

NAND4xp25_ASAP7_75t_SL g1775 ( 
.A(n_1769),
.B(n_1699),
.C(n_1611),
.D(n_1622),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1772),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1773),
.Y(n_1777)
);

NOR2xp67_ASAP7_75t_L g1778 ( 
.A(n_1774),
.B(n_1768),
.Y(n_1778)
);

AOI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1775),
.A2(n_1766),
.B1(n_1761),
.B2(n_1765),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_SL g1780 ( 
.A(n_1771),
.B(n_1611),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1772),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1776),
.Y(n_1782)
);

OAI221xp5_ASAP7_75t_SL g1783 ( 
.A1(n_1779),
.A2(n_1446),
.B1(n_1622),
.B2(n_1580),
.C(n_1576),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1781),
.B(n_1576),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1777),
.B(n_1593),
.Y(n_1785)
);

OAI222xp33_ASAP7_75t_L g1786 ( 
.A1(n_1780),
.A2(n_1569),
.B1(n_1567),
.B2(n_1348),
.C1(n_1570),
.C2(n_1617),
.Y(n_1786)
);

AOI21xp5_ASAP7_75t_SL g1787 ( 
.A1(n_1782),
.A2(n_1778),
.B(n_1334),
.Y(n_1787)
);

HB1xp67_ASAP7_75t_L g1788 ( 
.A(n_1785),
.Y(n_1788)
);

INVx4_ASAP7_75t_L g1789 ( 
.A(n_1784),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1789),
.A2(n_1783),
.B1(n_1786),
.B2(n_1593),
.Y(n_1790)
);

NOR4xp75_ASAP7_75t_L g1791 ( 
.A(n_1790),
.B(n_1787),
.C(n_1788),
.D(n_1334),
.Y(n_1791)
);

OAI21xp33_ASAP7_75t_L g1792 ( 
.A1(n_1791),
.A2(n_1580),
.B(n_1617),
.Y(n_1792)
);

AOI221x1_ASAP7_75t_L g1793 ( 
.A1(n_1791),
.A2(n_1619),
.B1(n_1618),
.B2(n_1570),
.C(n_1348),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1793),
.Y(n_1794)
);

AOI22x1_ASAP7_75t_L g1795 ( 
.A1(n_1792),
.A2(n_1305),
.B1(n_1351),
.B2(n_1619),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1794),
.B(n_1618),
.Y(n_1796)
);

OAI21xp5_ASAP7_75t_SL g1797 ( 
.A1(n_1796),
.A2(n_1795),
.B(n_1351),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1797),
.Y(n_1798)
);

AOI22xp33_ASAP7_75t_L g1799 ( 
.A1(n_1798),
.A2(n_1305),
.B1(n_1351),
.B2(n_1331),
.Y(n_1799)
);

AOI211xp5_ASAP7_75t_L g1800 ( 
.A1(n_1799),
.A2(n_1446),
.B(n_1351),
.C(n_1580),
.Y(n_1800)
);


endmodule