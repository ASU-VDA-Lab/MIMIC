module real_aes_1039_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_227;
wire n_564;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_478;
wire n_356;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_250;
wire n_85;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_552;
wire n_402;
wire n_87;
wire n_171;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g541 ( .A(n_0), .Y(n_541) );
AO22x2_ASAP7_75t_L g103 ( .A1(n_1), .A2(n_56), .B1(n_93), .B2(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g181 ( .A(n_2), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g153 ( .A1(n_3), .A2(n_63), .B1(n_154), .B2(n_160), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_4), .B(n_224), .Y(n_320) );
INVx1_ASAP7_75t_L g233 ( .A(n_5), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_6), .Y(n_124) );
AO22x2_ASAP7_75t_L g100 ( .A1(n_7), .A2(n_18), .B1(n_93), .B2(n_101), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_8), .Y(n_250) );
INVx2_ASAP7_75t_L g197 ( .A(n_9), .Y(n_197) );
INVx1_ASAP7_75t_L g329 ( .A(n_10), .Y(n_329) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_11), .Y(n_131) );
AOI22xp5_ASAP7_75t_L g143 ( .A1(n_12), .A2(n_70), .B1(n_144), .B2(n_149), .Y(n_143) );
INVx1_ASAP7_75t_L g326 ( .A(n_13), .Y(n_326) );
INVx1_ASAP7_75t_SL g291 ( .A(n_14), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_15), .B(n_212), .Y(n_312) );
AOI33xp33_ASAP7_75t_L g262 ( .A1(n_16), .A2(n_42), .A3(n_202), .B1(n_210), .B2(n_263), .B3(n_264), .Y(n_262) );
INVx1_ASAP7_75t_L g242 ( .A(n_17), .Y(n_242) );
OAI221xp5_ASAP7_75t_L g549 ( .A1(n_18), .A2(n_56), .B1(n_59), .B2(n_550), .C(n_552), .Y(n_549) );
OA21x2_ASAP7_75t_L g196 ( .A1(n_19), .A2(n_71), .B(n_197), .Y(n_196) );
OR2x2_ASAP7_75t_L g225 ( .A(n_19), .B(n_71), .Y(n_225) );
AND2x2_ASAP7_75t_L g85 ( .A(n_20), .B(n_86), .Y(n_85) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_21), .B(n_220), .Y(n_288) );
INVx3_ASAP7_75t_L g93 ( .A(n_22), .Y(n_93) );
OAI22xp5_ASAP7_75t_SL g533 ( .A1(n_23), .A2(n_38), .B1(n_534), .B2(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g535 ( .A(n_23), .Y(n_535) );
INVx1_ASAP7_75t_SL g94 ( .A(n_24), .Y(n_94) );
AO22x1_ASAP7_75t_L g105 ( .A1(n_25), .A2(n_49), .B1(n_106), .B2(n_112), .Y(n_105) );
INVx1_ASAP7_75t_L g183 ( .A(n_26), .Y(n_183) );
AND2x2_ASAP7_75t_L g218 ( .A(n_26), .B(n_181), .Y(n_218) );
AND2x2_ASAP7_75t_L g223 ( .A(n_26), .B(n_204), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g245 ( .A(n_27), .Y(n_245) );
OAI22xp5_ASAP7_75t_SL g79 ( .A1(n_28), .A2(n_80), .B1(n_81), .B2(n_177), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_28), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_29), .B(n_220), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g305 ( .A1(n_30), .A2(n_195), .B1(n_224), .B2(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_31), .B(n_314), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g164 ( .A1(n_32), .A2(n_41), .B1(n_165), .B2(n_168), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_33), .B(n_212), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_33), .A2(n_37), .B1(n_538), .B2(n_539), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_33), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g171 ( .A1(n_34), .A2(n_35), .B1(n_172), .B2(n_175), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_36), .B(n_230), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_37), .B(n_212), .Y(n_234) );
INVx1_ASAP7_75t_L g539 ( .A(n_37), .Y(n_539) );
INVx1_ASAP7_75t_L g534 ( .A(n_38), .Y(n_534) );
AO22x2_ASAP7_75t_L g96 ( .A1(n_39), .A2(n_59), .B1(n_93), .B2(n_97), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_40), .Y(n_309) );
INVx1_ASAP7_75t_L g556 ( .A(n_42), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_42), .A2(n_557), .B1(n_563), .B2(n_564), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_43), .B(n_212), .Y(n_274) );
INVx1_ASAP7_75t_L g206 ( .A(n_44), .Y(n_206) );
INVx1_ASAP7_75t_L g214 ( .A(n_44), .Y(n_214) );
AND2x2_ASAP7_75t_L g275 ( .A(n_45), .B(n_276), .Y(n_275) );
AOI221xp5_ASAP7_75t_L g231 ( .A1(n_46), .A2(n_61), .B1(n_200), .B2(n_220), .C(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_47), .B(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g95 ( .A(n_48), .Y(n_95) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_50), .B(n_195), .Y(n_252) );
AOI21xp5_ASAP7_75t_SL g199 ( .A1(n_51), .A2(n_200), .B(n_207), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_52), .A2(n_543), .B1(n_544), .B2(n_545), .Y(n_542) );
INVx1_ASAP7_75t_L g544 ( .A(n_52), .Y(n_544) );
INVx1_ASAP7_75t_L g323 ( .A(n_53), .Y(n_323) );
INVx1_ASAP7_75t_L g273 ( .A(n_54), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_55), .A2(n_200), .B(n_272), .Y(n_271) );
INVxp33_ASAP7_75t_L g554 ( .A(n_56), .Y(n_554) );
INVx1_ASAP7_75t_L g204 ( .A(n_57), .Y(n_204) );
INVx1_ASAP7_75t_L g216 ( .A(n_57), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_58), .Y(n_117) );
INVxp67_ASAP7_75t_L g553 ( .A(n_59), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_60), .B(n_220), .Y(n_265) );
INVx1_ASAP7_75t_L g570 ( .A(n_60), .Y(n_570) );
AND2x2_ASAP7_75t_L g293 ( .A(n_62), .B(n_194), .Y(n_293) );
INVx1_ASAP7_75t_L g324 ( .A(n_64), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_65), .A2(n_200), .B(n_290), .Y(n_289) );
A2O1A1Ixp33_ASAP7_75t_L g310 ( .A1(n_66), .A2(n_200), .B(n_257), .C(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_SL g193 ( .A(n_67), .B(n_194), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_68), .A2(n_200), .B1(n_260), .B2(n_261), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_69), .Y(n_137) );
INVx1_ASAP7_75t_L g208 ( .A(n_72), .Y(n_208) );
INVx1_ASAP7_75t_L g543 ( .A(n_73), .Y(n_543) );
AND2x2_ASAP7_75t_L g266 ( .A(n_74), .B(n_194), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_75), .A2(n_240), .B(n_241), .C(n_244), .Y(n_239) );
BUFx2_ASAP7_75t_SL g551 ( .A(n_76), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_77), .B(n_212), .Y(n_211) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_178), .B1(n_184), .B2(n_526), .C(n_528), .Y(n_78) );
OAI222xp33_ASAP7_75t_L g528 ( .A1(n_80), .A2(n_81), .B1(n_529), .B2(n_562), .C1(n_566), .C2(n_570), .Y(n_528) );
CKINVDCx16_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
NAND2xp5_ASAP7_75t_L g83 ( .A(n_84), .B(n_141), .Y(n_83) );
NOR4xp75_ASAP7_75t_L g84 ( .A(n_85), .B(n_105), .C(n_116), .D(n_130), .Y(n_84) );
INVx2_ASAP7_75t_SL g86 ( .A(n_87), .Y(n_86) );
BUFx2_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx6_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
AND2x2_ASAP7_75t_L g89 ( .A(n_90), .B(n_98), .Y(n_89) );
AND2x4_ASAP7_75t_L g127 ( .A(n_90), .B(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g139 ( .A(n_90), .B(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g90 ( .A(n_91), .B(n_96), .Y(n_90) );
AND2x2_ASAP7_75t_L g110 ( .A(n_91), .B(n_111), .Y(n_110) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_91), .Y(n_115) );
INVx2_ASAP7_75t_L g136 ( .A(n_91), .Y(n_136) );
OAI22x1_ASAP7_75t_L g91 ( .A1(n_92), .A2(n_93), .B1(n_94), .B2(n_95), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g97 ( .A(n_93), .Y(n_97) );
INVx2_ASAP7_75t_L g101 ( .A(n_93), .Y(n_101) );
INVx1_ASAP7_75t_L g104 ( .A(n_93), .Y(n_104) );
INVx2_ASAP7_75t_L g111 ( .A(n_96), .Y(n_111) );
AND2x2_ASAP7_75t_L g135 ( .A(n_96), .B(n_136), .Y(n_135) );
BUFx2_ASAP7_75t_L g152 ( .A(n_96), .Y(n_152) );
AND2x4_ASAP7_75t_L g158 ( .A(n_98), .B(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g167 ( .A(n_98), .B(n_135), .Y(n_167) );
AND2x4_ASAP7_75t_L g174 ( .A(n_98), .B(n_110), .Y(n_174) );
AND2x4_ASAP7_75t_L g98 ( .A(n_99), .B(n_102), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
AND2x4_ASAP7_75t_L g109 ( .A(n_100), .B(n_102), .Y(n_109) );
AND2x2_ASAP7_75t_L g114 ( .A(n_100), .B(n_103), .Y(n_114) );
INVx1_ASAP7_75t_L g123 ( .A(n_100), .Y(n_123) );
INVxp67_ASAP7_75t_L g140 ( .A(n_102), .Y(n_140) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_L g122 ( .A(n_103), .B(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
AND2x4_ASAP7_75t_L g134 ( .A(n_109), .B(n_135), .Y(n_134) );
AND2x4_ASAP7_75t_L g170 ( .A(n_109), .B(n_159), .Y(n_170) );
AND2x2_ASAP7_75t_L g121 ( .A(n_110), .B(n_122), .Y(n_121) );
AND2x4_ASAP7_75t_L g159 ( .A(n_111), .B(n_136), .Y(n_159) );
BUFx12f_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
AND2x4_ASAP7_75t_L g151 ( .A(n_114), .B(n_152), .Y(n_151) );
AND2x4_ASAP7_75t_L g176 ( .A(n_114), .B(n_159), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_118), .B1(n_124), .B2(n_125), .Y(n_116) );
INVx2_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
INVx4_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_L g148 ( .A(n_122), .B(n_135), .Y(n_148) );
AND2x4_ASAP7_75t_L g162 ( .A(n_122), .B(n_159), .Y(n_162) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_123), .Y(n_129) );
BUFx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OAI22xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_132), .B1(n_137), .B2(n_138), .Y(n_130) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx6_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_142), .B(n_163), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_153), .Y(n_142) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx5_ASAP7_75t_SL g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx4_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx8_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx8_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_164), .B(n_171), .Y(n_163) );
INVx2_ASAP7_75t_SL g165 ( .A(n_166), .Y(n_165) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx6_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
BUFx2_ASAP7_75t_SL g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
OR2x2_ASAP7_75t_SL g179 ( .A(n_180), .B(n_182), .Y(n_179) );
AND2x2_ASAP7_75t_L g221 ( .A(n_180), .B(n_210), .Y(n_221) );
INVx1_ASAP7_75t_L g555 ( .A(n_180), .Y(n_555) );
HB1xp67_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g205 ( .A(n_181), .B(n_206), .Y(n_205) );
AND3x1_ASAP7_75t_SL g548 ( .A(n_182), .B(n_549), .C(n_555), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_182), .B(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NOR2x1p5_ASAP7_75t_L g201 ( .A(n_183), .B(n_202), .Y(n_201) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
BUFx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NAND3x1_ASAP7_75t_L g186 ( .A(n_187), .B(n_416), .C(n_481), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_370), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_315), .B(n_343), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_190), .B(n_278), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_191), .B(n_226), .Y(n_190) );
AOI21xp33_ASAP7_75t_L g417 ( .A1(n_191), .A2(n_418), .B(n_429), .Y(n_417) );
AND2x2_ASAP7_75t_SL g452 ( .A(n_191), .B(n_359), .Y(n_452) );
AND2x2_ASAP7_75t_L g467 ( .A(n_191), .B(n_468), .Y(n_467) );
OR2x6_ASAP7_75t_L g477 ( .A(n_191), .B(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g479 ( .A(n_191), .B(n_469), .Y(n_479) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g353 ( .A(n_192), .Y(n_353) );
AND2x2_ASAP7_75t_L g366 ( .A(n_192), .B(n_367), .Y(n_366) );
INVx4_ASAP7_75t_L g385 ( .A(n_192), .Y(n_385) );
AND2x2_ASAP7_75t_L g388 ( .A(n_192), .B(n_304), .Y(n_388) );
NOR2x1_ASAP7_75t_SL g391 ( .A(n_192), .B(n_319), .Y(n_391) );
AND2x4_ASAP7_75t_L g403 ( .A(n_192), .B(n_401), .Y(n_403) );
OR2x2_ASAP7_75t_L g413 ( .A(n_192), .B(n_285), .Y(n_413) );
NAND2xp5_ASAP7_75t_SL g430 ( .A(n_192), .B(n_425), .Y(n_430) );
OR2x6_ASAP7_75t_L g192 ( .A(n_193), .B(n_198), .Y(n_192) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_194), .A2(n_239), .B1(n_245), .B2(n_246), .Y(n_238) );
INVx3_ASAP7_75t_L g246 ( .A(n_194), .Y(n_246) );
INVx4_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_195), .B(n_249), .Y(n_248) );
INVx3_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
BUFx4f_ASAP7_75t_L g230 ( .A(n_196), .Y(n_230) );
AND2x4_ASAP7_75t_L g224 ( .A(n_197), .B(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_SL g277 ( .A(n_197), .B(n_225), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_219), .B(n_224), .Y(n_198) );
INVxp67_ASAP7_75t_L g251 ( .A(n_200), .Y(n_251) );
AND2x4_ASAP7_75t_L g200 ( .A(n_201), .B(n_205), .Y(n_200) );
INVx1_ASAP7_75t_L g264 ( .A(n_202), .Y(n_264) );
INVx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
OR2x6_ASAP7_75t_L g209 ( .A(n_203), .B(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x6_ASAP7_75t_L g328 ( .A(n_204), .B(n_213), .Y(n_328) );
INVx2_ASAP7_75t_L g210 ( .A(n_206), .Y(n_210) );
AND2x4_ASAP7_75t_L g331 ( .A(n_206), .B(n_215), .Y(n_331) );
O2A1O1Ixp33_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_211), .C(n_217), .Y(n_207) );
O2A1O1Ixp33_ASAP7_75t_SL g232 ( .A1(n_209), .A2(n_217), .B(n_233), .C(n_234), .Y(n_232) );
INVxp67_ASAP7_75t_L g240 ( .A(n_209), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_L g272 ( .A1(n_209), .A2(n_217), .B(n_273), .C(n_274), .Y(n_272) );
O2A1O1Ixp33_ASAP7_75t_SL g290 ( .A1(n_209), .A2(n_217), .B(n_291), .C(n_292), .Y(n_290) );
INVx2_ASAP7_75t_L g314 ( .A(n_209), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_209), .A2(n_243), .B1(n_323), .B2(n_324), .Y(n_322) );
INVxp33_ASAP7_75t_L g263 ( .A(n_210), .Y(n_263) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_210), .Y(n_568) );
INVx1_ASAP7_75t_L g243 ( .A(n_212), .Y(n_243) );
AND2x4_ASAP7_75t_L g212 ( .A(n_213), .B(n_215), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g260 ( .A(n_217), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_217), .A2(n_312), .B(n_313), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_217), .B(n_224), .Y(n_332) );
INVx5_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_218), .Y(n_244) );
INVx1_ASAP7_75t_L g253 ( .A(n_220), .Y(n_253) );
AND2x4_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
INVx1_ASAP7_75t_L g307 ( .A(n_221), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_222), .Y(n_308) );
BUFx3_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_226), .A2(n_359), .B1(n_454), .B2(n_455), .Y(n_453) );
INVx1_ASAP7_75t_SL g497 ( .A(n_226), .Y(n_497) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_254), .Y(n_226) );
INVx2_ASAP7_75t_L g428 ( .A(n_227), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_227), .B(n_374), .Y(n_500) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_236), .Y(n_227) );
BUFx3_ASAP7_75t_L g346 ( .A(n_228), .Y(n_346) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g339 ( .A(n_229), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_229), .B(n_256), .Y(n_361) );
AND2x4_ASAP7_75t_L g378 ( .A(n_229), .B(n_379), .Y(n_378) );
INVxp67_ASAP7_75t_L g394 ( .A(n_229), .Y(n_394) );
INVx2_ASAP7_75t_L g451 ( .A(n_229), .Y(n_451) );
OA21x2_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_235), .Y(n_229) );
INVx2_ASAP7_75t_SL g257 ( .A(n_230), .Y(n_257) );
AND2x2_ASAP7_75t_L g369 ( .A(n_236), .B(n_335), .Y(n_369) );
NOR2xp67_ASAP7_75t_L g415 ( .A(n_236), .B(n_338), .Y(n_415) );
AND2x2_ASAP7_75t_L g434 ( .A(n_236), .B(n_338), .Y(n_434) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g296 ( .A(n_237), .Y(n_296) );
INVx1_ASAP7_75t_L g377 ( .A(n_237), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_237), .B(n_268), .Y(n_396) );
AND2x4_ASAP7_75t_L g450 ( .A(n_237), .B(n_451), .Y(n_450) );
OR2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_247), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
AO21x2_ASAP7_75t_L g268 ( .A1(n_246), .A2(n_269), .B(n_275), .Y(n_268) );
AO21x2_ASAP7_75t_L g338 ( .A1(n_246), .A2(n_269), .B(n_275), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_251), .B1(n_252), .B2(n_253), .Y(n_247) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_253), .Y(n_527) );
INVx1_ASAP7_75t_L g409 ( .A(n_254), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_254), .B(n_467), .Y(n_466) );
AND2x4_ASAP7_75t_L g254 ( .A(n_255), .B(n_267), .Y(n_254) );
AND2x2_ASAP7_75t_L g393 ( .A(n_255), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g433 ( .A(n_255), .Y(n_433) );
AND2x2_ASAP7_75t_L g438 ( .A(n_255), .B(n_338), .Y(n_438) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_256), .B(n_268), .Y(n_298) );
AO21x2_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_258), .B(n_266), .Y(n_256) );
AO21x2_ASAP7_75t_L g335 ( .A1(n_257), .A2(n_258), .B(n_266), .Y(n_335) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_259), .B(n_265), .Y(n_258) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx3_ASAP7_75t_L g374 ( .A(n_267), .Y(n_374) );
NAND2x1p5_ASAP7_75t_L g492 ( .A(n_267), .B(n_346), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_267), .B(n_296), .Y(n_513) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_268), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_276), .Y(n_286) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OAI21xp33_ASAP7_75t_SL g278 ( .A1(n_279), .A2(n_294), .B(n_299), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_281), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g351 ( .A(n_282), .Y(n_351) );
AND2x2_ASAP7_75t_L g365 ( .A(n_282), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g399 ( .A(n_282), .B(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g465 ( .A(n_282), .B(n_383), .Y(n_465) );
NOR3xp33_ASAP7_75t_L g511 ( .A(n_282), .B(n_512), .C(n_513), .Y(n_511) );
INVx3_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_283), .Y(n_342) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g358 ( .A(n_285), .Y(n_358) );
AND2x2_ASAP7_75t_L g364 ( .A(n_285), .B(n_319), .Y(n_364) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_285), .Y(n_375) );
AND2x2_ASAP7_75t_L g420 ( .A(n_285), .B(n_318), .Y(n_420) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_285), .Y(n_443) );
INVx1_ASAP7_75t_L g460 ( .A(n_285), .Y(n_460) );
AO21x2_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_287), .B(n_293), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx1_ASAP7_75t_L g502 ( .A(n_294), .Y(n_502) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_295), .B(n_373), .Y(n_474) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g336 ( .A(n_296), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AOI211x1_ASAP7_75t_L g370 ( .A1(n_300), .A2(n_371), .B(n_380), .C(n_397), .Y(n_370) );
INVx2_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_SL g363 ( .A(n_301), .B(n_364), .Y(n_363) );
AND2x4_ASAP7_75t_L g423 ( .A(n_301), .B(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g359 ( .A(n_303), .B(n_318), .Y(n_359) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x4_ASAP7_75t_L g317 ( .A(n_304), .B(n_318), .Y(n_317) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_304), .Y(n_384) );
INVx1_ASAP7_75t_L g401 ( .A(n_304), .Y(n_401) );
AND2x2_ASAP7_75t_L g469 ( .A(n_304), .B(n_319), .Y(n_469) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_310), .Y(n_304) );
NOR3xp33_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .C(n_309), .Y(n_306) );
INVxp67_ASAP7_75t_L g569 ( .A(n_308), .Y(n_569) );
OAI21xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_333), .B(n_340), .Y(n_315) );
NOR2x1_ASAP7_75t_L g488 ( .A(n_316), .B(n_385), .Y(n_488) );
INVx2_ASAP7_75t_L g520 ( .A(n_316), .Y(n_520) );
INVx4_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g352 ( .A(n_317), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g425 ( .A(n_318), .Y(n_425) );
INVx3_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g367 ( .A(n_319), .Y(n_367) );
AND2x4_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
OAI21xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_325), .B(n_332), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_327), .B1(n_329), .B2(n_330), .Y(n_325) );
INVxp67_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVxp67_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
OR2x2_ASAP7_75t_L g427 ( .A(n_334), .B(n_428), .Y(n_427) );
NAND2x1_ASAP7_75t_SL g449 ( .A(n_334), .B(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x4_ASAP7_75t_L g349 ( .A(n_335), .B(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g379 ( .A(n_335), .Y(n_379) );
INVx1_ASAP7_75t_L g503 ( .A(n_336), .Y(n_503) );
AND2x2_ASAP7_75t_L g368 ( .A(n_337), .B(n_369), .Y(n_368) );
NOR2x1_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx2_ASAP7_75t_L g350 ( .A(n_338), .Y(n_350) );
INVxp33_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g407 ( .A(n_342), .B(n_400), .Y(n_407) );
OAI211xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_347), .B(n_354), .C(n_362), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g431 ( .A(n_345), .B(n_432), .Y(n_431) );
NOR2xp67_ASAP7_75t_SL g436 ( .A(n_345), .B(n_437), .Y(n_436) );
INVx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_346), .B(n_433), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g347 ( .A(n_348), .B(n_352), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .Y(n_348) );
AND2x2_ASAP7_75t_L g480 ( .A(n_349), .B(n_450), .Y(n_480) );
AOI222xp33_ASAP7_75t_L g498 ( .A1(n_352), .A2(n_499), .B1(n_501), .B2(n_504), .C1(n_505), .C2(n_508), .Y(n_498) );
INVx1_ASAP7_75t_L g462 ( .A(n_353), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_360), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_358), .Y(n_389) );
AND2x4_ASAP7_75t_SL g424 ( .A(n_358), .B(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g478 ( .A(n_359), .Y(n_478) );
AND2x2_ASAP7_75t_L g523 ( .A(n_359), .B(n_375), .Y(n_523) );
AND2x2_ASAP7_75t_L g404 ( .A(n_360), .B(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g517 ( .A(n_361), .B(n_396), .Y(n_517) );
OAI21xp33_ASAP7_75t_SL g362 ( .A1(n_363), .A2(n_365), .B(n_368), .Y(n_362) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_363), .A2(n_383), .B(n_424), .Y(n_484) );
AND2x2_ASAP7_75t_L g508 ( .A(n_364), .B(n_385), .Y(n_508) );
NOR2xp33_ASAP7_75t_SL g518 ( .A(n_364), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g456 ( .A(n_367), .Y(n_456) );
NOR2x1_ASAP7_75t_L g461 ( .A(n_367), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g491 ( .A(n_369), .Y(n_491) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_376), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
AND2x2_ASAP7_75t_L g494 ( .A(n_374), .B(n_378), .Y(n_494) );
BUFx2_ASAP7_75t_L g382 ( .A(n_375), .Y(n_382) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
INVx1_ASAP7_75t_L g405 ( .A(n_377), .Y(n_405) );
INVx2_ASAP7_75t_L g411 ( .A(n_377), .Y(n_411) );
AND2x2_ASAP7_75t_L g447 ( .A(n_377), .B(n_438), .Y(n_447) );
AND2x4_ASAP7_75t_L g414 ( .A(n_378), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g454 ( .A(n_378), .B(n_411), .Y(n_454) );
AND2x2_ASAP7_75t_L g505 ( .A(n_378), .B(n_506), .Y(n_505) );
AOI31xp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_386), .A3(n_390), .B(n_392), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
AND2x2_ASAP7_75t_L g402 ( .A(n_382), .B(n_403), .Y(n_402) );
AND2x4_ASAP7_75t_SL g383 ( .A(n_384), .B(n_385), .Y(n_383) );
AND2x4_ASAP7_75t_L g400 ( .A(n_385), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_388), .A2(n_440), .B1(n_471), .B2(n_474), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_388), .B(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g525 ( .A(n_388), .B(n_441), .Y(n_525) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g440 ( .A(n_391), .B(n_441), .Y(n_440) );
NAND2x1p5_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
AND2x2_ASAP7_75t_L g463 ( .A(n_393), .B(n_434), .Y(n_463) );
INVx1_ASAP7_75t_L g473 ( .A(n_395), .Y(n_473) );
INVx2_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_406), .Y(n_397) );
OAI21xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_402), .B(n_404), .Y(n_398) );
INVx1_ASAP7_75t_L g496 ( .A(n_399), .Y(n_496) );
AND2x2_ASAP7_75t_L g504 ( .A(n_400), .B(n_456), .Y(n_504) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_400), .Y(n_510) );
AND2x2_ASAP7_75t_L g455 ( .A(n_403), .B(n_456), .Y(n_455) );
AOI22xp33_ASAP7_75t_SL g406 ( .A1(n_407), .A2(n_408), .B1(n_412), .B2(n_414), .Y(n_406) );
NOR2xp33_ASAP7_75t_SL g408 ( .A(n_409), .B(n_410), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_409), .A2(n_428), .B1(n_522), .B2(n_524), .Y(n_521) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx2_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g421 ( .A(n_414), .Y(n_421) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_444), .Y(n_416) );
OAI21xp33_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_421), .B(n_422), .Y(n_418) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
OAI21xp33_ASAP7_75t_L g422 ( .A1(n_420), .A2(n_423), .B(n_426), .Y(n_422) );
AOI22xp33_ASAP7_75t_SL g446 ( .A1(n_423), .A2(n_447), .B1(n_448), .B2(n_452), .Y(n_446) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_431), .B1(n_435), .B2(n_439), .Y(n_429) );
INVx1_ASAP7_75t_L g464 ( .A(n_432), .Y(n_464) );
NAND2x1p5_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NOR2xp67_ASAP7_75t_L g444 ( .A(n_445), .B(n_457), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_453), .Y(n_445) );
INVx2_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
NAND2xp33_ASAP7_75t_SL g499 ( .A(n_449), .B(n_500), .Y(n_499) );
INVx3_ASAP7_75t_L g472 ( .A(n_450), .Y(n_472) );
INVx3_ASAP7_75t_L g486 ( .A(n_454), .Y(n_486) );
INVxp67_ASAP7_75t_L g515 ( .A(n_455), .Y(n_515) );
NAND4xp25_ASAP7_75t_L g457 ( .A(n_458), .B(n_466), .C(n_470), .D(n_475), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_463), .B1(n_464), .B2(n_465), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
AND2x2_ASAP7_75t_L g468 ( .A(n_460), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g516 ( .A(n_464), .Y(n_516) );
NAND2xp33_ASAP7_75t_SL g471 ( .A(n_472), .B(n_473), .Y(n_471) );
OAI21xp33_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_479), .B(n_480), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND3x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_498), .C(n_509), .Y(n_481) );
AOI221x1_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_485), .B1(n_487), .B2(n_489), .C(n_495), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND2xp33_ASAP7_75t_SL g489 ( .A(n_490), .B(n_493), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
NAND2xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AOI211xp5_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_511), .B(n_514), .C(n_521), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B1(n_517), .B2(n_518), .Y(n_514) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
CKINVDCx16_ASAP7_75t_R g526 ( .A(n_527), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_548), .B1(n_556), .B2(n_557), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g563 ( .A(n_530), .Y(n_563) );
XOR2x2_ASAP7_75t_SL g530 ( .A(n_531), .B(n_540), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .B1(n_536), .B2(n_537), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_533), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_537), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .B1(n_546), .B2(n_547), .Y(n_540) );
INVx1_ASAP7_75t_L g546 ( .A(n_541), .Y(n_546) );
CKINVDCx16_ASAP7_75t_R g547 ( .A(n_542), .Y(n_547) );
INVx1_ASAP7_75t_L g545 ( .A(n_543), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_548), .Y(n_565) );
INVxp67_ASAP7_75t_L g561 ( .A(n_549), .Y(n_561) );
CKINVDCx8_ASAP7_75t_R g550 ( .A(n_551), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
CKINVDCx16_ASAP7_75t_R g559 ( .A(n_555), .Y(n_559) );
AOI21xp33_ASAP7_75t_L g567 ( .A1(n_555), .A2(n_568), .B(n_569), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_558), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
endmodule