module fake_aes_1024_n_38 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_38);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_7), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
CKINVDCx16_ASAP7_75t_R g13 ( .A(n_10), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
INVx3_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_2), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_3), .Y(n_17) );
INVx1_ASAP7_75t_SL g18 ( .A(n_17), .Y(n_18) );
INVx2_ASAP7_75t_SL g19 ( .A(n_15), .Y(n_19) );
INVx3_ASAP7_75t_L g20 ( .A(n_15), .Y(n_20) );
HB1xp67_ASAP7_75t_L g21 ( .A(n_17), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_14), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_19), .B(n_13), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_19), .B(n_20), .Y(n_24) );
NOR2x1_ASAP7_75t_SL g25 ( .A(n_22), .B(n_14), .Y(n_25) );
BUFx2_ASAP7_75t_L g26 ( .A(n_21), .Y(n_26) );
OAI33xp33_ASAP7_75t_L g27 ( .A1(n_23), .A2(n_22), .A3(n_12), .B1(n_16), .B2(n_11), .B3(n_18), .Y(n_27) );
AOI33xp33_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_20), .A3(n_1), .B1(n_2), .B2(n_3), .B3(n_0), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_24), .Y(n_29) );
INVx2_ASAP7_75t_L g30 ( .A(n_29), .Y(n_30) );
AND2x2_ASAP7_75t_L g31 ( .A(n_29), .B(n_25), .Y(n_31) );
NOR2xp33_ASAP7_75t_L g32 ( .A(n_31), .B(n_27), .Y(n_32) );
AND2x2_ASAP7_75t_L g33 ( .A(n_30), .B(n_28), .Y(n_33) );
NAND4xp25_ASAP7_75t_L g34 ( .A(n_32), .B(n_15), .C(n_20), .D(n_8), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_33), .Y(n_35) );
NOR3xp33_ASAP7_75t_L g36 ( .A(n_34), .B(n_35), .C(n_20), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_36), .Y(n_37) );
AOI22xp33_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_4), .B1(n_6), .B2(n_9), .Y(n_38) );
endmodule