module real_jpeg_24123_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_249;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_105;
wire n_40;
wire n_173;
wire n_243;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_198;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_202;
wire n_213;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx8_ASAP7_75t_SL g64 ( 
.A(n_3),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_4),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_4),
.B(n_70),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_4),
.B(n_27),
.C(n_43),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_105),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_4),
.B(n_113),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_4),
.A2(n_24),
.B1(n_210),
.B2(n_213),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_5),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_48),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_5),
.A2(n_48),
.B1(n_65),
.B2(n_66),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_6),
.A2(n_35),
.B1(n_45),
.B2(n_46),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_6),
.A2(n_35),
.B1(n_65),
.B2(n_66),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_7),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_7),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_7),
.A2(n_60),
.B1(n_65),
.B2(n_66),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_7),
.A2(n_45),
.B1(n_46),
.B2(n_60),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_60),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_8),
.A2(n_58),
.B1(n_69),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_8),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_8),
.A2(n_65),
.B1(n_66),
.B2(n_72),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_72),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_8),
.A2(n_45),
.B1(n_46),
.B2(n_72),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_9),
.A2(n_32),
.B1(n_45),
.B2(n_46),
.Y(n_94)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

NAND3xp33_ASAP7_75t_L g107 ( 
.A(n_10),
.B(n_64),
.C(n_65),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_11),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_12),
.A2(n_65),
.B1(n_66),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_12),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_80),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_12),
.A2(n_58),
.B1(n_69),
.B2(n_80),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_12),
.A2(n_45),
.B1(n_46),
.B2(n_80),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_13),
.A2(n_59),
.B1(n_106),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_13),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_13),
.A2(n_65),
.B1(n_66),
.B2(n_117),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_117),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_117),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_15),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_147),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_146),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_119),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_20),
.B(n_119),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_83),
.C(n_96),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_21),
.B(n_83),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_55),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_22),
.B(n_56),
.C(n_73),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_23),
.B(n_40),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_33),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_24),
.A2(n_89),
.B(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_24),
.A2(n_86),
.B(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_24),
.A2(n_37),
.B1(n_203),
.B2(n_210),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_24),
.A2(n_33),
.B(n_89),
.Y(n_229)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_25),
.B(n_34),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_25),
.A2(n_31),
.B1(n_36),
.B2(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_25),
.A2(n_36),
.B1(n_202),
.B2(n_204),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_26),
.A2(n_27),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_26),
.B(n_216),
.Y(n_215)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_29),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_39),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_39),
.A2(n_90),
.B(n_102),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_44),
.B(n_49),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_41),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_41),
.B(n_54),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_41),
.A2(n_51),
.B1(n_189),
.B2(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_41),
.B(n_105),
.Y(n_208)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_42),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_44),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_45),
.A2(n_46),
.B1(n_76),
.B2(n_77),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_45),
.A2(n_77),
.B(n_225),
.C(n_227),
.Y(n_224)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_46),
.B(n_185),
.Y(n_184)
);

NOR3xp33_ASAP7_75t_L g227 ( 
.A(n_46),
.B(n_65),
.C(n_76),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_50),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_50),
.A2(n_128),
.B(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_50),
.A2(n_93),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_50),
.A2(n_93),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_51),
.A2(n_126),
.B(n_127),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_51),
.A2(n_248),
.B(n_249),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_73),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_61),
.B1(n_70),
.B2(n_71),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_57),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_63),
.B1(n_64),
.B2(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_59),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_61),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_61),
.A2(n_70),
.B1(n_158),
.B2(n_160),
.Y(n_157)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_68),
.Y(n_61)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_62),
.A2(n_115),
.B1(n_116),
.B2(n_118),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_63),
.A2(n_66),
.B(n_104),
.C(n_107),
.Y(n_103)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_66),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

HAxp5_ASAP7_75t_SL g226 ( 
.A(n_66),
.B(n_105),
.CON(n_226),
.SN(n_226)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_70),
.B(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_71),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_79),
.B(n_81),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_74),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_74),
.B(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_74),
.A2(n_110),
.B1(n_113),
.B2(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_74),
.A2(n_113),
.B1(n_175),
.B2(n_226),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_78),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_78),
.A2(n_111),
.B1(n_174),
.B2(n_176),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_79),
.B(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_91),
.B2(n_95),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_95),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_93),
.B(n_154),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_94),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_96),
.B(n_262),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_108),
.C(n_114),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_97),
.A2(n_98),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_99),
.A2(n_100),
.B1(n_103),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_103),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_104),
.A2(n_105),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_105),
.B(n_124),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_108),
.B(n_114),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_111),
.B(n_112),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_134),
.B(n_135),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_116),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_145),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_130),
.B1(n_143),
.B2(n_144),
.Y(n_120)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_125),
.B2(n_129),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_137),
.B1(n_138),
.B2(n_142),
.Y(n_132)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_177),
.B(n_259),
.C(n_263),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_164),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_149),
.B(n_164),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_161),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_151),
.B(n_152),
.C(n_161),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.C(n_157),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_155),
.Y(n_166)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.C(n_169),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_165),
.B(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_167),
.B(n_169),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.C(n_173),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_170),
.Y(n_243)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_173),
.B(n_242),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_258),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_253),
.B(n_257),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_237),
.B(n_252),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_220),
.B(n_236),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_199),
.B(n_219),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_190),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_190),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_186),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_191),
.B(n_194),
.C(n_197),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_192),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_198),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_206),
.B(n_218),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_205),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_205),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_211),
.B(n_217),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_209),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_235),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_235),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_230),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_231),
.C(n_232),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_228),
.B2(n_229),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_229),
.Y(n_246)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_234),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_239),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_244),
.B2(n_245),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_247),
.C(n_250),
.Y(n_256)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_250),
.B2(n_251),
.Y(n_245)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_246),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_247),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_256),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_260),
.B(n_261),
.Y(n_263)
);


endmodule