module fake_jpeg_5533_n_179 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_152;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_SL g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_25),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_34),
.Y(n_42)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_1),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_1),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_49),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_41),
.B1(n_32),
.B2(n_39),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_21),
.B1(n_33),
.B2(n_30),
.Y(n_74)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_56),
.Y(n_77)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_65),
.Y(n_90)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_60),
.Y(n_86)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_62),
.Y(n_93)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_22),
.B1(n_41),
.B2(n_31),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_64),
.A2(n_79),
.B1(n_1),
.B2(n_3),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_38),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_39),
.B(n_32),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_66),
.A2(n_3),
.B(n_4),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_38),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_72),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_54),
.A2(n_22),
.B1(n_21),
.B2(n_23),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_69),
.A2(n_78),
.B1(n_17),
.B2(n_2),
.Y(n_97)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_71),
.Y(n_95)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_30),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_40),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_27),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_76),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_27),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_41),
.B1(n_33),
.B2(n_35),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_56),
.A2(n_24),
.B1(n_40),
.B2(n_33),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_34),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_24),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_83),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_47),
.B(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_37),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_37),
.C(n_35),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_89),
.Y(n_109)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_76),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_SL g94 ( 
.A(n_58),
.B(n_19),
.C(n_26),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_96),
.C(n_71),
.Y(n_110)
);

AO21x1_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_18),
.B(n_16),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_99),
.B1(n_12),
.B2(n_6),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_75),
.B(n_6),
.Y(n_114)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

O2A1O1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_62),
.B1(n_61),
.B2(n_68),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_4),
.Y(n_104)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_83),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_84),
.Y(n_129)
);

NOR3xp33_ASAP7_75t_SL g106 ( 
.A(n_94),
.B(n_65),
.C(n_67),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_112),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_SL g108 ( 
.A1(n_100),
.A2(n_78),
.B(n_77),
.C(n_63),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_108),
.A2(n_115),
.B(n_90),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_110),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_92),
.B(n_102),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_60),
.B(n_59),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_91),
.A2(n_70),
.B1(n_68),
.B2(n_11),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_117),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_5),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_92),
.C(n_98),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_88),
.B(n_84),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_120),
.Y(n_134)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

INVxp33_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_108),
.A2(n_103),
.B1(n_98),
.B2(n_88),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_108),
.B1(n_96),
.B2(n_87),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_126),
.A2(n_128),
.B(n_137),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_106),
.C(n_112),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_113),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_105),
.B(n_118),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_130),
.B(n_109),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_115),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_110),
.C(n_108),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_89),
.B(n_96),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_116),
.Y(n_138)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_146),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_143),
.C(n_144),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_134),
.B(n_111),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_141),
.B(n_145),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_121),
.C(n_95),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_6),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_148),
.B(n_149),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_136),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_153),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_126),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_142),
.A2(n_123),
.B1(n_137),
.B2(n_125),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_156),
.A2(n_125),
.B1(n_128),
.B2(n_131),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_160),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_130),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_146),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_162),
.C(n_163),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_132),
.C(n_133),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_113),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_87),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_152),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_156),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_170),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_158),
.C(n_154),
.Y(n_171)
);

NOR2x1_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_155),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_174),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_164),
.C(n_73),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_173),
.A2(n_170),
.B(n_166),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_73),
.Y(n_174)
);

AOI31xp33_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_172),
.A3(n_167),
.B(n_73),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_175),
.C(n_8),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_7),
.Y(n_179)
);


endmodule