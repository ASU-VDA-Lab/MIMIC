module fake_netlist_5_458_n_1658 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1658);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1658;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_150;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_152;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_146;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1637;
wire n_1419;
wire n_338;
wire n_149;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_151;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_148;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_147;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g146 ( 
.A(n_32),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_23),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_94),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_0),
.Y(n_149)
);

INVxp67_ASAP7_75t_SL g150 ( 
.A(n_56),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_102),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_21),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_59),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_2),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_43),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_109),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_83),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_54),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_86),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_67),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_62),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_43),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_80),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_70),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_32),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_142),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_101),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_87),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_37),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_112),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_103),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_140),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_125),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_26),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_128),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_110),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_26),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_18),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_91),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_130),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_134),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_66),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_99),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_89),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_104),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_92),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_68),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_6),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_75),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_28),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_2),
.Y(n_191)
);

BUFx10_ASAP7_75t_L g192 ( 
.A(n_23),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_105),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_28),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_4),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_51),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_100),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_113),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_131),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_31),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_31),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_15),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_5),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_129),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_120),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_133),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_3),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_21),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_117),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_114),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_121),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_24),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_119),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_111),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_88),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_3),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_14),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_106),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_71),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_98),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_63),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_33),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_24),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_122),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_118),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_136),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_126),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_35),
.Y(n_228)
);

INVxp67_ASAP7_75t_SL g229 ( 
.A(n_33),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_116),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_11),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_135),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_18),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_84),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_5),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_115),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_27),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_93),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_12),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_27),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_123),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_50),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_20),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_40),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_55),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_47),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_65),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_85),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_10),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_29),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_95),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_132),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_13),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_13),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_46),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_17),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_141),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_78),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_29),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_60),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_1),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_48),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_44),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_45),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_41),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_81),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_14),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_137),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_49),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_36),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_145),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_11),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_61),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_76),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_69),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_38),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_38),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_96),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_6),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_90),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_44),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_12),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_127),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_72),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_107),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_0),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_19),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_57),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_58),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_74),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_15),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_52),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_97),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_82),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_139),
.Y(n_295)
);

BUFx8_ASAP7_75t_SL g296 ( 
.A(n_124),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_45),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_191),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_185),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_224),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_191),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_280),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_296),
.Y(n_303)
);

INVxp33_ASAP7_75t_SL g304 ( 
.A(n_149),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_191),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_219),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_191),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_191),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_194),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_194),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_194),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_194),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_194),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_192),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_162),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_162),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_179),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_181),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_182),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_231),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_149),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_192),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_231),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_186),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_192),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_208),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_199),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_146),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_263),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_147),
.Y(n_330)
);

INVxp33_ASAP7_75t_SL g331 ( 
.A(n_155),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_208),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_152),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_190),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_187),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_189),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_148),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_195),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_203),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_193),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_197),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_212),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_209),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_204),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_216),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_225),
.Y(n_346)
);

INVxp33_ASAP7_75t_L g347 ( 
.A(n_228),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_156),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_205),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_210),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_258),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_211),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_243),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_168),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_175),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_244),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_168),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_259),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_262),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_285),
.Y(n_360)
);

INVxp33_ASAP7_75t_SL g361 ( 
.A(n_155),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_272),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_279),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g364 ( 
.A(n_263),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_282),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_287),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_165),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_165),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_348),
.B(n_198),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_298),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_354),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_298),
.Y(n_372)
);

OA21x2_ASAP7_75t_L g373 ( 
.A1(n_301),
.A2(n_206),
.B(n_159),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_337),
.B(n_198),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_354),
.Y(n_375)
);

NOR2x1_ASAP7_75t_L g376 ( 
.A(n_301),
.B(n_159),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_354),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_354),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_354),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g380 ( 
.A(n_321),
.B(n_229),
.Y(n_380)
);

NAND2xp33_ASAP7_75t_L g381 ( 
.A(n_354),
.B(n_168),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_305),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_299),
.B(n_154),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_357),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_327),
.A2(n_291),
.B1(n_188),
.B2(n_256),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_305),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_357),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_307),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_357),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_357),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_357),
.Y(n_391)
);

AND2x6_ASAP7_75t_L g392 ( 
.A(n_357),
.B(n_168),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_317),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_307),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_306),
.B(n_294),
.Y(n_395)
);

BUFx12f_ASAP7_75t_L g396 ( 
.A(n_303),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_308),
.B(n_294),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_308),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_337),
.Y(n_399)
);

OAI21x1_ASAP7_75t_L g400 ( 
.A1(n_309),
.A2(n_220),
.B(n_206),
.Y(n_400)
);

NAND2xp33_ASAP7_75t_R g401 ( 
.A(n_304),
.B(n_169),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_309),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_318),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_310),
.Y(n_404)
);

AND2x4_ASAP7_75t_L g405 ( 
.A(n_337),
.B(n_220),
.Y(n_405)
);

INVx4_ASAP7_75t_L g406 ( 
.A(n_355),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_343),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_310),
.B(n_151),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_311),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_346),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_355),
.B(n_260),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_319),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_311),
.B(n_151),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_312),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_312),
.B(n_153),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_351),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_313),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_300),
.B(n_263),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_313),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_355),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_323),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_323),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_328),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_315),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_328),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_326),
.B(n_260),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_330),
.Y(n_427)
);

AND2x6_ASAP7_75t_L g428 ( 
.A(n_315),
.B(n_168),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_316),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_316),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_330),
.B(n_274),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_320),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_320),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_395),
.A2(n_302),
.B1(n_300),
.B2(n_361),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_384),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_370),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_406),
.B(n_324),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_383),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_384),
.Y(n_439)
);

INVx4_ASAP7_75t_L g440 ( 
.A(n_384),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_418),
.B(n_360),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_395),
.B(n_335),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_394),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_384),
.Y(n_444)
);

AOI22xp33_ASAP7_75t_L g445 ( 
.A1(n_369),
.A2(n_331),
.B1(n_295),
.B2(n_274),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_393),
.B(n_336),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g447 ( 
.A(n_399),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_401),
.Y(n_448)
);

OR2x6_ASAP7_75t_L g449 ( 
.A(n_396),
.B(n_364),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_384),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_394),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_402),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_383),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_402),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_370),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_372),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_407),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_403),
.B(n_340),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_372),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_382),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_382),
.Y(n_461)
);

AND2x6_ASAP7_75t_L g462 ( 
.A(n_374),
.B(n_295),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_402),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_409),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_406),
.B(n_341),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_409),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_426),
.B(n_326),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_406),
.B(n_344),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_386),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_386),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_406),
.B(n_349),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_409),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_384),
.Y(n_473)
);

NOR2x1p5_ASAP7_75t_L g474 ( 
.A(n_412),
.B(n_169),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_388),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_SL g476 ( 
.A1(n_418),
.A2(n_329),
.B1(n_314),
.B2(n_364),
.Y(n_476)
);

NAND2xp33_ASAP7_75t_SL g477 ( 
.A(n_380),
.B(n_222),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_388),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_398),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_380),
.B(n_350),
.Y(n_480)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_384),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_401),
.Y(n_482)
);

OAI22xp33_ASAP7_75t_L g483 ( 
.A1(n_380),
.A2(n_314),
.B1(n_329),
.B2(n_246),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_407),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_399),
.B(n_352),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_398),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_404),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_404),
.Y(n_488)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_387),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_414),
.Y(n_490)
);

INVx4_ASAP7_75t_L g491 ( 
.A(n_387),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_399),
.Y(n_492)
);

AO21x2_ASAP7_75t_L g493 ( 
.A1(n_400),
.A2(n_180),
.B(n_176),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_414),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_420),
.Y(n_495)
);

OAI22xp33_ASAP7_75t_L g496 ( 
.A1(n_408),
.A2(n_255),
.B1(n_254),
.B2(n_217),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_420),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_387),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_417),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_417),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_420),
.Y(n_501)
);

BUFx6f_ASAP7_75t_SL g502 ( 
.A(n_405),
.Y(n_502)
);

NAND3xp33_ASAP7_75t_L g503 ( 
.A(n_408),
.B(n_415),
.C(n_413),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_387),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_369),
.B(n_322),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_369),
.A2(n_405),
.B1(n_411),
.B2(n_431),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_413),
.B(n_325),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_426),
.B(n_332),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_424),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_424),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_410),
.Y(n_511)
);

AND3x2_ASAP7_75t_L g512 ( 
.A(n_374),
.B(n_150),
.C(n_184),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_426),
.B(n_332),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_415),
.B(n_153),
.Y(n_514)
);

INVxp33_ASAP7_75t_L g515 ( 
.A(n_383),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_374),
.Y(n_516)
);

OR2x2_ASAP7_75t_L g517 ( 
.A(n_405),
.B(n_347),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_424),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_397),
.B(n_423),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_419),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_424),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_423),
.B(n_425),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_419),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_405),
.B(n_157),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_424),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_405),
.B(n_167),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_419),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_431),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_387),
.Y(n_529)
);

INVx5_ASAP7_75t_L g530 ( 
.A(n_392),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_411),
.B(n_214),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_411),
.B(n_157),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_424),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_411),
.A2(n_183),
.B1(n_273),
.B2(n_334),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_425),
.B(n_367),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_431),
.B(n_368),
.Y(n_536)
);

INVxp33_ASAP7_75t_L g537 ( 
.A(n_385),
.Y(n_537)
);

NAND2xp33_ASAP7_75t_L g538 ( 
.A(n_392),
.B(n_183),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_427),
.B(n_368),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_431),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_431),
.B(n_158),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_410),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_424),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_419),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_424),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_430),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_430),
.Y(n_547)
);

BUFx10_ASAP7_75t_L g548 ( 
.A(n_427),
.Y(n_548)
);

INVx5_ASAP7_75t_L g549 ( 
.A(n_392),
.Y(n_549)
);

OAI22xp33_ASAP7_75t_L g550 ( 
.A1(n_396),
.A2(n_261),
.B1(n_235),
.B2(n_223),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_430),
.Y(n_551)
);

AND2x6_ASAP7_75t_L g552 ( 
.A(n_376),
.B(n_183),
.Y(n_552)
);

INVx4_ASAP7_75t_SL g553 ( 
.A(n_392),
.Y(n_553)
);

BUFx2_ASAP7_75t_L g554 ( 
.A(n_416),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_430),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_419),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_376),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_385),
.B(n_158),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_387),
.Y(n_559)
);

AND2x6_ASAP7_75t_L g560 ( 
.A(n_375),
.B(n_183),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_429),
.B(n_160),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_371),
.B(n_390),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_396),
.A2(n_173),
.B1(n_172),
.B2(n_293),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_387),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_371),
.B(n_218),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_430),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_SL g567 ( 
.A1(n_416),
.A2(n_222),
.B1(n_276),
.B2(n_277),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_430),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_400),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_430),
.B(n_160),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_421),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_373),
.Y(n_572)
);

NAND2x1p5_ASAP7_75t_L g573 ( 
.A(n_373),
.B(n_196),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_430),
.B(n_161),
.Y(n_574)
);

CKINVDCx14_ASAP7_75t_R g575 ( 
.A(n_433),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_387),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_516),
.B(n_448),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_516),
.B(n_333),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_503),
.B(n_371),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_540),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_478),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_478),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_506),
.B(n_183),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_557),
.B(n_273),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_486),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_540),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_442),
.A2(n_232),
.B1(n_230),
.B2(n_227),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_557),
.B(n_371),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_519),
.B(n_371),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_486),
.Y(n_590)
);

INVx8_ASAP7_75t_L g591 ( 
.A(n_449),
.Y(n_591)
);

INVxp67_ASAP7_75t_L g592 ( 
.A(n_480),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_495),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_528),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_505),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_528),
.B(n_273),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_487),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_487),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_495),
.B(n_334),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_507),
.B(n_161),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_447),
.B(n_273),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_536),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_501),
.B(n_273),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_492),
.B(n_163),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_572),
.A2(n_381),
.B(n_391),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_572),
.B(n_390),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_455),
.B(n_390),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_469),
.B(n_475),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_488),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_457),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_479),
.B(n_436),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_436),
.B(n_433),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_492),
.B(n_213),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_456),
.B(n_433),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_488),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_500),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_497),
.B(n_215),
.Y(n_617)
);

AO221x1_ASAP7_75t_L g618 ( 
.A1(n_496),
.A2(n_236),
.B1(n_245),
.B2(n_252),
.C(n_269),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_497),
.B(n_163),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_500),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_456),
.Y(n_621)
);

NOR3xp33_ASAP7_75t_L g622 ( 
.A(n_476),
.B(n_333),
.C(n_338),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_459),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_441),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_459),
.B(n_433),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_460),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_514),
.A2(n_221),
.B1(n_226),
.B2(n_234),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_517),
.B(n_338),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_460),
.B(n_433),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_434),
.B(n_164),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_461),
.Y(n_631)
);

O2A1O1Ixp33_ASAP7_75t_L g632 ( 
.A1(n_526),
.A2(n_381),
.B(n_339),
.C(n_345),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_461),
.B(n_433),
.Y(n_633)
);

NOR3xp33_ASAP7_75t_L g634 ( 
.A(n_558),
.B(n_342),
.C(n_353),
.Y(n_634)
);

NAND3xp33_ASAP7_75t_L g635 ( 
.A(n_445),
.B(n_239),
.C(n_240),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_470),
.B(n_490),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_470),
.B(n_433),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_490),
.Y(n_638)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_438),
.B(n_342),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_494),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_499),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_467),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_499),
.B(n_433),
.Y(n_643)
);

AO221x1_ASAP7_75t_L g644 ( 
.A1(n_483),
.A2(n_550),
.B1(n_569),
.B2(n_275),
.C(n_278),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_437),
.B(n_421),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_467),
.Y(n_646)
);

BUFx12f_ASAP7_75t_L g647 ( 
.A(n_449),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_443),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_435),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_530),
.B(n_284),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_443),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_451),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_530),
.B(n_549),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_530),
.B(n_238),
.Y(n_654)
);

BUFx5_ASAP7_75t_L g655 ( 
.A(n_569),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_508),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_451),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_530),
.B(n_241),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_508),
.B(n_339),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_452),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_482),
.B(n_164),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_513),
.Y(n_662)
);

OAI221xp5_ASAP7_75t_L g663 ( 
.A1(n_477),
.A2(n_362),
.B1(n_366),
.B2(n_365),
.C(n_363),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_517),
.B(n_353),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_513),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_522),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_485),
.B(n_166),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_520),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_452),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_482),
.B(n_446),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_454),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_462),
.A2(n_242),
.B1(n_247),
.B2(n_248),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_465),
.B(n_421),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_523),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_454),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_463),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_527),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_544),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_530),
.B(n_251),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_468),
.B(n_421),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_458),
.B(n_166),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_502),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_556),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_549),
.B(n_257),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_512),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_548),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_502),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_471),
.B(n_421),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_463),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_561),
.B(n_422),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_464),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_502),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_531),
.B(n_422),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_462),
.B(n_422),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_462),
.B(n_422),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_549),
.B(n_266),
.Y(n_696)
);

INVxp67_ASAP7_75t_SL g697 ( 
.A(n_435),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_548),
.Y(n_698)
);

NOR2x1p5_ASAP7_75t_L g699 ( 
.A(n_449),
.B(n_276),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_464),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_462),
.B(n_422),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_534),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_462),
.B(n_375),
.Y(n_703)
);

INVxp67_ASAP7_75t_SL g704 ( 
.A(n_435),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_549),
.B(n_268),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_524),
.A2(n_170),
.B1(n_171),
.B2(n_293),
.Y(n_706)
);

NOR3xp33_ASAP7_75t_L g707 ( 
.A(n_453),
.B(n_356),
.C(n_366),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_548),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_477),
.A2(n_373),
.B1(n_281),
.B2(n_286),
.Y(n_709)
);

NOR2xp67_ASAP7_75t_L g710 ( 
.A(n_563),
.B(n_535),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_575),
.B(n_377),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_532),
.A2(n_173),
.B1(n_271),
.B2(n_290),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_457),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_474),
.B(n_567),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_511),
.B(n_542),
.Y(n_715)
);

NAND3xp33_ASAP7_75t_L g716 ( 
.A(n_541),
.B(n_174),
.C(n_178),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_466),
.Y(n_717)
);

INVxp67_ASAP7_75t_SL g718 ( 
.A(n_435),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_573),
.B(n_377),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_573),
.B(n_378),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_537),
.B(n_271),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_571),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_484),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_466),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_549),
.B(n_283),
.Y(n_725)
);

AND2x6_ASAP7_75t_L g726 ( 
.A(n_509),
.B(n_510),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_472),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_472),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_565),
.B(n_283),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_562),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_450),
.B(n_379),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_435),
.Y(n_732)
);

O2A1O1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_570),
.A2(n_345),
.B(n_359),
.C(n_358),
.Y(n_733)
);

BUFx5_ASAP7_75t_L g734 ( 
.A(n_560),
.Y(n_734)
);

OAI22xp33_ASAP7_75t_L g735 ( 
.A1(n_624),
.A2(n_449),
.B1(n_515),
.B2(n_542),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_577),
.B(n_511),
.Y(n_736)
);

BUFx4f_ASAP7_75t_SL g737 ( 
.A(n_723),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_592),
.B(n_554),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_594),
.Y(n_739)
);

OR2x4_ASAP7_75t_L g740 ( 
.A(n_630),
.B(n_539),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_621),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_580),
.Y(n_742)
);

INVxp67_ASAP7_75t_L g743 ( 
.A(n_639),
.Y(n_743)
);

NOR2x1_ASAP7_75t_R g744 ( 
.A(n_647),
.B(n_554),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_666),
.B(n_498),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_580),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_610),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_638),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_638),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_642),
.B(n_553),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_600),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_661),
.B(n_484),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_715),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_721),
.B(n_574),
.Y(n_754)
);

INVx3_ASAP7_75t_L g755 ( 
.A(n_593),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_628),
.B(n_356),
.Y(n_756)
);

O2A1O1Ixp33_ASAP7_75t_L g757 ( 
.A1(n_602),
.A2(n_538),
.B(n_568),
.C(n_566),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_641),
.B(n_504),
.Y(n_758)
);

NOR2x1p5_ASAP7_75t_L g759 ( 
.A(n_708),
.B(n_698),
.Y(n_759)
);

OR2x4_ASAP7_75t_L g760 ( 
.A(n_630),
.B(n_358),
.Y(n_760)
);

NOR2xp67_ASAP7_75t_L g761 ( 
.A(n_686),
.B(n_359),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_667),
.B(n_504),
.Y(n_762)
);

A2O1A1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_600),
.A2(n_521),
.B(n_568),
.C(n_566),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_667),
.B(n_504),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_713),
.Y(n_765)
);

INVxp67_ASAP7_75t_L g766 ( 
.A(n_721),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_578),
.B(n_623),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_583),
.A2(n_493),
.B1(n_552),
.B2(n_510),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_626),
.B(n_529),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_641),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_649),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_581),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_581),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_599),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_599),
.B(n_553),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_659),
.B(n_553),
.Y(n_776)
);

INVx2_ASAP7_75t_SL g777 ( 
.A(n_659),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_670),
.B(n_708),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_670),
.B(n_595),
.Y(n_779)
);

NAND2x1p5_ASAP7_75t_L g780 ( 
.A(n_682),
.B(n_687),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_649),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_655),
.B(n_529),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_685),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_582),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_593),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_664),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_585),
.Y(n_787)
);

OR2x6_ASAP7_75t_L g788 ( 
.A(n_591),
.B(n_362),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_591),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_649),
.Y(n_790)
);

BUFx4f_ASAP7_75t_L g791 ( 
.A(n_591),
.Y(n_791)
);

OR2x6_ASAP7_75t_L g792 ( 
.A(n_682),
.B(n_365),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_646),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_655),
.B(n_529),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_649),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_655),
.B(n_636),
.Y(n_796)
);

INVx2_ASAP7_75t_SL g797 ( 
.A(n_656),
.Y(n_797)
);

NOR3xp33_ASAP7_75t_SL g798 ( 
.A(n_663),
.B(n_281),
.C(n_286),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_710),
.B(n_553),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_655),
.B(n_564),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_662),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_665),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_585),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_714),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_655),
.B(n_564),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_687),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_655),
.B(n_730),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_692),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_590),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_597),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_631),
.B(n_564),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_640),
.B(n_576),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_611),
.B(n_576),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_729),
.A2(n_552),
.B1(n_493),
.B2(n_509),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_597),
.Y(n_815)
);

A2O1A1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_681),
.A2(n_525),
.B(n_555),
.C(n_551),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_598),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_692),
.Y(n_818)
);

CKINVDCx20_ASAP7_75t_R g819 ( 
.A(n_681),
.Y(n_819)
);

OAI21xp5_ASAP7_75t_L g820 ( 
.A1(n_606),
.A2(n_576),
.B(n_546),
.Y(n_820)
);

BUFx4f_ASAP7_75t_L g821 ( 
.A(n_586),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_604),
.B(n_288),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_729),
.B(n_440),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_604),
.B(n_288),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_716),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_608),
.B(n_619),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_619),
.B(n_440),
.Y(n_827)
);

INVx4_ASAP7_75t_L g828 ( 
.A(n_726),
.Y(n_828)
);

OR2x6_ASAP7_75t_L g829 ( 
.A(n_699),
.B(n_518),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_609),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_587),
.B(n_289),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_627),
.B(n_289),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_613),
.B(n_290),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_609),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_589),
.B(n_473),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_615),
.Y(n_836)
);

OAI221xp5_ASAP7_75t_L g837 ( 
.A1(n_622),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.C(n_207),
.Y(n_837)
);

INVxp67_ASAP7_75t_L g838 ( 
.A(n_707),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_616),
.B(n_439),
.Y(n_839)
);

BUFx3_ASAP7_75t_L g840 ( 
.A(n_722),
.Y(n_840)
);

NOR2x1p5_ASAP7_75t_L g841 ( 
.A(n_635),
.B(n_177),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_616),
.B(n_439),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_620),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_620),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_668),
.B(n_439),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_726),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_583),
.A2(n_493),
.B1(n_552),
.B2(n_555),
.Y(n_847)
);

INVxp67_ASAP7_75t_L g848 ( 
.A(n_613),
.Y(n_848)
);

OR2x6_ASAP7_75t_L g849 ( 
.A(n_617),
.B(n_518),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_726),
.Y(n_850)
);

BUFx12f_ASAP7_75t_L g851 ( 
.A(n_726),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_644),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_617),
.B(n_473),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_674),
.B(n_444),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_677),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_709),
.A2(n_552),
.B1(n_521),
.B2(n_545),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_579),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_709),
.A2(n_552),
.B1(n_546),
.B2(n_543),
.Y(n_858)
);

NAND2x1_ASAP7_75t_L g859 ( 
.A(n_726),
.B(n_732),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_732),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_678),
.B(n_444),
.Y(n_861)
);

BUFx10_ASAP7_75t_L g862 ( 
.A(n_683),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_588),
.B(n_444),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_648),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_648),
.B(n_444),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_706),
.B(n_292),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_711),
.Y(n_867)
);

OR2x2_ASAP7_75t_L g868 ( 
.A(n_712),
.B(n_233),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_719),
.A2(n_491),
.B(n_473),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_634),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_651),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_651),
.B(n_652),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_652),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_672),
.B(n_292),
.Y(n_874)
);

INVx4_ASAP7_75t_L g875 ( 
.A(n_657),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_657),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_660),
.B(n_669),
.Y(n_877)
);

NAND2x1p5_ASAP7_75t_L g878 ( 
.A(n_653),
.B(n_481),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_703),
.B(n_525),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_618),
.A2(n_552),
.B1(n_533),
.B2(n_547),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_660),
.B(n_559),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_694),
.Y(n_882)
);

INVxp67_ASAP7_75t_L g883 ( 
.A(n_702),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_669),
.B(n_559),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_671),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_675),
.B(n_559),
.Y(n_886)
);

AOI21x1_ASAP7_75t_L g887 ( 
.A1(n_605),
.A2(n_545),
.B(n_533),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_675),
.Y(n_888)
);

INVx5_ASAP7_75t_L g889 ( 
.A(n_676),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_697),
.B(n_481),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_676),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_704),
.B(n_489),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_725),
.A2(n_551),
.B1(n_547),
.B2(n_543),
.Y(n_893)
);

A2O1A1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_693),
.A2(n_538),
.B(n_432),
.C(n_429),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_689),
.Y(n_895)
);

BUFx8_ASAP7_75t_SL g896 ( 
.A(n_607),
.Y(n_896)
);

INVxp67_ASAP7_75t_SL g897 ( 
.A(n_718),
.Y(n_897)
);

INVx5_ASAP7_75t_L g898 ( 
.A(n_689),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_724),
.A2(n_373),
.B1(n_428),
.B2(n_560),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_691),
.B(n_559),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_691),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_700),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_695),
.Y(n_903)
);

NAND3xp33_ASAP7_75t_SL g904 ( 
.A(n_733),
.B(n_237),
.C(n_249),
.Y(n_904)
);

NOR2xp67_ASAP7_75t_L g905 ( 
.A(n_727),
.B(n_73),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_766),
.B(n_701),
.Y(n_906)
);

NOR3xp33_ASAP7_75t_SL g907 ( 
.A(n_735),
.B(n_264),
.C(n_253),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_753),
.Y(n_908)
);

NOR3xp33_ASAP7_75t_SL g909 ( 
.A(n_752),
.B(n_265),
.C(n_267),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_779),
.B(n_720),
.Y(n_910)
);

O2A1O1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_754),
.A2(n_584),
.B(n_596),
.C(n_601),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_826),
.B(n_700),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_741),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_857),
.B(n_717),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_796),
.A2(n_673),
.B(n_688),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_767),
.B(n_717),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_751),
.A2(n_680),
.B(n_645),
.C(n_632),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_786),
.B(n_734),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_883),
.A2(n_643),
.B(n_612),
.C(n_614),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_749),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_SL g921 ( 
.A1(n_819),
.A2(n_297),
.B1(n_270),
.B2(n_250),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_796),
.A2(n_653),
.B(n_690),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_756),
.B(n_867),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_736),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_743),
.B(n_725),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_867),
.B(n_728),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_867),
.B(n_728),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_777),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_822),
.A2(n_584),
.B(n_596),
.C(n_603),
.Y(n_929)
);

NOR2x1_ASAP7_75t_R g930 ( 
.A(n_747),
.B(n_601),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_L g931 ( 
.A1(n_852),
.A2(n_684),
.B1(n_654),
.B2(n_658),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_739),
.B(n_625),
.Y(n_932)
);

CKINVDCx20_ASAP7_75t_R g933 ( 
.A(n_737),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_748),
.Y(n_934)
);

NAND2x1p5_ASAP7_75t_L g935 ( 
.A(n_828),
.B(n_603),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_821),
.B(n_734),
.Y(n_936)
);

INVx4_ASAP7_75t_L g937 ( 
.A(n_775),
.Y(n_937)
);

O2A1O1Ixp5_ASAP7_75t_SL g938 ( 
.A1(n_778),
.A2(n_684),
.B(n_696),
.C(n_705),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_823),
.A2(n_491),
.B(n_489),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_774),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_807),
.A2(n_629),
.B1(n_637),
.B2(n_633),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_821),
.B(n_734),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_770),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_745),
.B(n_731),
.Y(n_944)
);

NAND3xp33_ASAP7_75t_L g945 ( 
.A(n_738),
.B(n_824),
.C(n_838),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_807),
.A2(n_705),
.B(n_696),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_783),
.Y(n_947)
);

BUFx2_ASAP7_75t_R g948 ( 
.A(n_789),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_890),
.A2(n_679),
.B(n_658),
.Y(n_949)
);

O2A1O1Ixp33_ASAP7_75t_SL g950 ( 
.A1(n_799),
.A2(n_679),
.B(n_654),
.C(n_650),
.Y(n_950)
);

OR2x6_ASAP7_75t_L g951 ( 
.A(n_788),
.B(n_650),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_804),
.Y(n_952)
);

O2A1O1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_837),
.A2(n_429),
.B(n_432),
.C(n_389),
.Y(n_953)
);

AO32x2_ASAP7_75t_L g954 ( 
.A1(n_875),
.A2(n_1),
.A3(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_954)
);

O2A1O1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_866),
.A2(n_432),
.B(n_389),
.C(n_9),
.Y(n_955)
);

AOI22xp33_ASAP7_75t_L g956 ( 
.A1(n_831),
.A2(n_734),
.B1(n_560),
.B2(n_428),
.Y(n_956)
);

OAI21x1_ASAP7_75t_L g957 ( 
.A1(n_887),
.A2(n_389),
.B(n_734),
.Y(n_957)
);

INVx8_ASAP7_75t_L g958 ( 
.A(n_851),
.Y(n_958)
);

INVx4_ASAP7_75t_L g959 ( 
.A(n_775),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_772),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_891),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_776),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_848),
.B(n_734),
.Y(n_963)
);

BUFx2_ASAP7_75t_L g964 ( 
.A(n_792),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_892),
.A2(n_391),
.B(n_392),
.Y(n_965)
);

BUFx2_ASAP7_75t_L g966 ( 
.A(n_792),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_776),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_771),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_760),
.A2(n_740),
.B1(n_856),
.B2(n_858),
.Y(n_969)
);

NAND2xp33_ASAP7_75t_L g970 ( 
.A(n_806),
.B(n_560),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_820),
.A2(n_560),
.B(n_428),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_870),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_SL g973 ( 
.A(n_765),
.B(n_560),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_841),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_L g975 ( 
.A1(n_760),
.A2(n_391),
.B1(n_16),
.B2(n_17),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_L g976 ( 
.A1(n_740),
.A2(n_391),
.B1(n_16),
.B2(n_19),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_793),
.B(n_392),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_797),
.B(n_392),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_750),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_840),
.B(n_391),
.Y(n_980)
);

OA22x2_ASAP7_75t_L g981 ( 
.A1(n_801),
.A2(n_10),
.B1(n_20),
.B2(n_22),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_771),
.Y(n_982)
);

O2A1O1Ixp5_ASAP7_75t_L g983 ( 
.A1(n_827),
.A2(n_64),
.B(n_144),
.C(n_143),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_802),
.B(n_392),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_782),
.A2(n_391),
.B(n_53),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_765),
.B(n_868),
.Y(n_986)
);

INVx4_ASAP7_75t_L g987 ( 
.A(n_806),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_750),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_792),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_R g990 ( 
.A(n_791),
.B(n_138),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_896),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_897),
.B(n_25),
.Y(n_992)
);

OAI321xp33_ASAP7_75t_L g993 ( 
.A1(n_833),
.A2(n_25),
.A3(n_30),
.B1(n_34),
.B2(n_35),
.C(n_36),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_771),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_825),
.B(n_30),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_745),
.B(n_428),
.Y(n_996)
);

BUFx2_ASAP7_75t_L g997 ( 
.A(n_788),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_794),
.A2(n_800),
.B(n_805),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_781),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_SL g1000 ( 
.A(n_791),
.B(n_428),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_829),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_862),
.B(n_806),
.Y(n_1002)
);

AOI221xp5_ASAP7_75t_L g1003 ( 
.A1(n_832),
.A2(n_34),
.B1(n_37),
.B2(n_39),
.C(n_40),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_855),
.B(n_39),
.Y(n_1004)
);

CKINVDCx16_ASAP7_75t_R g1005 ( 
.A(n_788),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_874),
.A2(n_428),
.B1(n_42),
.B2(n_46),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_755),
.B(n_41),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_805),
.A2(n_77),
.B(n_79),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_835),
.A2(n_108),
.B(n_428),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_784),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_862),
.B(n_42),
.Y(n_1011)
);

AOI21x1_ASAP7_75t_L g1012 ( 
.A1(n_762),
.A2(n_764),
.B(n_863),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_798),
.A2(n_47),
.B(n_48),
.C(n_428),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_755),
.B(n_428),
.Y(n_1014)
);

OR2x6_ASAP7_75t_L g1015 ( 
.A(n_829),
.B(n_428),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_785),
.B(n_813),
.Y(n_1016)
);

OAI21xp33_ASAP7_75t_L g1017 ( 
.A1(n_808),
.A2(n_853),
.B(n_761),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_814),
.A2(n_757),
.B(n_813),
.C(n_879),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_882),
.B(n_903),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_882),
.B(n_903),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_818),
.Y(n_1021)
);

OA21x2_ASAP7_75t_L g1022 ( 
.A1(n_820),
.A2(n_816),
.B(n_763),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_781),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_818),
.B(n_785),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_882),
.B(n_903),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_873),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_768),
.A2(n_847),
.B1(n_828),
.B2(n_746),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_742),
.B(n_746),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_742),
.B(n_875),
.Y(n_1029)
);

NAND3xp33_ASAP7_75t_L g1030 ( 
.A(n_849),
.B(n_880),
.C(n_879),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_869),
.A2(n_863),
.B(n_842),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_889),
.A2(n_898),
.B1(n_899),
.B2(n_846),
.Y(n_1032)
);

AOI21x1_ASAP7_75t_L g1033 ( 
.A1(n_946),
.A2(n_845),
.B(n_854),
.Y(n_1033)
);

AOI221x1_ASAP7_75t_L g1034 ( 
.A1(n_976),
.A2(n_975),
.B1(n_969),
.B2(n_1027),
.C(n_1031),
.Y(n_1034)
);

NAND3xp33_ASAP7_75t_L g1035 ( 
.A(n_995),
.B(n_849),
.C(n_894),
.Y(n_1035)
);

AO31x2_ASAP7_75t_L g1036 ( 
.A1(n_1018),
.A2(n_854),
.A3(n_861),
.B(n_845),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_908),
.Y(n_1037)
);

NOR2xp67_ASAP7_75t_SL g1038 ( 
.A(n_993),
.B(n_846),
.Y(n_1038)
);

OAI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_922),
.A2(n_758),
.B(n_893),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_933),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_924),
.B(n_759),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_939),
.A2(n_877),
.B(n_872),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_1032),
.A2(n_898),
.B(n_889),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_986),
.B(n_744),
.Y(n_1044)
);

AO31x2_ASAP7_75t_L g1045 ( 
.A1(n_1027),
.A2(n_861),
.A3(n_812),
.B(n_811),
.Y(n_1045)
);

OA22x2_ASAP7_75t_L g1046 ( 
.A1(n_975),
.A2(n_976),
.B1(n_921),
.B2(n_952),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_960),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_1032),
.A2(n_839),
.B(n_842),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_923),
.B(n_846),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_910),
.B(n_844),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_912),
.B(n_830),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_945),
.B(n_850),
.Y(n_1052)
);

NOR2xp67_ASAP7_75t_SL g1053 ( 
.A(n_1005),
.B(n_850),
.Y(n_1053)
);

AOI21x1_ASAP7_75t_L g1054 ( 
.A1(n_1012),
.A2(n_812),
.B(n_811),
.Y(n_1054)
);

AO31x2_ASAP7_75t_L g1055 ( 
.A1(n_917),
.A2(n_941),
.A3(n_969),
.B(n_919),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_912),
.B(n_834),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_916),
.B(n_810),
.Y(n_1057)
);

NAND2x1p5_ASAP7_75t_L g1058 ( 
.A(n_987),
.B(n_795),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_947),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_938),
.A2(n_900),
.B(n_886),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_916),
.B(n_815),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_1019),
.B(n_809),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_937),
.B(n_850),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1010),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_962),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_1019),
.B(n_787),
.Y(n_1066)
);

AOI21x1_ASAP7_75t_L g1067 ( 
.A1(n_941),
.A2(n_905),
.B(n_769),
.Y(n_1067)
);

AO32x2_ASAP7_75t_L g1068 ( 
.A1(n_974),
.A2(n_904),
.A3(n_849),
.B1(n_836),
.B2(n_817),
.Y(n_1068)
);

INVxp67_ASAP7_75t_SL g1069 ( 
.A(n_1029),
.Y(n_1069)
);

AOI211x1_ASAP7_75t_L g1070 ( 
.A1(n_1004),
.A2(n_803),
.B(n_895),
.C(n_885),
.Y(n_1070)
);

OAI21x1_ASAP7_75t_L g1071 ( 
.A1(n_965),
.A2(n_886),
.B(n_884),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_944),
.A2(n_881),
.B(n_865),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_1016),
.A2(n_985),
.B(n_971),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_950),
.A2(n_859),
.B(n_781),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_911),
.A2(n_790),
.B(n_795),
.Y(n_1075)
);

AOI21x1_ASAP7_75t_L g1076 ( 
.A1(n_1022),
.A2(n_902),
.B(n_876),
.Y(n_1076)
);

AO21x1_ASAP7_75t_L g1077 ( 
.A1(n_955),
.A2(n_871),
.B(n_864),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_1030),
.A2(n_795),
.B(n_790),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_971),
.A2(n_773),
.B(n_843),
.Y(n_1079)
);

NOR2x1_ASAP7_75t_SL g1080 ( 
.A(n_936),
.B(n_790),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_935),
.A2(n_888),
.B(n_901),
.Y(n_1081)
);

OA21x2_ASAP7_75t_L g1082 ( 
.A1(n_983),
.A2(n_878),
.B(n_780),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_SL g1083 ( 
.A(n_948),
.B(n_860),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_925),
.A2(n_860),
.B(n_929),
.C(n_907),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1020),
.B(n_1025),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_913),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_1011),
.A2(n_972),
.B(n_1013),
.C(n_1003),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_962),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_964),
.B(n_966),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1020),
.A2(n_1025),
.B(n_1017),
.Y(n_1090)
);

OA22x2_ASAP7_75t_L g1091 ( 
.A1(n_989),
.A2(n_1001),
.B1(n_997),
.B2(n_940),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_932),
.A2(n_906),
.B(n_942),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_928),
.B(n_930),
.Y(n_1093)
);

INVx2_ASAP7_75t_SL g1094 ( 
.A(n_1021),
.Y(n_1094)
);

INVx4_ASAP7_75t_L g1095 ( 
.A(n_968),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_968),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_920),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_926),
.B(n_927),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_931),
.A2(n_909),
.B(n_992),
.C(n_1007),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_963),
.A2(n_1028),
.B(n_918),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_996),
.A2(n_1028),
.B(n_914),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_914),
.A2(n_1009),
.B(n_996),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_934),
.Y(n_1103)
);

AND3x4_ASAP7_75t_L g1104 ( 
.A(n_991),
.B(n_958),
.C(n_1026),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_943),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_979),
.B(n_988),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_979),
.B(n_988),
.Y(n_1107)
);

AOI21xp33_ASAP7_75t_L g1108 ( 
.A1(n_981),
.A2(n_953),
.B(n_1006),
.Y(n_1108)
);

NAND3xp33_ASAP7_75t_L g1109 ( 
.A(n_1008),
.B(n_951),
.C(n_1002),
.Y(n_1109)
);

INVx4_ASAP7_75t_L g1110 ( 
.A(n_968),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_961),
.A2(n_1024),
.B(n_980),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_967),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_958),
.Y(n_1113)
);

BUFx4_ASAP7_75t_SL g1114 ( 
.A(n_951),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_967),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_970),
.A2(n_1014),
.B(n_973),
.Y(n_1116)
);

INVxp67_ASAP7_75t_L g1117 ( 
.A(n_981),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_958),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_937),
.B(n_959),
.Y(n_1119)
);

AO21x1_ASAP7_75t_L g1120 ( 
.A1(n_954),
.A2(n_977),
.B(n_978),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_951),
.A2(n_1015),
.B1(n_959),
.B2(n_954),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_987),
.B(n_1015),
.Y(n_1122)
);

NOR2xp67_ASAP7_75t_SL g1123 ( 
.A(n_982),
.B(n_994),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1015),
.A2(n_954),
.B1(n_956),
.B2(n_982),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_982),
.B(n_994),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_994),
.Y(n_1126)
);

NAND3xp33_ASAP7_75t_L g1127 ( 
.A(n_984),
.B(n_1000),
.C(n_999),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_999),
.A2(n_1023),
.B(n_990),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_999),
.B(n_1023),
.Y(n_1129)
);

AOI221x1_ASAP7_75t_L g1130 ( 
.A1(n_976),
.A2(n_975),
.B1(n_969),
.B2(n_1027),
.C(n_1031),
.Y(n_1130)
);

A2O1A1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_910),
.A2(n_754),
.B(n_751),
.C(n_779),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_960),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_910),
.B(n_912),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_SL g1134 ( 
.A1(n_963),
.A2(n_799),
.B(n_969),
.C(n_942),
.Y(n_1134)
);

O2A1O1Ixp33_ASAP7_75t_SL g1135 ( 
.A1(n_963),
.A2(n_799),
.B(n_969),
.C(n_942),
.Y(n_1135)
);

OAI21xp5_ASAP7_75t_SL g1136 ( 
.A1(n_995),
.A2(n_537),
.B(n_751),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_924),
.B(n_766),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_915),
.A2(n_796),
.B(n_823),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_910),
.B(n_912),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_R g1140 ( 
.A(n_933),
.B(n_407),
.Y(n_1140)
);

AOI221x1_ASAP7_75t_L g1141 ( 
.A1(n_976),
.A2(n_975),
.B1(n_969),
.B2(n_1027),
.C(n_1031),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_986),
.B(n_766),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_957),
.A2(n_887),
.B(n_1031),
.Y(n_1143)
);

OAI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1018),
.A2(n_915),
.B(n_998),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_910),
.B(n_912),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_957),
.A2(n_887),
.B(n_1031),
.Y(n_1146)
);

AOI21x1_ASAP7_75t_L g1147 ( 
.A1(n_946),
.A2(n_949),
.B(n_1012),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_910),
.B(n_912),
.Y(n_1148)
);

AO21x2_ASAP7_75t_L g1149 ( 
.A1(n_1012),
.A2(n_1031),
.B(n_1018),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_910),
.B(n_912),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1018),
.A2(n_915),
.B(n_998),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_910),
.B(n_912),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_910),
.B(n_912),
.Y(n_1153)
);

NOR2xp67_ASAP7_75t_L g1154 ( 
.A(n_945),
.B(n_743),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_957),
.A2(n_887),
.B(n_1031),
.Y(n_1155)
);

OR2x2_ASAP7_75t_L g1156 ( 
.A(n_924),
.B(n_766),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_957),
.A2(n_887),
.B(n_1031),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_910),
.B(n_912),
.Y(n_1158)
);

AO31x2_ASAP7_75t_L g1159 ( 
.A1(n_1018),
.A2(n_1027),
.A3(n_1031),
.B(n_816),
.Y(n_1159)
);

AO21x2_ASAP7_75t_L g1160 ( 
.A1(n_1144),
.A2(n_1151),
.B(n_1147),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_1059),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1143),
.A2(n_1155),
.B(n_1146),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_SL g1163 ( 
.A1(n_1046),
.A2(n_1142),
.B1(n_1121),
.B2(n_1144),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_1046),
.A2(n_1038),
.B1(n_1108),
.B2(n_1117),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1157),
.A2(n_1071),
.B(n_1042),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1131),
.A2(n_1099),
.B(n_1087),
.Y(n_1166)
);

INVx3_ASAP7_75t_SL g1167 ( 
.A(n_1040),
.Y(n_1167)
);

OR2x2_ASAP7_75t_L g1168 ( 
.A(n_1085),
.B(n_1156),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1076),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1137),
.B(n_1089),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1047),
.Y(n_1171)
);

NAND2x1p5_ASAP7_75t_L g1172 ( 
.A(n_1053),
.B(n_1123),
.Y(n_1172)
);

NAND3xp33_ASAP7_75t_L g1173 ( 
.A(n_1136),
.B(n_1154),
.C(n_1084),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1133),
.A2(n_1150),
.B1(n_1158),
.B2(n_1153),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1133),
.A2(n_1150),
.B1(n_1158),
.B2(n_1153),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_1096),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1139),
.A2(n_1152),
.B1(n_1145),
.B2(n_1148),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1139),
.B(n_1145),
.Y(n_1178)
);

OAI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1034),
.A2(n_1130),
.B1(n_1141),
.B2(n_1152),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1085),
.B(n_1041),
.Y(n_1180)
);

AOI21x1_ASAP7_75t_SL g1181 ( 
.A1(n_1148),
.A2(n_1050),
.B(n_1051),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1050),
.B(n_1069),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_1037),
.Y(n_1183)
);

BUFx12f_ASAP7_75t_L g1184 ( 
.A(n_1118),
.Y(n_1184)
);

OA21x2_ASAP7_75t_L g1185 ( 
.A1(n_1151),
.A2(n_1060),
.B(n_1138),
.Y(n_1185)
);

AO21x1_ASAP7_75t_L g1186 ( 
.A1(n_1052),
.A2(n_1121),
.B(n_1108),
.Y(n_1186)
);

OR2x6_ASAP7_75t_L g1187 ( 
.A(n_1090),
.B(n_1078),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1064),
.Y(n_1188)
);

O2A1O1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_1134),
.A2(n_1135),
.B(n_1044),
.C(n_1093),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_1128),
.Y(n_1190)
);

OA21x2_ASAP7_75t_L g1191 ( 
.A1(n_1060),
.A2(n_1073),
.B(n_1039),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1033),
.A2(n_1074),
.B(n_1102),
.Y(n_1192)
);

INVxp67_ASAP7_75t_L g1193 ( 
.A(n_1094),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1122),
.B(n_1065),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_SL g1195 ( 
.A(n_1083),
.B(n_1104),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1098),
.B(n_1062),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1035),
.A2(n_1109),
.B1(n_1091),
.B2(n_1105),
.Y(n_1197)
);

OA21x2_ASAP7_75t_L g1198 ( 
.A1(n_1039),
.A2(n_1067),
.B(n_1048),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1092),
.A2(n_1100),
.B(n_1075),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1079),
.A2(n_1054),
.B(n_1101),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1062),
.B(n_1066),
.Y(n_1201)
);

OA21x2_ASAP7_75t_L g1202 ( 
.A1(n_1077),
.A2(n_1120),
.B(n_1072),
.Y(n_1202)
);

BUFx12f_ASAP7_75t_L g1203 ( 
.A(n_1113),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_1106),
.B(n_1107),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_1122),
.B(n_1065),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1066),
.B(n_1056),
.Y(n_1206)
);

OA21x2_ASAP7_75t_L g1207 ( 
.A1(n_1043),
.A2(n_1051),
.B(n_1056),
.Y(n_1207)
);

NAND2x1p5_ASAP7_75t_L g1208 ( 
.A(n_1049),
.B(n_1088),
.Y(n_1208)
);

AOI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1091),
.A2(n_1083),
.B1(n_1119),
.B2(n_1127),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1086),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1116),
.A2(n_1111),
.B(n_1061),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1057),
.A2(n_1061),
.B(n_1081),
.Y(n_1212)
);

NAND2x1p5_ASAP7_75t_L g1213 ( 
.A(n_1088),
.B(n_1063),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1063),
.B(n_1115),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1082),
.A2(n_1124),
.B(n_1057),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_1112),
.B(n_1106),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_1140),
.Y(n_1217)
);

INVx3_ASAP7_75t_L g1218 ( 
.A(n_1095),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1082),
.A2(n_1124),
.B(n_1107),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1097),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_SL g1221 ( 
.A1(n_1080),
.A2(n_1132),
.B(n_1125),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1103),
.Y(n_1222)
);

CKINVDCx16_ASAP7_75t_R g1223 ( 
.A(n_1110),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1068),
.A2(n_1149),
.A3(n_1159),
.B(n_1055),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_1114),
.Y(n_1225)
);

O2A1O1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1129),
.A2(n_1126),
.B(n_1125),
.C(n_1058),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1070),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1058),
.A2(n_1036),
.B(n_1159),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1036),
.A2(n_1068),
.B(n_1045),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1159),
.A2(n_1045),
.B(n_1068),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1055),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1055),
.A2(n_1131),
.B(n_1136),
.C(n_751),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1045),
.A2(n_1146),
.B(n_1143),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_1096),
.Y(n_1234)
);

BUFx6f_ASAP7_75t_L g1235 ( 
.A(n_1096),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1046),
.A2(n_754),
.B1(n_819),
.B2(n_1003),
.Y(n_1236)
);

NAND2x1p5_ASAP7_75t_L g1237 ( 
.A(n_1053),
.B(n_1123),
.Y(n_1237)
);

OR2x6_ASAP7_75t_L g1238 ( 
.A(n_1090),
.B(n_1078),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1137),
.B(n_766),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1046),
.A2(n_754),
.B1(n_819),
.B2(n_1003),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1047),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1137),
.B(n_766),
.Y(n_1242)
);

BUFx3_ASAP7_75t_L g1243 ( 
.A(n_1059),
.Y(n_1243)
);

INVx6_ASAP7_75t_L g1244 ( 
.A(n_1059),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_SL g1245 ( 
.A1(n_1080),
.A2(n_1077),
.B(n_1043),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1137),
.B(n_766),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1142),
.B(n_766),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1059),
.Y(n_1248)
);

AO31x2_ASAP7_75t_L g1249 ( 
.A1(n_1034),
.A2(n_1141),
.A3(n_1130),
.B(n_1120),
.Y(n_1249)
);

NAND2x1p5_ASAP7_75t_L g1250 ( 
.A(n_1053),
.B(n_1123),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1047),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1143),
.A2(n_1146),
.B(n_1155),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1142),
.B(n_766),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1131),
.A2(n_754),
.B(n_1087),
.C(n_1144),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1046),
.A2(n_754),
.B1(n_819),
.B2(n_1003),
.Y(n_1255)
);

AO21x2_ASAP7_75t_L g1256 ( 
.A1(n_1144),
.A2(n_1151),
.B(n_1147),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1143),
.A2(n_1146),
.B(n_1155),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1047),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1143),
.A2(n_1146),
.B(n_1155),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_1122),
.B(n_1085),
.Y(n_1260)
);

OR2x2_ASAP7_75t_L g1261 ( 
.A(n_1085),
.B(n_1156),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_R g1262 ( 
.A(n_1083),
.B(n_933),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1131),
.B(n_1133),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1047),
.Y(n_1264)
);

NAND3xp33_ASAP7_75t_L g1265 ( 
.A(n_1131),
.B(n_442),
.C(n_754),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1142),
.A2(n_819),
.B1(n_482),
.B2(n_1131),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1144),
.A2(n_1151),
.B(n_1138),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1122),
.B(n_1085),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1059),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1047),
.Y(n_1270)
);

AO21x1_ASAP7_75t_L g1271 ( 
.A1(n_1087),
.A2(n_976),
.B(n_975),
.Y(n_1271)
);

AO21x2_ASAP7_75t_L g1272 ( 
.A1(n_1144),
.A2(n_1151),
.B(n_1147),
.Y(n_1272)
);

A2O1A1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1131),
.A2(n_754),
.B(n_1087),
.C(n_1144),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1144),
.A2(n_1151),
.B(n_1138),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1143),
.A2(n_1146),
.B(n_1155),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1144),
.A2(n_1151),
.B(n_1138),
.Y(n_1276)
);

BUFx12f_ASAP7_75t_L g1277 ( 
.A(n_1040),
.Y(n_1277)
);

INVx8_ASAP7_75t_L g1278 ( 
.A(n_1234),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_SL g1279 ( 
.A1(n_1254),
.A2(n_1273),
.B(n_1265),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1236),
.A2(n_1255),
.B1(n_1240),
.B2(n_1163),
.Y(n_1280)
);

O2A1O1Ixp33_ASAP7_75t_L g1281 ( 
.A1(n_1254),
.A2(n_1273),
.B(n_1166),
.C(n_1189),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1236),
.A2(n_1255),
.B1(n_1240),
.B2(n_1163),
.Y(n_1282)
);

O2A1O1Ixp5_ASAP7_75t_L g1283 ( 
.A1(n_1271),
.A2(n_1179),
.B(n_1263),
.C(n_1186),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_SL g1284 ( 
.A1(n_1172),
.A2(n_1250),
.B(n_1237),
.Y(n_1284)
);

NOR2xp67_ASAP7_75t_L g1285 ( 
.A(n_1173),
.B(n_1193),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1168),
.B(n_1261),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1174),
.B(n_1175),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1164),
.A2(n_1179),
.B1(n_1247),
.B2(n_1253),
.Y(n_1288)
);

O2A1O1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1263),
.A2(n_1266),
.B(n_1232),
.C(n_1177),
.Y(n_1289)
);

OA22x2_ASAP7_75t_L g1290 ( 
.A1(n_1209),
.A2(n_1221),
.B1(n_1268),
.B2(n_1260),
.Y(n_1290)
);

NAND2x1p5_ASAP7_75t_L g1291 ( 
.A(n_1190),
.B(n_1207),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1260),
.B(n_1268),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1164),
.A2(n_1253),
.B1(n_1247),
.B2(n_1206),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1201),
.B(n_1196),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1244),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1204),
.B(n_1268),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1188),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1197),
.A2(n_1250),
.B1(n_1172),
.B2(n_1237),
.Y(n_1298)
);

O2A1O1Ixp5_ASAP7_75t_L g1299 ( 
.A1(n_1267),
.A2(n_1276),
.B(n_1274),
.C(n_1199),
.Y(n_1299)
);

INVx1_ASAP7_75t_SL g1300 ( 
.A(n_1239),
.Y(n_1300)
);

OA22x2_ASAP7_75t_L g1301 ( 
.A1(n_1171),
.A2(n_1270),
.B1(n_1251),
.B2(n_1210),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1242),
.B(n_1246),
.Y(n_1302)
);

NOR2x1_ASAP7_75t_SL g1303 ( 
.A(n_1187),
.B(n_1238),
.Y(n_1303)
);

O2A1O1Ixp33_ASAP7_75t_L g1304 ( 
.A1(n_1195),
.A2(n_1193),
.B(n_1245),
.C(n_1187),
.Y(n_1304)
);

AND2x4_ASAP7_75t_SL g1305 ( 
.A(n_1194),
.B(n_1205),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1161),
.Y(n_1306)
);

O2A1O1Ixp5_ASAP7_75t_L g1307 ( 
.A1(n_1211),
.A2(n_1229),
.B(n_1212),
.C(n_1231),
.Y(n_1307)
);

INVxp67_ASAP7_75t_SL g1308 ( 
.A(n_1204),
.Y(n_1308)
);

NAND2xp33_ASAP7_75t_SL g1309 ( 
.A(n_1262),
.B(n_1225),
.Y(n_1309)
);

INVx1_ASAP7_75t_SL g1310 ( 
.A(n_1183),
.Y(n_1310)
);

OA22x2_ASAP7_75t_L g1311 ( 
.A1(n_1241),
.A2(n_1258),
.B1(n_1264),
.B2(n_1222),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1220),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1194),
.B(n_1205),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_1205),
.B(n_1183),
.Y(n_1314)
);

CKINVDCx16_ASAP7_75t_R g1315 ( 
.A(n_1262),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1220),
.A2(n_1227),
.B1(n_1217),
.B2(n_1225),
.Y(n_1316)
);

BUFx3_ASAP7_75t_L g1317 ( 
.A(n_1244),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_SL g1318 ( 
.A1(n_1226),
.A2(n_1187),
.B(n_1238),
.Y(n_1318)
);

O2A1O1Ixp33_ASAP7_75t_L g1319 ( 
.A1(n_1238),
.A2(n_1208),
.B(n_1167),
.C(n_1213),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_SL g1320 ( 
.A(n_1277),
.B(n_1167),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1216),
.B(n_1249),
.Y(n_1321)
);

AOI221xp5_ASAP7_75t_L g1322 ( 
.A1(n_1160),
.A2(n_1272),
.B1(n_1256),
.B2(n_1214),
.C(n_1269),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1208),
.B(n_1235),
.Y(n_1323)
);

OA21x2_ASAP7_75t_L g1324 ( 
.A1(n_1233),
.A2(n_1192),
.B(n_1200),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1223),
.A2(n_1185),
.B1(n_1269),
.B2(n_1161),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1185),
.A2(n_1243),
.B1(n_1248),
.B2(n_1203),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1176),
.B(n_1235),
.Y(n_1327)
);

AOI21x1_ASAP7_75t_SL g1328 ( 
.A1(n_1181),
.A2(n_1190),
.B(n_1249),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1218),
.B(n_1235),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1203),
.A2(n_1218),
.B1(n_1184),
.B2(n_1198),
.Y(n_1330)
);

OA21x2_ASAP7_75t_L g1331 ( 
.A1(n_1230),
.A2(n_1165),
.B(n_1215),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1184),
.A2(n_1198),
.B1(n_1235),
.B2(n_1176),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1176),
.B(n_1228),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1198),
.A2(n_1176),
.B1(n_1202),
.B2(n_1169),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1224),
.B(n_1219),
.Y(n_1335)
);

AOI21x1_ASAP7_75t_SL g1336 ( 
.A1(n_1191),
.A2(n_1162),
.B(n_1275),
.Y(n_1336)
);

AOI21x1_ASAP7_75t_SL g1337 ( 
.A1(n_1252),
.A2(n_1257),
.B(n_1259),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1236),
.A2(n_1255),
.B1(n_1240),
.B2(n_1163),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1178),
.B(n_1182),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1180),
.B(n_1170),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_SL g1341 ( 
.A1(n_1254),
.A2(n_1273),
.B(n_1131),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1236),
.A2(n_1255),
.B1(n_1240),
.B2(n_1163),
.Y(n_1342)
);

A2O1A1Ixp33_ASAP7_75t_SL g1343 ( 
.A1(n_1166),
.A2(n_630),
.B(n_670),
.C(n_995),
.Y(n_1343)
);

A2O1A1Ixp33_ASAP7_75t_L g1344 ( 
.A1(n_1265),
.A2(n_1166),
.B(n_754),
.C(n_1254),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1180),
.B(n_1170),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1180),
.B(n_1170),
.Y(n_1346)
);

OA21x2_ASAP7_75t_L g1347 ( 
.A1(n_1233),
.A2(n_1199),
.B(n_1130),
.Y(n_1347)
);

NOR2x1_ASAP7_75t_SL g1348 ( 
.A(n_1187),
.B(n_1238),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1161),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1174),
.B(n_1175),
.Y(n_1350)
);

INVxp67_ASAP7_75t_SL g1351 ( 
.A(n_1206),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1178),
.B(n_1182),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_SL g1353 ( 
.A1(n_1254),
.A2(n_1273),
.B(n_1131),
.Y(n_1353)
);

OAI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1344),
.A2(n_1279),
.B(n_1281),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1351),
.B(n_1308),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1288),
.B(n_1293),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_1295),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1341),
.A2(n_1353),
.B(n_1289),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1301),
.Y(n_1359)
);

INVx3_ASAP7_75t_L g1360 ( 
.A(n_1331),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1331),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1311),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1335),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1334),
.Y(n_1364)
);

INVx2_ASAP7_75t_SL g1365 ( 
.A(n_1333),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1324),
.Y(n_1366)
);

INVxp67_ASAP7_75t_L g1367 ( 
.A(n_1321),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1297),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1291),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1312),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_SL g1371 ( 
.A1(n_1319),
.A2(n_1338),
.B(n_1280),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1299),
.A2(n_1307),
.B(n_1283),
.Y(n_1372)
);

BUFx2_ASAP7_75t_L g1373 ( 
.A(n_1322),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1324),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1303),
.B(n_1348),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1347),
.B(n_1325),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1326),
.B(n_1296),
.Y(n_1377)
);

NAND3xp33_ASAP7_75t_L g1378 ( 
.A(n_1343),
.B(n_1288),
.C(n_1280),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_1317),
.Y(n_1379)
);

OA21x2_ASAP7_75t_L g1380 ( 
.A1(n_1287),
.A2(n_1350),
.B(n_1332),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1287),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1292),
.Y(n_1382)
);

OR2x2_ASAP7_75t_L g1383 ( 
.A(n_1326),
.B(n_1330),
.Y(n_1383)
);

INVx2_ASAP7_75t_SL g1384 ( 
.A(n_1330),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1318),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1286),
.Y(n_1386)
);

OA21x2_ASAP7_75t_L g1387 ( 
.A1(n_1282),
.A2(n_1342),
.B(n_1338),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1290),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1290),
.B(n_1346),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1294),
.Y(n_1390)
);

INVxp67_ASAP7_75t_SL g1391 ( 
.A(n_1304),
.Y(n_1391)
);

INVx3_ASAP7_75t_L g1392 ( 
.A(n_1323),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1339),
.B(n_1352),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1294),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1336),
.A2(n_1337),
.B(n_1328),
.Y(n_1395)
);

AO21x2_ASAP7_75t_L g1396 ( 
.A1(n_1282),
.A2(n_1342),
.B(n_1316),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1316),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_SL g1398 ( 
.A(n_1293),
.B(n_1298),
.Y(n_1398)
);

AND2x4_ASAP7_75t_L g1399 ( 
.A(n_1375),
.B(n_1327),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1381),
.B(n_1345),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1367),
.B(n_1363),
.Y(n_1401)
);

INVx4_ASAP7_75t_SL g1402 ( 
.A(n_1388),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1382),
.B(n_1340),
.Y(n_1403)
);

INVx5_ASAP7_75t_L g1404 ( 
.A(n_1360),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1367),
.B(n_1300),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1375),
.Y(n_1406)
);

OAI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1378),
.A2(n_1315),
.B1(n_1285),
.B2(n_1298),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1375),
.B(n_1313),
.Y(n_1408)
);

BUFx12f_ASAP7_75t_L g1409 ( 
.A(n_1357),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1361),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1363),
.B(n_1310),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1382),
.B(n_1302),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1356),
.A2(n_1309),
.B1(n_1314),
.B2(n_1320),
.Y(n_1413)
);

INVxp67_ASAP7_75t_L g1414 ( 
.A(n_1377),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1389),
.B(n_1305),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1389),
.B(n_1329),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1368),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1356),
.A2(n_1349),
.B1(n_1306),
.B2(n_1278),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1368),
.Y(n_1419)
);

BUFx2_ASAP7_75t_L g1420 ( 
.A(n_1369),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1370),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1365),
.B(n_1349),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1361),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1381),
.B(n_1284),
.Y(n_1424)
);

BUFx3_ASAP7_75t_L g1425 ( 
.A(n_1409),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1399),
.B(n_1375),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1417),
.Y(n_1427)
);

INVx3_ASAP7_75t_R g1428 ( 
.A(n_1405),
.Y(n_1428)
);

NAND3xp33_ASAP7_75t_L g1429 ( 
.A(n_1414),
.B(n_1378),
.C(n_1358),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1409),
.B(n_1386),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1414),
.B(n_1386),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_R g1432 ( 
.A(n_1409),
.B(n_1357),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1417),
.Y(n_1433)
);

NAND3xp33_ASAP7_75t_L g1434 ( 
.A(n_1407),
.B(n_1358),
.C(n_1354),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1412),
.B(n_1355),
.Y(n_1435)
);

AOI222xp33_ASAP7_75t_L g1436 ( 
.A1(n_1407),
.A2(n_1354),
.B1(n_1398),
.B2(n_1391),
.C1(n_1373),
.C2(n_1388),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1411),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1399),
.B(n_1392),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_R g1439 ( 
.A(n_1424),
.B(n_1379),
.Y(n_1439)
);

AOI222xp33_ASAP7_75t_L g1440 ( 
.A1(n_1400),
.A2(n_1398),
.B1(n_1391),
.B2(n_1373),
.C1(n_1388),
.C2(n_1397),
.Y(n_1440)
);

NAND3xp33_ASAP7_75t_L g1441 ( 
.A(n_1413),
.B(n_1371),
.C(n_1387),
.Y(n_1441)
);

AO31x2_ASAP7_75t_L g1442 ( 
.A1(n_1420),
.A2(n_1373),
.A3(n_1361),
.B(n_1366),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1418),
.A2(n_1387),
.B1(n_1388),
.B2(n_1383),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1399),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_SL g1445 ( 
.A1(n_1416),
.A2(n_1387),
.B1(n_1396),
.B2(n_1383),
.Y(n_1445)
);

CKINVDCx16_ASAP7_75t_R g1446 ( 
.A(n_1415),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1401),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1419),
.Y(n_1448)
);

OAI31xp33_ASAP7_75t_SL g1449 ( 
.A1(n_1408),
.A2(n_1385),
.A3(n_1375),
.B(n_1387),
.Y(n_1449)
);

OR2x6_ASAP7_75t_L g1450 ( 
.A(n_1411),
.B(n_1385),
.Y(n_1450)
);

OAI33xp33_ASAP7_75t_L g1451 ( 
.A1(n_1400),
.A2(n_1359),
.A3(n_1362),
.B1(n_1390),
.B2(n_1394),
.B3(n_1393),
.Y(n_1451)
);

NAND3xp33_ASAP7_75t_L g1452 ( 
.A(n_1421),
.B(n_1377),
.C(n_1364),
.Y(n_1452)
);

NAND2xp33_ASAP7_75t_R g1453 ( 
.A(n_1422),
.B(n_1379),
.Y(n_1453)
);

INVx5_ASAP7_75t_L g1454 ( 
.A(n_1404),
.Y(n_1454)
);

AO21x2_ASAP7_75t_L g1455 ( 
.A1(n_1410),
.A2(n_1374),
.B(n_1366),
.Y(n_1455)
);

OR2x6_ASAP7_75t_L g1456 ( 
.A(n_1406),
.B(n_1385),
.Y(n_1456)
);

OAI221xp5_ASAP7_75t_L g1457 ( 
.A1(n_1406),
.A2(n_1393),
.B1(n_1385),
.B2(n_1384),
.C(n_1362),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_SL g1458 ( 
.A1(n_1416),
.A2(n_1396),
.B1(n_1384),
.B2(n_1380),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1427),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1433),
.Y(n_1460)
);

INVxp67_ASAP7_75t_SL g1461 ( 
.A(n_1429),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1455),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1448),
.Y(n_1463)
);

BUFx2_ASAP7_75t_L g1464 ( 
.A(n_1442),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1442),
.B(n_1410),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1454),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1447),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1439),
.B(n_1402),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1431),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1454),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1454),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1452),
.B(n_1410),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1450),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1443),
.A2(n_1360),
.B(n_1395),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1450),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1450),
.Y(n_1476)
);

OA21x2_ASAP7_75t_L g1477 ( 
.A1(n_1457),
.A2(n_1374),
.B(n_1423),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1456),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1428),
.Y(n_1479)
);

NAND3xp33_ASAP7_75t_SL g1480 ( 
.A(n_1436),
.B(n_1376),
.C(n_1394),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1437),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1437),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1437),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1456),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1465),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1461),
.B(n_1469),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1461),
.B(n_1440),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1478),
.B(n_1426),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1459),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1479),
.B(n_1478),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1465),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1480),
.A2(n_1434),
.B1(n_1396),
.B2(n_1441),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1461),
.B(n_1458),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1479),
.B(n_1426),
.Y(n_1494)
);

BUFx2_ASAP7_75t_L g1495 ( 
.A(n_1478),
.Y(n_1495)
);

NOR2xp67_ASAP7_75t_L g1496 ( 
.A(n_1466),
.B(n_1404),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1459),
.Y(n_1497)
);

INVx3_ASAP7_75t_SL g1498 ( 
.A(n_1468),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1459),
.Y(n_1499)
);

INVx1_ASAP7_75t_SL g1500 ( 
.A(n_1481),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1460),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1467),
.B(n_1435),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1478),
.B(n_1444),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1465),
.Y(n_1504)
);

BUFx2_ASAP7_75t_L g1505 ( 
.A(n_1478),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1460),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1484),
.B(n_1446),
.Y(n_1507)
);

NOR2x1_ASAP7_75t_L g1508 ( 
.A(n_1480),
.B(n_1425),
.Y(n_1508)
);

AOI221xp5_ASAP7_75t_L g1509 ( 
.A1(n_1480),
.A2(n_1441),
.B1(n_1451),
.B2(n_1445),
.C(n_1430),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1484),
.B(n_1438),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1460),
.Y(n_1511)
);

INVx5_ASAP7_75t_L g1512 ( 
.A(n_1466),
.Y(n_1512)
);

NAND2x1p5_ASAP7_75t_L g1513 ( 
.A(n_1466),
.B(n_1372),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1465),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1462),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1467),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1473),
.B(n_1449),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1469),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1472),
.B(n_1401),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1481),
.B(n_1403),
.Y(n_1520)
);

NOR2x1_ASAP7_75t_R g1521 ( 
.A(n_1468),
.B(n_1306),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1463),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1462),
.Y(n_1523)
);

NAND3xp33_ASAP7_75t_L g1524 ( 
.A(n_1477),
.B(n_1372),
.C(n_1364),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1515),
.Y(n_1525)
);

NOR2x1_ASAP7_75t_L g1526 ( 
.A(n_1508),
.B(n_1466),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1487),
.B(n_1481),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1516),
.B(n_1472),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1498),
.B(n_1482),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1489),
.Y(n_1530)
);

INVx2_ASAP7_75t_SL g1531 ( 
.A(n_1512),
.Y(n_1531)
);

NOR2xp67_ASAP7_75t_L g1532 ( 
.A(n_1512),
.B(n_1473),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1490),
.B(n_1509),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1489),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1498),
.B(n_1475),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1497),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1498),
.B(n_1475),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1490),
.B(n_1475),
.Y(n_1538)
);

NAND4xp75_ASAP7_75t_L g1539 ( 
.A(n_1508),
.B(n_1477),
.C(n_1470),
.D(n_1471),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1497),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1507),
.B(n_1475),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1493),
.B(n_1492),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1499),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_SL g1544 ( 
.A(n_1493),
.B(n_1432),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1515),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1486),
.B(n_1472),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1486),
.B(n_1472),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1499),
.Y(n_1548)
);

NOR2x1_ASAP7_75t_L g1549 ( 
.A(n_1495),
.B(n_1466),
.Y(n_1549)
);

INVxp67_ASAP7_75t_L g1550 ( 
.A(n_1495),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1501),
.Y(n_1551)
);

NOR3xp33_ASAP7_75t_L g1552 ( 
.A(n_1505),
.B(n_1466),
.C(n_1474),
.Y(n_1552)
);

NOR2x1_ASAP7_75t_L g1553 ( 
.A(n_1505),
.B(n_1466),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1501),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1506),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1506),
.Y(n_1556)
);

INVx2_ASAP7_75t_SL g1557 ( 
.A(n_1512),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1511),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1507),
.B(n_1482),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1535),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1530),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1533),
.B(n_1494),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1534),
.Y(n_1563)
);

INVxp67_ASAP7_75t_L g1564 ( 
.A(n_1529),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1541),
.B(n_1494),
.Y(n_1565)
);

NOR2x1_ASAP7_75t_L g1566 ( 
.A(n_1526),
.B(n_1500),
.Y(n_1566)
);

INVxp67_ASAP7_75t_L g1567 ( 
.A(n_1529),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1541),
.B(n_1510),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1535),
.B(n_1537),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1550),
.B(n_1517),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1528),
.B(n_1518),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1536),
.Y(n_1572)
);

CKINVDCx16_ASAP7_75t_R g1573 ( 
.A(n_1537),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1540),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1543),
.Y(n_1575)
);

INVx4_ASAP7_75t_L g1576 ( 
.A(n_1531),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_1544),
.Y(n_1577)
);

INVxp67_ASAP7_75t_SL g1578 ( 
.A(n_1549),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1538),
.B(n_1510),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1548),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1551),
.Y(n_1581)
);

AOI221xp5_ASAP7_75t_L g1582 ( 
.A1(n_1542),
.A2(n_1524),
.B1(n_1517),
.B2(n_1464),
.C(n_1500),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1538),
.B(n_1503),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1554),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1571),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1577),
.B(n_1544),
.Y(n_1586)
);

AOI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1573),
.A2(n_1539),
.B1(n_1559),
.B2(n_1527),
.Y(n_1587)
);

NOR2x1_ASAP7_75t_L g1588 ( 
.A(n_1566),
.B(n_1576),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1576),
.Y(n_1589)
);

O2A1O1Ixp5_ASAP7_75t_L g1590 ( 
.A1(n_1578),
.A2(n_1546),
.B(n_1547),
.C(n_1528),
.Y(n_1590)
);

AO22x1_ASAP7_75t_L g1591 ( 
.A1(n_1569),
.A2(n_1553),
.B1(n_1512),
.B2(n_1552),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1576),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1571),
.Y(n_1593)
);

AOI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1582),
.A2(n_1503),
.B1(n_1488),
.B2(n_1532),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1569),
.B(n_1560),
.Y(n_1595)
);

AOI211xp5_ASAP7_75t_L g1596 ( 
.A1(n_1562),
.A2(n_1521),
.B(n_1546),
.C(n_1547),
.Y(n_1596)
);

OAI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1570),
.A2(n_1524),
.B1(n_1453),
.B2(n_1557),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1572),
.Y(n_1598)
);

OAI21xp5_ASAP7_75t_SL g1599 ( 
.A1(n_1564),
.A2(n_1488),
.B(n_1557),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1572),
.Y(n_1600)
);

INVx1_ASAP7_75t_SL g1601 ( 
.A(n_1583),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1567),
.B(n_1555),
.Y(n_1602)
);

AOI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1565),
.A2(n_1488),
.B1(n_1396),
.B2(n_1531),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1588),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1601),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1601),
.B(n_1565),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1585),
.B(n_1583),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1593),
.B(n_1568),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1595),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1589),
.B(n_1568),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1592),
.B(n_1579),
.Y(n_1611)
);

INVx1_ASAP7_75t_SL g1612 ( 
.A(n_1586),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1598),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1596),
.B(n_1579),
.Y(n_1614)
);

INVxp67_ASAP7_75t_L g1615 ( 
.A(n_1602),
.Y(n_1615)
);

OAI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1615),
.A2(n_1590),
.B(n_1594),
.Y(n_1616)
);

O2A1O1Ixp33_ASAP7_75t_L g1617 ( 
.A1(n_1604),
.A2(n_1602),
.B(n_1597),
.C(n_1600),
.Y(n_1617)
);

AOI221xp5_ASAP7_75t_L g1618 ( 
.A1(n_1612),
.A2(n_1587),
.B1(n_1591),
.B2(n_1599),
.C(n_1575),
.Y(n_1618)
);

O2A1O1Ixp33_ASAP7_75t_L g1619 ( 
.A1(n_1604),
.A2(n_1574),
.B(n_1581),
.C(n_1561),
.Y(n_1619)
);

AOI211xp5_ASAP7_75t_L g1620 ( 
.A1(n_1606),
.A2(n_1563),
.B(n_1584),
.C(n_1580),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1610),
.B(n_1580),
.Y(n_1621)
);

OAI31xp33_ASAP7_75t_L g1622 ( 
.A1(n_1614),
.A2(n_1584),
.A3(n_1464),
.B(n_1471),
.Y(n_1622)
);

AOI322xp5_ASAP7_75t_L g1623 ( 
.A1(n_1615),
.A2(n_1603),
.A3(n_1464),
.B1(n_1556),
.B2(n_1558),
.C1(n_1485),
.C2(n_1504),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1608),
.Y(n_1624)
);

AOI211xp5_ASAP7_75t_L g1625 ( 
.A1(n_1616),
.A2(n_1605),
.B(n_1609),
.C(n_1611),
.Y(n_1625)
);

OAI21xp5_ASAP7_75t_SL g1626 ( 
.A1(n_1618),
.A2(n_1607),
.B(n_1611),
.Y(n_1626)
);

NAND5xp2_ASAP7_75t_L g1627 ( 
.A(n_1617),
.B(n_1613),
.C(n_1610),
.D(n_1513),
.E(n_1482),
.Y(n_1627)
);

INVxp33_ASAP7_75t_SL g1628 ( 
.A(n_1624),
.Y(n_1628)
);

AOI211xp5_ASAP7_75t_L g1629 ( 
.A1(n_1622),
.A2(n_1610),
.B(n_1521),
.C(n_1496),
.Y(n_1629)
);

NAND2x1p5_ASAP7_75t_L g1630 ( 
.A(n_1628),
.B(n_1621),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1629),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1625),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1626),
.B(n_1620),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1627),
.B(n_1619),
.Y(n_1634)
);

OAI311xp33_ASAP7_75t_L g1635 ( 
.A1(n_1626),
.A2(n_1623),
.A3(n_1519),
.B1(n_1502),
.C1(n_1483),
.Y(n_1635)
);

BUFx3_ASAP7_75t_L g1636 ( 
.A(n_1630),
.Y(n_1636)
);

NAND4xp25_ASAP7_75t_SL g1637 ( 
.A(n_1634),
.B(n_1545),
.C(n_1525),
.D(n_1470),
.Y(n_1637)
);

CKINVDCx20_ASAP7_75t_R g1638 ( 
.A(n_1633),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1632),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1632),
.B(n_1512),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1636),
.Y(n_1641)
);

NAND4xp75_ASAP7_75t_L g1642 ( 
.A(n_1640),
.B(n_1631),
.C(n_1635),
.D(n_1496),
.Y(n_1642)
);

NOR4xp75_ASAP7_75t_SL g1643 ( 
.A(n_1637),
.B(n_1512),
.C(n_1520),
.D(n_1525),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1641),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1644),
.B(n_1639),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1645),
.Y(n_1646)
);

AOI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1646),
.A2(n_1638),
.B(n_1643),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1647),
.Y(n_1648)
);

CKINVDCx20_ASAP7_75t_R g1649 ( 
.A(n_1648),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1648),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1650),
.A2(n_1642),
.B1(n_1545),
.B2(n_1523),
.Y(n_1651)
);

AOI221xp5_ASAP7_75t_L g1652 ( 
.A1(n_1649),
.A2(n_1523),
.B1(n_1515),
.B2(n_1485),
.C(n_1504),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1651),
.B(n_1470),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1652),
.A2(n_1491),
.B1(n_1485),
.B2(n_1504),
.Y(n_1654)
);

AOI22x1_ASAP7_75t_L g1655 ( 
.A1(n_1653),
.A2(n_1523),
.B1(n_1349),
.B2(n_1491),
.Y(n_1655)
);

AOI322xp5_ASAP7_75t_L g1656 ( 
.A1(n_1654),
.A2(n_1491),
.A3(n_1514),
.B1(n_1470),
.B2(n_1471),
.C1(n_1464),
.C2(n_1476),
.Y(n_1656)
);

AOI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1655),
.A2(n_1514),
.B1(n_1488),
.B2(n_1522),
.Y(n_1657)
);

AOI211xp5_ASAP7_75t_L g1658 ( 
.A1(n_1657),
.A2(n_1656),
.B(n_1470),
.C(n_1471),
.Y(n_1658)
);


endmodule