module fake_ariane_1982_n_382 (n_8, n_56, n_24, n_7, n_22, n_43, n_1, n_49, n_6, n_13, n_20, n_27, n_48, n_29, n_17, n_4, n_41, n_50, n_38, n_55, n_2, n_47, n_18, n_32, n_28, n_37, n_58, n_9, n_51, n_45, n_11, n_34, n_26, n_3, n_46, n_14, n_0, n_52, n_36, n_33, n_44, n_19, n_30, n_39, n_40, n_31, n_42, n_57, n_16, n_5, n_12, n_15, n_53, n_21, n_23, n_35, n_10, n_54, n_25, n_382);

input n_8;
input n_56;
input n_24;
input n_7;
input n_22;
input n_43;
input n_1;
input n_49;
input n_6;
input n_13;
input n_20;
input n_27;
input n_48;
input n_29;
input n_17;
input n_4;
input n_41;
input n_50;
input n_38;
input n_55;
input n_2;
input n_47;
input n_18;
input n_32;
input n_28;
input n_37;
input n_58;
input n_9;
input n_51;
input n_45;
input n_11;
input n_34;
input n_26;
input n_3;
input n_46;
input n_14;
input n_0;
input n_52;
input n_36;
input n_33;
input n_44;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_42;
input n_57;
input n_16;
input n_5;
input n_12;
input n_15;
input n_53;
input n_21;
input n_23;
input n_35;
input n_10;
input n_54;
input n_25;

output n_382;

wire n_295;
wire n_356;
wire n_170;
wire n_190;
wire n_160;
wire n_64;
wire n_180;
wire n_119;
wire n_124;
wire n_307;
wire n_332;
wire n_294;
wire n_197;
wire n_176;
wire n_172;
wire n_347;
wire n_183;
wire n_373;
wire n_299;
wire n_133;
wire n_66;
wire n_205;
wire n_341;
wire n_71;
wire n_109;
wire n_245;
wire n_96;
wire n_319;
wire n_283;
wire n_187;
wire n_367;
wire n_345;
wire n_374;
wire n_318;
wire n_103;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_370;
wire n_189;
wire n_286;
wire n_72;
wire n_117;
wire n_139;
wire n_85;
wire n_130;
wire n_349;
wire n_346;
wire n_214;
wire n_348;
wire n_379;
wire n_138;
wire n_162;
wire n_264;
wire n_137;
wire n_122;
wire n_198;
wire n_232;
wire n_73;
wire n_327;
wire n_77;
wire n_372;
wire n_377;
wire n_87;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_59;
wire n_336;
wire n_315;
wire n_311;
wire n_239;
wire n_272;
wire n_339;
wire n_167;
wire n_90;
wire n_153;
wire n_269;
wire n_75;
wire n_158;
wire n_69;
wire n_259;
wire n_95;
wire n_143;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_173;
wire n_242;
wire n_309;
wire n_331;
wire n_115;
wire n_320;
wire n_267;
wire n_335;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_62;
wire n_210;
wire n_200;
wire n_166;
wire n_253;
wire n_218;
wire n_79;
wire n_271;
wire n_247;
wire n_91;
wire n_240;
wire n_369;
wire n_128;
wire n_224;
wire n_82;
wire n_222;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_330;
wire n_129;
wire n_126;
wire n_282;
wire n_328;
wire n_368;
wire n_301;
wire n_248;
wire n_277;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_93;
wire n_108;
wire n_303;
wire n_168;
wire n_81;
wire n_206;
wire n_352;
wire n_238;
wire n_365;
wire n_136;
wire n_334;
wire n_192;
wire n_300;
wire n_163;
wire n_88;
wire n_141;
wire n_104;
wire n_314;
wire n_273;
wire n_305;
wire n_312;
wire n_233;
wire n_60;
wire n_333;
wire n_376;
wire n_221;
wire n_321;
wire n_86;
wire n_361;
wire n_89;
wire n_149;
wire n_237;
wire n_175;
wire n_74;
wire n_181;
wire n_260;
wire n_362;
wire n_310;
wire n_236;
wire n_281;
wire n_209;
wire n_262;
wire n_225;
wire n_235;
wire n_297;
wire n_290;
wire n_84;
wire n_371;
wire n_199;
wire n_107;
wire n_217;
wire n_178;
wire n_308;
wire n_201;
wire n_70;
wire n_343;
wire n_287;
wire n_302;
wire n_380;
wire n_94;
wire n_284;
wire n_249;
wire n_65;
wire n_123;
wire n_212;
wire n_355;
wire n_278;
wire n_255;
wire n_257;
wire n_148;
wire n_135;
wire n_171;
wire n_61;
wire n_102;
wire n_182;
wire n_316;
wire n_196;
wire n_125;
wire n_254;
wire n_219;
wire n_231;
wire n_366;
wire n_234;
wire n_280;
wire n_215;
wire n_252;
wire n_161;
wire n_298;
wire n_68;
wire n_78;
wire n_63;
wire n_99;
wire n_216;
wire n_223;
wire n_83;
wire n_288;
wire n_179;
wire n_195;
wire n_213;
wire n_110;
wire n_304;
wire n_67;
wire n_306;
wire n_313;
wire n_92;
wire n_203;
wire n_378;
wire n_150;
wire n_98;
wire n_375;
wire n_113;
wire n_114;
wire n_324;
wire n_337;
wire n_111;
wire n_274;
wire n_296;
wire n_265;
wire n_208;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_100;
wire n_132;
wire n_147;
wire n_204;
wire n_76;
wire n_342;
wire n_246;
wire n_159;
wire n_358;
wire n_105;
wire n_131;
wire n_263;
wire n_360;
wire n_229;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_101;
wire n_243;
wire n_134;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_112;
wire n_268;
wire n_266;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_364;
wire n_258;
wire n_118;
wire n_121;
wire n_353;
wire n_241;
wire n_357;
wire n_191;
wire n_80;
wire n_211;
wire n_97;
wire n_322;
wire n_251;
wire n_116;
wire n_351;
wire n_359;
wire n_155;
wire n_127;

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_17),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_23),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

CKINVDCx5p33_ASAP7_75t_R g69 ( 
.A(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_12),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

CKINVDCx5p33_ASAP7_75t_R g75 ( 
.A(n_15),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

INVxp67_ASAP7_75t_SL g77 ( 
.A(n_13),
.Y(n_77)
);

INVxp33_ASAP7_75t_SL g78 ( 
.A(n_41),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_14),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

CKINVDCx5p33_ASAP7_75t_R g82 ( 
.A(n_14),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_16),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_12),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_33),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_6),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVxp67_ASAP7_75t_SL g88 ( 
.A(n_2),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_47),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_34),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_11),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_0),
.Y(n_95)
);

INVxp33_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

INVxp67_ASAP7_75t_SL g98 ( 
.A(n_57),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_27),
.Y(n_99)
);

CKINVDCx5p33_ASAP7_75t_R g100 ( 
.A(n_55),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_30),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_32),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_13),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_9),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_0),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_29),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_11),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_3),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_46),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_44),
.Y(n_111)
);

CKINVDCx5p33_ASAP7_75t_R g112 ( 
.A(n_85),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_85),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_74),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_91),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_102),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_R g120 ( 
.A(n_62),
.B(n_18),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g121 ( 
.A(n_75),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_83),
.Y(n_122)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_82),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_104),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_69),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_100),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_74),
.B(n_64),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_65),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

AND3x2_ASAP7_75t_L g134 ( 
.A(n_72),
.B(n_1),
.C(n_4),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_101),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_89),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_99),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_78),
.Y(n_138)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_72),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_60),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_107),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_60),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_63),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_66),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_111),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_111),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_68),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_68),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_110),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_70),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_70),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_71),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_66),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_110),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_71),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_79),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_79),
.B(n_1),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_81),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_81),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_87),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_87),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_117),
.Y(n_162)
);

NAND2x1p5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_97),
.Y(n_163)
);

AO22x2_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_73),
.B1(n_105),
.B2(n_95),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

NAND2x1p5_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_97),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_118),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_103),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_118),
.Y(n_169)
);

AOI22x1_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_88),
.B1(n_77),
.B2(n_108),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_121),
.Y(n_171)
);

AND2x4_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_103),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_108),
.C(n_73),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_96),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_127),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_127),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_131),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_132),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_133),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_123),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_115),
.A2(n_98),
.B1(n_90),
.B2(n_92),
.Y(n_182)
);

NAND2x1_ASAP7_75t_L g183 ( 
.A(n_131),
.B(n_106),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_112),
.Y(n_184)
);

AND2x6_ASAP7_75t_L g185 ( 
.A(n_133),
.B(n_106),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_125),
.B(n_90),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_139),
.B(n_105),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_149),
.B(n_59),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_112),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_131),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_113),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_119),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_131),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_142),
.Y(n_194)
);

AO22x2_ASAP7_75t_L g195 ( 
.A1(n_114),
.A2(n_84),
.B1(n_95),
.B2(n_93),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_147),
.Y(n_196)
);

AND2x4_ASAP7_75t_L g197 ( 
.A(n_147),
.B(n_84),
.Y(n_197)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_115),
.B(n_80),
.C(n_93),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_113),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_136),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_144),
.Y(n_201)
);

NOR2xp67_ASAP7_75t_L g202 ( 
.A(n_126),
.B(n_106),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_135),
.Y(n_203)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_185),
.Y(n_204)
);

AOI222xp33_ASAP7_75t_L g205 ( 
.A1(n_195),
.A2(n_80),
.B1(n_76),
.B2(n_153),
.C1(n_158),
.C2(n_156),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_186),
.A2(n_67),
.B(n_155),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_188),
.Y(n_207)
);

AO32x1_ASAP7_75t_L g208 ( 
.A1(n_177),
.A2(n_155),
.A3(n_92),
.B1(n_94),
.B2(n_59),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_138),
.Y(n_209)
);

NOR2xp67_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_145),
.Y(n_210)
);

O2A1O1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_194),
.A2(n_201),
.B(n_188),
.C(n_162),
.Y(n_211)
);

AO21x2_ASAP7_75t_L g212 ( 
.A1(n_202),
.A2(n_120),
.B(n_94),
.Y(n_212)
);

AND2x6_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_76),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_175),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_159),
.Y(n_215)
);

AOI221xp5_ASAP7_75t_L g216 ( 
.A1(n_195),
.A2(n_146),
.B1(n_148),
.B2(n_154),
.C(n_152),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_139),
.B(n_137),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_190),
.A2(n_139),
.B(n_130),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_192),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_165),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_203),
.B(n_161),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_165),
.Y(n_224)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_185),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_171),
.B(n_160),
.Y(n_226)
);

AO21x2_ASAP7_75t_L g227 ( 
.A1(n_173),
.A2(n_134),
.B(n_150),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_178),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_L g229 ( 
.A1(n_182),
.A2(n_151),
.B(n_143),
.C(n_7),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_178),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_181),
.Y(n_231)
);

O2A1O1Ixp33_ASAP7_75t_L g232 ( 
.A1(n_187),
.A2(n_4),
.B(n_5),
.C(n_7),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_179),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_184),
.B(n_116),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_163),
.B(n_5),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_179),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_180),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_191),
.B(n_124),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_193),
.A2(n_35),
.B(n_56),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_180),
.A2(n_26),
.B(n_51),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_196),
.A2(n_20),
.B(n_43),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_196),
.B(n_166),
.Y(n_242)
);

AO32x1_ASAP7_75t_L g243 ( 
.A1(n_167),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_16),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_199),
.B(n_122),
.Y(n_244)
);

AND2x4_ASAP7_75t_L g245 ( 
.A(n_168),
.B(n_8),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_169),
.Y(n_246)
);

HAxp5_ASAP7_75t_L g247 ( 
.A(n_198),
.B(n_10),
.CON(n_247),
.SN(n_247)
);

OR2x6_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_166),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_207),
.B(n_163),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

OAI21x1_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_170),
.B(n_187),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_209),
.B(n_189),
.Y(n_252)
);

OA21x2_ASAP7_75t_L g253 ( 
.A1(n_242),
.A2(n_197),
.B(n_172),
.Y(n_253)
);

CKINVDCx6p67_ASAP7_75t_R g254 ( 
.A(n_220),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_226),
.A2(n_189),
.B1(n_197),
.B2(n_172),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_215),
.B(n_168),
.Y(n_257)
);

OAI21x1_ASAP7_75t_L g258 ( 
.A1(n_239),
.A2(n_185),
.B(n_195),
.Y(n_258)
);

AOI221x1_ASAP7_75t_L g259 ( 
.A1(n_235),
.A2(n_164),
.B1(n_195),
.B2(n_172),
.C(n_185),
.Y(n_259)
);

OAI21x1_ASAP7_75t_L g260 ( 
.A1(n_206),
.A2(n_185),
.B(n_164),
.Y(n_260)
);

NAND2xp33_ASAP7_75t_R g261 ( 
.A(n_231),
.B(n_164),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_228),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_211),
.A2(n_215),
.B(n_214),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_213),
.Y(n_264)
);

AO31x2_ASAP7_75t_L g265 ( 
.A1(n_236),
.A2(n_38),
.A3(n_39),
.B(n_246),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_218),
.Y(n_266)
);

AO21x2_ASAP7_75t_L g267 ( 
.A1(n_219),
.A2(n_212),
.B(n_217),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_205),
.A2(n_216),
.B1(n_213),
.B2(n_245),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_238),
.Y(n_269)
);

OA21x2_ASAP7_75t_L g270 ( 
.A1(n_240),
.A2(n_241),
.B(n_229),
.Y(n_270)
);

OAI21x1_ASAP7_75t_L g271 ( 
.A1(n_223),
.A2(n_232),
.B(n_210),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_222),
.B(n_244),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_205),
.A2(n_213),
.B1(n_228),
.B2(n_227),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_213),
.B(n_212),
.Y(n_274)
);

AOI221xp5_ASAP7_75t_L g275 ( 
.A1(n_238),
.A2(n_234),
.B1(n_247),
.B2(n_227),
.C(n_223),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_228),
.Y(n_276)
);

NAND3x1_ASAP7_75t_L g277 ( 
.A(n_243),
.B(n_208),
.C(n_204),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_221),
.Y(n_278)
);

OAI21x1_ASAP7_75t_L g279 ( 
.A1(n_208),
.A2(n_204),
.B(n_225),
.Y(n_279)
);

INVxp33_ASAP7_75t_SL g280 ( 
.A(n_204),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_224),
.B(n_204),
.Y(n_281)
);

CKINVDCx6p67_ASAP7_75t_R g282 ( 
.A(n_225),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_L g283 ( 
.A1(n_224),
.A2(n_207),
.B1(n_216),
.B2(n_182),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_213),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_228),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_233),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_230),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_207),
.B(n_210),
.Y(n_288)
);

OA21x2_ASAP7_75t_L g289 ( 
.A1(n_242),
.A2(n_237),
.B(n_233),
.Y(n_289)
);

OR2x6_ASAP7_75t_L g290 ( 
.A(n_248),
.B(n_264),
.Y(n_290)
);

NAND2xp33_ASAP7_75t_R g291 ( 
.A(n_266),
.B(n_252),
.Y(n_291)
);

NAND2xp33_ASAP7_75t_R g292 ( 
.A(n_266),
.B(n_272),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_R g293 ( 
.A(n_254),
.B(n_261),
.Y(n_293)
);

O2A1O1Ixp33_ASAP7_75t_SL g294 ( 
.A1(n_288),
.A2(n_249),
.B(n_263),
.C(n_264),
.Y(n_294)
);

NAND2xp33_ASAP7_75t_SL g295 ( 
.A(n_268),
.B(n_288),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_L g296 ( 
.A1(n_248),
.A2(n_272),
.B1(n_283),
.B2(n_269),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_287),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_254),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_248),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_257),
.B(n_273),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_253),
.B(n_275),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_255),
.B(n_278),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_287),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_250),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_284),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_276),
.Y(n_306)
);

NOR3xp33_ASAP7_75t_SL g307 ( 
.A(n_256),
.B(n_286),
.C(n_274),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_L g308 ( 
.A1(n_259),
.A2(n_285),
.B1(n_262),
.B2(n_276),
.Y(n_308)
);

AND2x2_ASAP7_75t_SL g309 ( 
.A(n_276),
.B(n_270),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_262),
.A2(n_285),
.B1(n_276),
.B2(n_280),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_289),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_271),
.B(n_260),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_289),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_289),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g315 ( 
.A1(n_267),
.A2(n_270),
.B1(n_251),
.B2(n_258),
.Y(n_315)
);

NOR2x1_ASAP7_75t_SL g316 ( 
.A(n_267),
.B(n_281),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_303),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_303),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_267),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_297),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_296),
.B(n_270),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_297),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_309),
.Y(n_323)
);

NAND2xp33_ASAP7_75t_SL g324 ( 
.A(n_291),
.B(n_280),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_309),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g326 ( 
.A(n_290),
.B(n_279),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_300),
.B(n_295),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_301),
.B(n_282),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_309),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_290),
.B(n_279),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_292),
.Y(n_331)
);

OAI211xp5_ASAP7_75t_L g332 ( 
.A1(n_302),
.A2(n_277),
.B(n_265),
.C(n_282),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_290),
.B(n_265),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_304),
.A2(n_265),
.B1(n_277),
.B2(n_290),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_301),
.B(n_265),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_322),
.Y(n_336)
);

OR2x2_ASAP7_75t_L g337 ( 
.A(n_327),
.B(n_314),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_323),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_317),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_327),
.B(n_319),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_319),
.B(n_304),
.Y(n_341)
);

NOR3xp33_ASAP7_75t_L g342 ( 
.A(n_324),
.B(n_298),
.C(n_294),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_323),
.B(n_314),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_317),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_318),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_331),
.B(n_299),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_318),
.B(n_293),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_320),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_320),
.B(n_305),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_321),
.A2(n_298),
.B1(n_305),
.B2(n_307),
.Y(n_350)
);

OAI33xp33_ASAP7_75t_L g351 ( 
.A1(n_347),
.A2(n_334),
.A3(n_308),
.B1(n_335),
.B2(n_310),
.B3(n_328),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_339),
.Y(n_352)
);

OAI33xp33_ASAP7_75t_L g353 ( 
.A1(n_346),
.A2(n_334),
.A3(n_335),
.B1(n_328),
.B2(n_313),
.B3(n_311),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_341),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_344),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_341),
.B(n_340),
.Y(n_356)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_340),
.B(n_329),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_339),
.B(n_329),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_350),
.B(n_306),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_336),
.Y(n_360)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_356),
.B(n_337),
.Y(n_361)
);

AOI211x1_ASAP7_75t_L g362 ( 
.A1(n_355),
.A2(n_349),
.B(n_345),
.C(n_332),
.Y(n_362)
);

AOI322xp5_ASAP7_75t_L g363 ( 
.A1(n_359),
.A2(n_333),
.A3(n_342),
.B1(n_345),
.B2(n_348),
.C1(n_315),
.C2(n_330),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_354),
.Y(n_364)
);

NOR3xp33_ASAP7_75t_L g365 ( 
.A(n_364),
.B(n_351),
.C(n_353),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_361),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_362),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_363),
.Y(n_368)
);

AOI222xp33_ASAP7_75t_L g369 ( 
.A1(n_368),
.A2(n_332),
.B1(n_333),
.B2(n_358),
.C1(n_352),
.C2(n_338),
.Y(n_369)
);

NOR4xp25_ASAP7_75t_L g370 ( 
.A(n_367),
.B(n_352),
.C(n_358),
.D(n_337),
.Y(n_370)
);

AOI221xp5_ASAP7_75t_L g371 ( 
.A1(n_365),
.A2(n_357),
.B1(n_330),
.B2(n_312),
.C(n_326),
.Y(n_371)
);

AOI211xp5_ASAP7_75t_L g372 ( 
.A1(n_366),
.A2(n_357),
.B(n_312),
.C(n_326),
.Y(n_372)
);

AOI222xp33_ASAP7_75t_L g373 ( 
.A1(n_371),
.A2(n_366),
.B1(n_370),
.B2(n_369),
.C1(n_372),
.C2(n_326),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_372),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_370),
.B(n_323),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_374),
.B(n_316),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_375),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_377),
.B(n_376),
.Y(n_378)
);

OAI322xp33_ASAP7_75t_L g379 ( 
.A1(n_378),
.A2(n_373),
.A3(n_375),
.B1(n_343),
.B2(n_325),
.C1(n_329),
.C2(n_360),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_L g380 ( 
.A1(n_379),
.A2(n_325),
.B1(n_360),
.B2(n_326),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_380),
.A2(n_325),
.B1(n_338),
.B2(n_322),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_381),
.A2(n_322),
.B1(n_311),
.B2(n_313),
.Y(n_382)
);


endmodule