module fake_jpeg_20503_n_328 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_23),
.Y(n_37)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NOR2xp67_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_15),
.Y(n_42)
);

NAND2xp33_ASAP7_75t_SL g46 ( 
.A(n_42),
.B(n_23),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NAND3xp33_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_30),
.C(n_29),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_17),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_36),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_17),
.B1(n_26),
.B2(n_22),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_17),
.B1(n_26),
.B2(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_46),
.A2(n_48),
.B(n_50),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_40),
.B1(n_39),
.B2(n_37),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_61),
.A2(n_71),
.B1(n_75),
.B2(n_54),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_51),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_64),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_63),
.A2(n_69),
.B1(n_79),
.B2(n_54),
.Y(n_99)
);

AND2x4_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_37),
.Y(n_65)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_65),
.B(n_74),
.Y(n_100)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_45),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_68),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_26),
.B1(n_16),
.B2(n_40),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_39),
.B1(n_26),
.B2(n_38),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_54),
.A2(n_16),
.B1(n_21),
.B2(n_22),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_43),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_38),
.B1(n_21),
.B2(n_29),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_45),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_76),
.Y(n_95)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_59),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_78),
.A2(n_85),
.B1(n_55),
.B2(n_21),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_52),
.A2(n_38),
.B1(n_21),
.B2(n_29),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_81),
.A2(n_27),
.B1(n_33),
.B2(n_24),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_55),
.Y(n_82)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_47),
.B(n_30),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_83),
.Y(n_107)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_35),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_35),
.Y(n_118)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_91),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_103),
.B1(n_104),
.B2(n_110),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_113),
.B1(n_115),
.B2(n_67),
.Y(n_126)
);

INVxp33_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_60),
.A2(n_65),
.B1(n_62),
.B2(n_64),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_74),
.A2(n_29),
.B1(n_22),
.B2(n_30),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_65),
.A2(n_22),
.B1(n_43),
.B2(n_41),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_77),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_118),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_65),
.A2(n_43),
.B1(n_41),
.B2(n_24),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_87),
.A2(n_19),
.B1(n_32),
.B2(n_31),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_120),
.B(n_31),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_126),
.A2(n_130),
.B1(n_145),
.B2(n_148),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_98),
.A2(n_79),
.B1(n_90),
.B2(n_84),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_127),
.A2(n_136),
.B1(n_94),
.B2(n_27),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_109),
.A2(n_101),
.B(n_100),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_129),
.A2(n_143),
.B(n_144),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_61),
.B1(n_71),
.B2(n_75),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_68),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_133),
.Y(n_174)
);

INVx5_ASAP7_75t_SL g132 ( 
.A(n_111),
.Y(n_132)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_76),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_80),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_134),
.B(n_135),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_88),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_100),
.A2(n_90),
.B1(n_91),
.B2(n_89),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_92),
.B(n_72),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_138),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_35),
.C(n_86),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_96),
.C(n_97),
.Y(n_151)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_114),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_146),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_101),
.A2(n_78),
.B(n_27),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_99),
.A2(n_86),
.B1(n_70),
.B2(n_85),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_92),
.B(n_35),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_113),
.A2(n_95),
.B1(n_112),
.B2(n_110),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_95),
.B(n_41),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_108),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_140),
.A2(n_120),
.B1(n_118),
.B2(n_117),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_150),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_151),
.B(n_164),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_138),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_153),
.Y(n_194)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_96),
.C(n_97),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_122),
.C(n_127),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_114),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_158),
.A2(n_143),
.B(n_140),
.Y(n_183)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_159),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_121),
.Y(n_160)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_126),
.A2(n_148),
.B1(n_130),
.B2(n_145),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_161),
.A2(n_142),
.B1(n_132),
.B2(n_125),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

INVx3_ASAP7_75t_SL g213 ( 
.A(n_162),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_124),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_166),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_119),
.Y(n_164)
);

OAI22x1_ASAP7_75t_SL g165 ( 
.A1(n_122),
.A2(n_105),
.B1(n_108),
.B2(n_82),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_125),
.B1(n_123),
.B2(n_111),
.Y(n_189)
);

AOI32xp33_ASAP7_75t_L g166 ( 
.A1(n_128),
.A2(n_106),
.A3(n_72),
.B1(n_82),
.B2(n_94),
.Y(n_166)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_124),
.Y(n_172)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_172),
.Y(n_211)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_173),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_106),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_175),
.A2(n_179),
.B(n_0),
.Y(n_204)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_176),
.A2(n_182),
.B1(n_169),
.B2(n_179),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_147),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_136),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_181),
.A2(n_165),
.B1(n_182),
.B2(n_158),
.Y(n_187)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_131),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_196),
.Y(n_217)
);

AOI322xp5_ASAP7_75t_L g184 ( 
.A1(n_180),
.A2(n_135),
.A3(n_122),
.B1(n_144),
.B2(n_127),
.C1(n_139),
.C2(n_142),
.Y(n_184)
);

MAJx2_ASAP7_75t_L g225 ( 
.A(n_184),
.B(n_208),
.C(n_214),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_157),
.C(n_163),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_187),
.A2(n_193),
.B1(n_195),
.B2(n_197),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_192),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_156),
.A2(n_123),
.B1(n_111),
.B2(n_33),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_156),
.A2(n_33),
.B1(n_32),
.B2(n_31),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_181),
.A2(n_32),
.B1(n_28),
.B2(n_19),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_158),
.A2(n_28),
.B1(n_19),
.B2(n_15),
.Y(n_195)
);

OAI32xp33_ASAP7_75t_L g196 ( 
.A1(n_174),
.A2(n_20),
.A3(n_25),
.B1(n_18),
.B2(n_23),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_161),
.A2(n_171),
.B1(n_162),
.B2(n_152),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_164),
.A2(n_28),
.B1(n_14),
.B2(n_13),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_198),
.A2(n_206),
.B1(n_207),
.B2(n_25),
.Y(n_237)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_212),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_174),
.A2(n_20),
.B1(n_25),
.B2(n_18),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_150),
.A2(n_25),
.B1(n_18),
.B2(n_2),
.Y(n_207)
);

XNOR2x2_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_25),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_151),
.B(n_25),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_154),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_178),
.A2(n_14),
.B(n_13),
.Y(n_212)
);

A2O1A1O1Ixp25_ASAP7_75t_L g214 ( 
.A1(n_177),
.A2(n_14),
.B(n_12),
.C(n_25),
.D(n_18),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_218),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_176),
.C(n_173),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_223),
.C(n_230),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_170),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_224),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_221),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_170),
.C(n_168),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_168),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_167),
.Y(n_227)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_205),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_207),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_194),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_232),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_186),
.B(n_167),
.C(n_155),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_155),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_234),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_211),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_153),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_185),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_235)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_235),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_25),
.C(n_18),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_238),
.C(n_18),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_203),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_18),
.C(n_12),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_187),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_239)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

NAND3xp33_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_212),
.C(n_201),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_258),
.Y(n_264)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_245),
.A2(n_244),
.B1(n_251),
.B2(n_247),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_228),
.A2(n_191),
.B(n_214),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_249),
.A2(n_3),
.B(n_4),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_221),
.B(n_198),
.Y(n_252)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_226),
.A2(n_188),
.B1(n_217),
.B2(n_231),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_253),
.A2(n_215),
.B1(n_218),
.B2(n_222),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_216),
.B(n_196),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_255),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_190),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_213),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_257),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_215),
.B(n_213),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_260),
.A2(n_11),
.B1(n_4),
.B2(n_5),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_219),
.C(n_220),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_262),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_246),
.C(n_255),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_223),
.C(n_224),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_268),
.Y(n_282)
);

XOR2x2_ASAP7_75t_SL g267 ( 
.A(n_254),
.B(n_225),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_267),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_236),
.C(n_206),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_238),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_272),
.Y(n_279)
);

OAI21xp33_ASAP7_75t_L g272 ( 
.A1(n_243),
.A2(n_225),
.B(n_195),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_192),
.C(n_193),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_275),
.Y(n_291)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_18),
.C(n_4),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_248),
.B(n_3),
.C(n_4),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_8),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_277),
.A2(n_249),
.B(n_240),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_263),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_287),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_280),
.Y(n_296)
);

AOI21xp33_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_256),
.B(n_257),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_283),
.A2(n_267),
.B(n_269),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_270),
.A2(n_253),
.B1(n_258),
.B2(n_5),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_285),
.A2(n_286),
.B1(n_8),
.B2(n_9),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_272),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_290),
.Y(n_298)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_264),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_289),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_7),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_8),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_295),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_262),
.C(n_261),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_269),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_300),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_268),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_290),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_265),
.C(n_9),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_304),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_303),
.A2(n_284),
.B1(n_292),
.B2(n_280),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_11),
.Y(n_304)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_308),
.Y(n_314)
);

NOR2x1_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_288),
.Y(n_309)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_309),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_279),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_310),
.B(n_312),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_279),
.Y(n_311)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_311),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_9),
.C(n_10),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_313),
.B(n_298),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_306),
.A2(n_296),
.B(n_300),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_319),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_317),
.A2(n_312),
.B(n_307),
.Y(n_321)
);

AOI21xp33_ASAP7_75t_L g323 ( 
.A1(n_321),
.A2(n_322),
.B(n_318),
.Y(n_323)
);

BUFx24_ASAP7_75t_SL g322 ( 
.A(n_314),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_323),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_320),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_315),
.B(n_299),
.Y(n_326)
);

O2A1O1Ixp33_ASAP7_75t_SL g327 ( 
.A1(n_326),
.A2(n_309),
.B(n_311),
.C(n_302),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_298),
.B1(n_305),
.B2(n_10),
.Y(n_328)
);


endmodule