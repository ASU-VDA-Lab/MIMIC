module fake_jpeg_5518_n_233 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_233);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_233;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_26),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_0),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_28),
.A2(n_20),
.B1(n_24),
.B2(n_14),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_45),
.B1(n_34),
.B2(n_32),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_30),
.B(n_20),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_48),
.Y(n_51)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_31),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_24),
.B1(n_13),
.B2(n_22),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_49),
.B(n_27),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_27),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_52),
.B(n_54),
.Y(n_79)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_34),
.B1(n_30),
.B2(n_28),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_57),
.B1(n_68),
.B2(n_37),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_30),
.B1(n_32),
.B2(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_29),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_33),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_36),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_60),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_40),
.B1(n_41),
.B2(n_32),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_19),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_50),
.B1(n_39),
.B2(n_32),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

OR2x2_ASAP7_75t_SL g66 ( 
.A(n_49),
.B(n_0),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_66),
.A2(n_67),
.B1(n_50),
.B2(n_46),
.Y(n_76)
);

OR2x2_ASAP7_75t_SL g67 ( 
.A(n_50),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_19),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_69),
.A2(n_78),
.B1(n_83),
.B2(n_88),
.Y(n_102)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_64),
.B(n_51),
.Y(n_107)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_45),
.B1(n_41),
.B2(n_40),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_80),
.A2(n_61),
.B1(n_64),
.B2(n_56),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_81),
.A2(n_68),
.B1(n_65),
.B2(n_51),
.Y(n_90)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

OAI21x1_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_67),
.B(n_51),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_32),
.C(n_41),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_58),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_37),
.B1(n_46),
.B2(n_16),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_57),
.A2(n_37),
.B1(n_46),
.B2(n_44),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_89),
.B(n_84),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_84),
.B1(n_69),
.B2(n_86),
.Y(n_116)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_92),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_70),
.B(n_54),
.Y(n_92)
);

AO21x1_ASAP7_75t_L g93 ( 
.A1(n_73),
.A2(n_51),
.B(n_63),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_93),
.A2(n_98),
.B1(n_100),
.B2(n_99),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_107),
.B1(n_72),
.B2(n_73),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_70),
.B(n_54),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

AND2x4_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_51),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_100),
.A2(n_74),
.B(n_62),
.Y(n_126)
);

BUFx4f_ASAP7_75t_SL g101 ( 
.A(n_73),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_71),
.B(n_60),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_103),
.Y(n_110)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_104),
.A2(n_82),
.B1(n_44),
.B2(n_71),
.Y(n_125)
);

INVxp33_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_74),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_101),
.Y(n_109)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_112),
.B(n_93),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_75),
.B1(n_78),
.B2(n_83),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_114),
.A2(n_116),
.B1(n_104),
.B2(n_97),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_89),
.C(n_87),
.Y(n_139)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_119),
.B(n_120),
.Y(n_127)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_94),
.A2(n_65),
.B1(n_79),
.B2(n_82),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_121),
.A2(n_124),
.B1(n_91),
.B2(n_106),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_79),
.B(n_76),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_122),
.A2(n_126),
.B(n_95),
.Y(n_137)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_125),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_107),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_139),
.C(n_140),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_114),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_118),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_134),
.Y(n_148)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_138),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_136),
.A2(n_142),
.B1(n_66),
.B2(n_29),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_67),
.B(n_109),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_111),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_89),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_53),
.C(n_52),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_143),
.C(n_145),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_119),
.A2(n_105),
.B1(n_95),
.B2(n_97),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_52),
.C(n_59),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_52),
.Y(n_144)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_144),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_52),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_113),
.B1(n_121),
.B2(n_110),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_149),
.B1(n_154),
.B2(n_158),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_146),
.A2(n_113),
.B1(n_126),
.B2(n_116),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_164),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_153),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_129),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_137),
.A2(n_131),
.B1(n_133),
.B2(n_139),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_133),
.A2(n_110),
.B1(n_120),
.B2(n_117),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_159),
.A2(n_160),
.B(n_21),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_128),
.A2(n_144),
.B(n_135),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_66),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_21),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_162),
.A2(n_35),
.B1(n_25),
.B2(n_22),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_134),
.A2(n_136),
.B1(n_142),
.B2(n_130),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_44),
.C(n_29),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_25),
.C(n_22),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_156),
.B(n_130),
.Y(n_166)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_168),
.A2(n_154),
.B1(n_18),
.B2(n_15),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_171),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_35),
.Y(n_170)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_21),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_165),
.C(n_157),
.Y(n_183)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_176),
.Y(n_184)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_178),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_1),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_174),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_149),
.A2(n_25),
.B1(n_18),
.B2(n_15),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_180),
.A2(n_162),
.B1(n_161),
.B2(n_159),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_185),
.C(n_187),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_155),
.C(n_157),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_155),
.C(n_153),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_188),
.A2(n_190),
.B1(n_177),
.B2(n_173),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_18),
.Y(n_190)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_1),
.B(n_2),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_180),
.Y(n_195)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_189),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_196),
.A2(n_199),
.B(n_203),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_167),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_197),
.B(n_201),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_178),
.C(n_177),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_184),
.A2(n_169),
.B(n_12),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_200),
.A2(n_191),
.B(n_192),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_11),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_1),
.C(n_2),
.Y(n_203)
);

NOR2x1_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_190),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_204),
.A2(n_206),
.B(n_209),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_212),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_181),
.Y(n_209)
);

BUFx24_ASAP7_75t_SL g210 ( 
.A(n_203),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_211),
.Y(n_217)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_199),
.Y(n_211)
);

BUFx24_ASAP7_75t_SL g212 ( 
.A(n_194),
.Y(n_212)
);

NOR2xp67_ASAP7_75t_SL g213 ( 
.A(n_208),
.B(n_194),
.Y(n_213)
);

NOR2xp67_ASAP7_75t_SL g221 ( 
.A(n_213),
.B(n_2),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_205),
.A2(n_181),
.B(n_187),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_216),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_205),
.B(n_11),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_205),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_218),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.Y(n_224)
);

A2O1A1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_214),
.A2(n_10),
.B(n_9),
.C(n_4),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_220),
.B(n_222),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_219),
.C(n_3),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_10),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_9),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_227),
.Y(n_229)
);

A2O1A1O1Ixp25_ASAP7_75t_L g228 ( 
.A1(n_225),
.A2(n_223),
.B(n_3),
.C(n_5),
.D(n_7),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_228),
.A2(n_2),
.B(n_3),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_229),
.Y(n_231)
);

OAI32xp33_ASAP7_75t_SL g232 ( 
.A1(n_231),
.A2(n_5),
.A3(n_8),
.B1(n_213),
.B2(n_221),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_232),
.Y(n_233)
);


endmodule