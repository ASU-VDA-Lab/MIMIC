module fake_netlist_1_5952_n_45 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_45);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_25;
wire n_30;
wire n_26;
wire n_16;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
NAND2xp5_ASAP7_75t_L g15 ( .A(n_4), .B(n_1), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_3), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_0), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_12), .Y(n_18) );
BUFx6f_ASAP7_75t_L g19 ( .A(n_10), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_1), .Y(n_20) );
INVx3_ASAP7_75t_L g21 ( .A(n_8), .Y(n_21) );
INVx3_ASAP7_75t_L g22 ( .A(n_7), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_6), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_18), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_21), .B(n_0), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_17), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_20), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g28 ( .A(n_21), .B(n_2), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_22), .B(n_2), .Y(n_29) );
INVx2_ASAP7_75t_L g30 ( .A(n_26), .Y(n_30) );
INVx6_ASAP7_75t_L g31 ( .A(n_27), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_25), .Y(n_32) );
OR2x2_ASAP7_75t_L g33 ( .A(n_32), .B(n_24), .Y(n_33) );
AND2x2_ASAP7_75t_L g34 ( .A(n_31), .B(n_24), .Y(n_34) );
NAND4xp25_ASAP7_75t_SL g35 ( .A(n_30), .B(n_29), .C(n_28), .D(n_15), .Y(n_35) );
NOR2xp33_ASAP7_75t_L g36 ( .A(n_33), .B(n_31), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_34), .Y(n_37) );
AND2x2_ASAP7_75t_L g38 ( .A(n_37), .B(n_15), .Y(n_38) );
O2A1O1Ixp33_ASAP7_75t_L g39 ( .A1(n_36), .A2(n_23), .B(n_35), .C(n_22), .Y(n_39) );
INVx2_ASAP7_75t_L g40 ( .A(n_38), .Y(n_40) );
NOR2xp33_ASAP7_75t_R g41 ( .A(n_39), .B(n_16), .Y(n_41) );
NAND2xp5_ASAP7_75t_L g42 ( .A(n_40), .B(n_19), .Y(n_42) );
OAI222xp33_ASAP7_75t_L g43 ( .A1(n_41), .A2(n_19), .B1(n_9), .B2(n_11), .C1(n_13), .C2(n_14), .Y(n_43) );
INVx1_ASAP7_75t_L g44 ( .A(n_42), .Y(n_44) );
AOI22xp33_ASAP7_75t_L g45 ( .A1(n_44), .A2(n_19), .B1(n_43), .B2(n_5), .Y(n_45) );
endmodule