module fake_ibex_1420_n_755 (n_85, n_128, n_84, n_64, n_3, n_73, n_65, n_103, n_95, n_55, n_130, n_63, n_98, n_129, n_29, n_106, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_120, n_93, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_88, n_133, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_22, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_105, n_126, n_1, n_111, n_25, n_36, n_104, n_41, n_45, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_50, n_11, n_92, n_101, n_113, n_96, n_68, n_117, n_79, n_81, n_35, n_132, n_31, n_56, n_23, n_91, n_54, n_19, n_755);

input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_103;
input n_95;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_106;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_120;
input n_93;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_88;
input n_133;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_22;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_105;
input n_126;
input n_1;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_50;
input n_11;
input n_92;
input n_101;
input n_113;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_132;
input n_31;
input n_56;
input n_23;
input n_91;
input n_54;
input n_19;

output n_755;

wire n_151;
wire n_599;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_638;
wire n_398;
wire n_304;
wire n_191;
wire n_593;
wire n_153;
wire n_545;
wire n_583;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_608;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_421;
wire n_738;
wire n_475;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_698;
wire n_187;
wire n_667;
wire n_154;
wire n_682;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_723;
wire n_144;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_561;
wire n_417;
wire n_471;
wire n_739;
wire n_265;
wire n_504;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_210;
wire n_348;
wire n_220;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_147;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_598;
wire n_143;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_732;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_168;
wire n_526;
wire n_155;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_515;
wire n_642;
wire n_150;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_750;
wire n_746;
wire n_136;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_355;
wire n_474;
wire n_636;
wire n_594;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_141;
wire n_487;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_454;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_438;
wire n_689;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_205;
wire n_618;
wire n_488;
wire n_139;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_347;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_262;
wire n_299;
wire n_433;
wire n_439;
wire n_704;
wire n_643;
wire n_137;
wire n_679;
wire n_338;
wire n_173;
wire n_696;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_257;
wire n_718;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_713;
wire n_307;
wire n_192;
wire n_140;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_392;
wire n_206;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_546;
wire n_199;
wire n_592;
wire n_495;
wire n_410;
wire n_308;
wire n_675;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_135;
wire n_520;
wire n_684;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_138;
wire n_650;
wire n_409;
wire n_582;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_332;
wire n_517;
wire n_211;
wire n_744;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_415;
wire n_597;
wire n_288;
wire n_285;
wire n_247;
wire n_320;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_148;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_616;
wire n_217;
wire n_324;
wire n_391;
wire n_537;
wire n_728;
wire n_670;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_752;
wire n_668;
wire n_266;
wire n_294;
wire n_485;
wire n_284;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_693;
wire n_311;
wire n_661;
wire n_406;
wire n_606;
wire n_737;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_149;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_687;
wire n_159;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_751;
wire n_160;
wire n_657;
wire n_184;
wire n_492;
wire n_649;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_559;
wire n_425;

INVx2_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_76),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_50),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_32),
.B(n_38),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_68),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_81),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_108),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_14),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_37),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_12),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_29),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_103),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_15),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_35),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_82),
.Y(n_149)
);

INVxp33_ASAP7_75t_SL g150 ( 
.A(n_70),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_4),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_77),
.Y(n_152)
);

BUFx8_ASAP7_75t_SL g153 ( 
.A(n_31),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_4),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_132),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_109),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_36),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_119),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_67),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_52),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_131),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_14),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_80),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_124),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_60),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_63),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_69),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_112),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_75),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_116),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_110),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_94),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_26),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_71),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_19),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_78),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_62),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_64),
.Y(n_181)
);

NOR2xp67_ASAP7_75t_L g182 ( 
.A(n_8),
.B(n_89),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_65),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_24),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_96),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_91),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_123),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_61),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_55),
.Y(n_189)
);

BUFx2_ASAP7_75t_SL g190 ( 
.A(n_15),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_134),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_66),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_90),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_97),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_114),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_53),
.Y(n_196)
);

INVxp33_ASAP7_75t_SL g197 ( 
.A(n_87),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_28),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_56),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_111),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_85),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_115),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_47),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_42),
.Y(n_204)
);

NOR2xp67_ASAP7_75t_L g205 ( 
.A(n_98),
.B(n_121),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_86),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_104),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_54),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_48),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_74),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_72),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_10),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_57),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_39),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_40),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_88),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_105),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_28),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_17),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_30),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_51),
.Y(n_221)
);

INVx4_ASAP7_75t_R g222 ( 
.A(n_133),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_13),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_43),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_18),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_122),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_106),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_59),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_73),
.Y(n_229)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_19),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_113),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_216),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_144),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_151),
.B(n_0),
.Y(n_234)
);

BUFx12f_ASAP7_75t_L g235 ( 
.A(n_149),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_155),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_145),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_161),
.Y(n_239)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_172),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_153),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_142),
.Y(n_243)
);

INVxp33_ASAP7_75t_SL g244 ( 
.A(n_147),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_146),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_245)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_136),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_162),
.Y(n_247)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_230),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

AOI22x1_ASAP7_75t_SL g250 ( 
.A1(n_184),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_218),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_161),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_153),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_230),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_230),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_135),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_135),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_148),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_168),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_164),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_177),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_146),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_163),
.A2(n_11),
.B1(n_16),
.B2(n_17),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_148),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_163),
.A2(n_16),
.B1(n_18),
.B2(n_20),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_139),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_173),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_175),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_140),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_152),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_154),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_173),
.B(n_21),
.Y(n_272)
);

AND2x4_ASAP7_75t_L g273 ( 
.A(n_180),
.B(n_21),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_180),
.B(n_186),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_186),
.B(n_22),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_176),
.B(n_23),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_194),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_191),
.Y(n_278)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_161),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_165),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_203),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_203),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_156),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_158),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_213),
.B(n_25),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_159),
.B(n_27),
.Y(n_286)
);

BUFx8_ASAP7_75t_L g287 ( 
.A(n_218),
.Y(n_287)
);

AND2x6_ASAP7_75t_L g288 ( 
.A(n_166),
.B(n_167),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_218),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_165),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_170),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_203),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_171),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_174),
.Y(n_294)
);

AND2x6_ASAP7_75t_L g295 ( 
.A(n_178),
.B(n_33),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_203),
.Y(n_296)
);

INVx5_ASAP7_75t_L g297 ( 
.A(n_222),
.Y(n_297)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_295),
.Y(n_298)
);

BUFx6f_ASAP7_75t_SL g299 ( 
.A(n_273),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_273),
.B(n_179),
.Y(n_300)
);

OAI22xp33_ASAP7_75t_L g301 ( 
.A1(n_245),
.A2(n_198),
.B1(n_212),
.B2(n_219),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_242),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_242),
.Y(n_303)
);

NAND2xp33_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_141),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_295),
.A2(n_197),
.B1(n_150),
.B2(n_228),
.Y(n_305)
);

BUFx6f_ASAP7_75t_SL g306 ( 
.A(n_232),
.Y(n_306)
);

OR2x6_ASAP7_75t_L g307 ( 
.A(n_241),
.B(n_190),
.Y(n_307)
);

BUFx6f_ASAP7_75t_SL g308 ( 
.A(n_294),
.Y(n_308)
);

OR2x6_ASAP7_75t_L g309 ( 
.A(n_263),
.B(n_182),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_254),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_255),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_266),
.B(n_181),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_239),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_269),
.B(n_183),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_236),
.B(n_223),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_247),
.Y(n_316)
);

AND3x2_ASAP7_75t_L g317 ( 
.A(n_236),
.B(n_138),
.C(n_229),
.Y(n_317)
);

INVx11_ASAP7_75t_L g318 ( 
.A(n_235),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_240),
.Y(n_319)
);

AND3x2_ASAP7_75t_L g320 ( 
.A(n_234),
.B(n_138),
.C(n_207),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_260),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_246),
.B(n_185),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_239),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_239),
.Y(n_324)
);

INVx8_ASAP7_75t_L g325 ( 
.A(n_297),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_268),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_246),
.B(n_225),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_287),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_287),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_274),
.B(n_143),
.Y(n_330)
);

INVx5_ASAP7_75t_L g331 ( 
.A(n_248),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g332 ( 
.A1(n_295),
.A2(n_202),
.B1(n_187),
.B2(n_226),
.Y(n_332)
);

AND2x6_ASAP7_75t_L g333 ( 
.A(n_275),
.B(n_188),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_270),
.B(n_189),
.Y(n_334)
);

INVx5_ASAP7_75t_L g335 ( 
.A(n_248),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_271),
.B(n_291),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_L g337 ( 
.A1(n_295),
.A2(n_204),
.B1(n_192),
.B2(n_224),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_256),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_R g339 ( 
.A(n_253),
.B(n_193),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_237),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_237),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_259),
.Y(n_342)
);

INVx4_ASAP7_75t_SL g343 ( 
.A(n_288),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_283),
.B(n_196),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_257),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_258),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_264),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_264),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_267),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_267),
.Y(n_350)
);

AND3x2_ASAP7_75t_L g351 ( 
.A(n_250),
.B(n_214),
.C(n_200),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_278),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_278),
.Y(n_353)
);

BUFx10_ASAP7_75t_L g354 ( 
.A(n_276),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_249),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_272),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_284),
.B(n_206),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_293),
.B(n_244),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_293),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g360 ( 
.A(n_243),
.B(n_210),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_286),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_252),
.Y(n_362)
);

NAND2xp33_ASAP7_75t_R g363 ( 
.A(n_277),
.B(n_157),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_252),
.Y(n_364)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_251),
.Y(n_365)
);

NAND2xp33_ASAP7_75t_L g366 ( 
.A(n_288),
.B(n_160),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_L g367 ( 
.A1(n_288),
.A2(n_215),
.B1(n_211),
.B2(n_221),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_252),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_285),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_285),
.A2(n_231),
.B1(n_227),
.B2(n_208),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_281),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_281),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_361),
.B(n_356),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_339),
.Y(n_374)
);

OR2x6_ASAP7_75t_L g375 ( 
.A(n_307),
.B(n_233),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_321),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_358),
.A2(n_227),
.B1(n_208),
.B2(n_231),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_319),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_340),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_358),
.A2(n_217),
.B1(n_262),
.B2(n_265),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_330),
.B(n_169),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_327),
.B(n_369),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_L g383 ( 
.A(n_326),
.B(n_280),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_340),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_315),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_341),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_369),
.B(n_137),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_341),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_339),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_359),
.Y(n_390)
);

OAI22x1_ASAP7_75t_SL g391 ( 
.A1(n_316),
.A2(n_253),
.B1(n_290),
.B2(n_217),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g392 ( 
.A1(n_333),
.A2(n_261),
.B1(n_238),
.B2(n_289),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_336),
.B(n_322),
.Y(n_393)
);

NAND2xp33_ASAP7_75t_L g394 ( 
.A(n_332),
.B(n_337),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_365),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_355),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_338),
.Y(n_397)
);

INVx4_ASAP7_75t_L g398 ( 
.A(n_325),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_333),
.A2(n_209),
.B1(n_199),
.B2(n_201),
.Y(n_399)
);

NAND2xp33_ASAP7_75t_L g400 ( 
.A(n_332),
.B(n_195),
.Y(n_400)
);

OR2x6_ASAP7_75t_L g401 ( 
.A(n_307),
.B(n_205),
.Y(n_401)
);

NAND2x1p5_ASAP7_75t_L g402 ( 
.A(n_328),
.B(n_279),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_308),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_347),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_R g405 ( 
.A(n_363),
.B(n_342),
.Y(n_405)
);

A2O1A1Ixp33_ASAP7_75t_L g406 ( 
.A1(n_344),
.A2(n_296),
.B(n_292),
.C(n_282),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_318),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_348),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_337),
.B(n_279),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_329),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_305),
.B(n_281),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_308),
.Y(n_412)
);

NOR2xp67_ASAP7_75t_L g413 ( 
.A(n_360),
.B(n_30),
.Y(n_413)
);

INVx2_ASAP7_75t_SL g414 ( 
.A(n_354),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_300),
.B(n_296),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_300),
.B(n_354),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_333),
.B(n_312),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_299),
.B(n_296),
.Y(n_418)
);

AND2x2_ASAP7_75t_SL g419 ( 
.A(n_304),
.B(n_367),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_L g420 ( 
.A1(n_333),
.A2(n_344),
.B1(n_349),
.B2(n_350),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_307),
.B(n_31),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_345),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_299),
.B(n_34),
.Y(n_423)
);

INVx2_ASAP7_75t_SL g424 ( 
.A(n_320),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_346),
.Y(n_425)
);

NOR2x1p5_ASAP7_75t_L g426 ( 
.A(n_306),
.B(n_41),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_314),
.B(n_44),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_334),
.B(n_45),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_352),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_334),
.B(n_46),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_353),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_370),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_367),
.B(n_49),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_L g434 ( 
.A1(n_357),
.A2(n_310),
.B1(n_302),
.B2(n_303),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_373),
.A2(n_420),
.B1(n_419),
.B2(n_376),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_373),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_382),
.B(n_393),
.Y(n_437)
);

O2A1O1Ixp5_ASAP7_75t_L g438 ( 
.A1(n_411),
.A2(n_311),
.B(n_302),
.C(n_303),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_382),
.B(n_320),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_376),
.B(n_301),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_387),
.B(n_416),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_387),
.B(n_317),
.Y(n_442)
);

NAND3xp33_ASAP7_75t_L g443 ( 
.A(n_394),
.B(n_363),
.C(n_366),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_383),
.A2(n_301),
.B1(n_309),
.B2(n_325),
.Y(n_444)
);

CKINVDCx10_ASAP7_75t_R g445 ( 
.A(n_375),
.Y(n_445)
);

O2A1O1Ixp33_ASAP7_75t_L g446 ( 
.A1(n_411),
.A2(n_309),
.B(n_311),
.C(n_310),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_378),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_414),
.B(n_385),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_396),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_398),
.B(n_343),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_417),
.A2(n_331),
.B(n_335),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_390),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_397),
.Y(n_453)
);

AOI21x1_ASAP7_75t_L g454 ( 
.A1(n_409),
.A2(n_372),
.B(n_371),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_L g455 ( 
.A1(n_419),
.A2(n_351),
.B1(n_343),
.B2(n_335),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_420),
.A2(n_331),
.B1(n_335),
.B2(n_351),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_398),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_407),
.B(n_313),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_392),
.A2(n_368),
.B1(n_364),
.B2(n_362),
.Y(n_459)
);

NAND2xp33_ASAP7_75t_SL g460 ( 
.A(n_405),
.B(n_362),
.Y(n_460)
);

BUFx8_ASAP7_75t_SL g461 ( 
.A(n_374),
.Y(n_461)
);

BUFx8_ASAP7_75t_L g462 ( 
.A(n_421),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_392),
.A2(n_324),
.B1(n_323),
.B2(n_313),
.Y(n_463)
);

OR2x6_ASAP7_75t_SL g464 ( 
.A(n_389),
.B(n_58),
.Y(n_464)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_410),
.Y(n_465)
);

OA22x2_ASAP7_75t_L g466 ( 
.A1(n_380),
.A2(n_375),
.B1(n_432),
.B2(n_424),
.Y(n_466)
);

AOI21x1_ASAP7_75t_L g467 ( 
.A1(n_427),
.A2(n_79),
.B(n_83),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_399),
.B(n_84),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_413),
.B(n_381),
.Y(n_469)
);

A2O1A1Ixp33_ASAP7_75t_L g470 ( 
.A1(n_422),
.A2(n_92),
.B(n_93),
.C(n_95),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_425),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_434),
.A2(n_100),
.B(n_101),
.Y(n_472)
);

OR2x6_ASAP7_75t_L g473 ( 
.A(n_375),
.B(n_102),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_429),
.B(n_431),
.Y(n_474)
);

NAND3xp33_ASAP7_75t_SL g475 ( 
.A(n_405),
.B(n_117),
.C(n_118),
.Y(n_475)
);

O2A1O1Ixp33_ASAP7_75t_L g476 ( 
.A1(n_400),
.A2(n_130),
.B(n_125),
.C(n_127),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_434),
.A2(n_120),
.B1(n_129),
.B2(n_404),
.Y(n_477)
);

AND2x2_ASAP7_75t_SL g478 ( 
.A(n_403),
.B(n_391),
.Y(n_478)
);

A2O1A1Ixp33_ASAP7_75t_L g479 ( 
.A1(n_415),
.A2(n_408),
.B(n_428),
.C(n_430),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_403),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_379),
.A2(n_388),
.B1(n_384),
.B2(n_386),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_401),
.B(n_412),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_412),
.A2(n_402),
.B1(n_426),
.B2(n_395),
.Y(n_483)
);

OAI21xp33_ASAP7_75t_L g484 ( 
.A1(n_423),
.A2(n_418),
.B(n_433),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_406),
.B(n_373),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_373),
.Y(n_486)
);

NAND3xp33_ASAP7_75t_L g487 ( 
.A(n_387),
.B(n_305),
.C(n_382),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_376),
.B(n_414),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_373),
.B(n_382),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_373),
.B(n_382),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_489),
.A2(n_490),
.B(n_437),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_436),
.Y(n_492)
);

INVx3_ASAP7_75t_SL g493 ( 
.A(n_478),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_479),
.A2(n_474),
.B(n_441),
.Y(n_494)
);

OR2x6_ASAP7_75t_SL g495 ( 
.A(n_445),
.B(n_483),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_457),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_486),
.B(n_440),
.Y(n_497)
);

AOI21xp33_ASAP7_75t_L g498 ( 
.A1(n_448),
.A2(n_488),
.B(n_442),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_480),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_447),
.B(n_452),
.Y(n_500)
);

AOI221x1_ASAP7_75t_L g501 ( 
.A1(n_443),
.A2(n_477),
.B1(n_484),
.B2(n_475),
.C(n_470),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_453),
.B(n_471),
.Y(n_502)
);

OAI21x1_ASAP7_75t_L g503 ( 
.A1(n_459),
.A2(n_463),
.B(n_451),
.Y(n_503)
);

AO22x2_ASAP7_75t_L g504 ( 
.A1(n_466),
.A2(n_445),
.B1(n_473),
.B2(n_439),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_461),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_444),
.B(n_455),
.Y(n_506)
);

INVxp33_ASAP7_75t_L g507 ( 
.A(n_482),
.Y(n_507)
);

AO32x2_ASAP7_75t_L g508 ( 
.A1(n_481),
.A2(n_456),
.A3(n_465),
.B1(n_464),
.B2(n_460),
.Y(n_508)
);

NOR2x1_ASAP7_75t_R g509 ( 
.A(n_465),
.B(n_450),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_462),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_458),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_489),
.A2(n_490),
.B(n_304),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_480),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_449),
.Y(n_514)
);

OR2x2_ASAP7_75t_L g515 ( 
.A(n_489),
.B(n_376),
.Y(n_515)
);

A2O1A1Ixp33_ASAP7_75t_L g516 ( 
.A1(n_437),
.A2(n_446),
.B(n_487),
.C(n_489),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_437),
.B(n_489),
.Y(n_517)
);

INVx6_ASAP7_75t_L g518 ( 
.A(n_465),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_454),
.A2(n_438),
.B(n_467),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_436),
.B(n_486),
.Y(n_520)
);

INVx2_ASAP7_75t_SL g521 ( 
.A(n_480),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_490),
.A2(n_489),
.B1(n_437),
.B2(n_486),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_486),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_489),
.A2(n_490),
.B(n_304),
.Y(n_524)
);

AO31x2_ASAP7_75t_L g525 ( 
.A1(n_435),
.A2(n_477),
.A3(n_470),
.B(n_485),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_440),
.B(n_376),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_437),
.B(n_489),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_SL g528 ( 
.A1(n_473),
.A2(n_298),
.B(n_477),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_437),
.B(n_489),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_436),
.Y(n_530)
);

BUFx12f_ASAP7_75t_L g531 ( 
.A(n_478),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_457),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_437),
.B(n_489),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_436),
.B(n_486),
.Y(n_534)
);

AO31x2_ASAP7_75t_L g535 ( 
.A1(n_435),
.A2(n_477),
.A3(n_470),
.B(n_485),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_437),
.B(n_489),
.Y(n_536)
);

AO32x2_ASAP7_75t_L g537 ( 
.A1(n_435),
.A2(n_477),
.A3(n_483),
.B1(n_481),
.B2(n_463),
.Y(n_537)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_489),
.B(n_376),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_436),
.Y(n_539)
);

O2A1O1Ixp5_ASAP7_75t_L g540 ( 
.A1(n_469),
.A2(n_411),
.B(n_468),
.C(n_460),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_486),
.B(n_373),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_436),
.B(n_486),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_440),
.B(n_376),
.Y(n_543)
);

NOR3xp33_ASAP7_75t_L g544 ( 
.A(n_489),
.B(n_490),
.C(n_437),
.Y(n_544)
);

AO21x1_ASAP7_75t_L g545 ( 
.A1(n_472),
.A2(n_476),
.B(n_477),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_436),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_486),
.B(n_373),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_437),
.B(n_489),
.Y(n_548)
);

INVx3_ASAP7_75t_SL g549 ( 
.A(n_478),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_436),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_437),
.B(n_489),
.Y(n_551)
);

AO32x2_ASAP7_75t_L g552 ( 
.A1(n_435),
.A2(n_477),
.A3(n_483),
.B1(n_481),
.B2(n_463),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_436),
.Y(n_553)
);

CKINVDCx6p67_ASAP7_75t_R g554 ( 
.A(n_445),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_490),
.A2(n_489),
.B1(n_437),
.B2(n_486),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_437),
.B(n_489),
.Y(n_556)
);

INVx5_ASAP7_75t_L g557 ( 
.A(n_457),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_437),
.A2(n_376),
.B1(n_377),
.B2(n_290),
.Y(n_558)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_457),
.Y(n_559)
);

OA21x2_ASAP7_75t_L g560 ( 
.A1(n_503),
.A2(n_501),
.B(n_519),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_522),
.A2(n_555),
.B1(n_536),
.B2(n_517),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_492),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_514),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_530),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_515),
.B(n_538),
.Y(n_565)
);

BUFx4_ASAP7_75t_R g566 ( 
.A(n_499),
.Y(n_566)
);

OA21x2_ASAP7_75t_L g567 ( 
.A1(n_545),
.A2(n_494),
.B(n_540),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_539),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_557),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_544),
.B(n_527),
.Y(n_570)
);

AO21x2_ASAP7_75t_L g571 ( 
.A1(n_528),
.A2(n_524),
.B(n_512),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_557),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_491),
.B(n_529),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_533),
.B(n_548),
.Y(n_574)
);

AO21x1_ASAP7_75t_L g575 ( 
.A1(n_511),
.A2(n_506),
.B(n_497),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g576 ( 
.A(n_551),
.B(n_556),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_557),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_546),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_520),
.B(n_542),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_518),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_526),
.B(n_543),
.Y(n_581)
);

AO31x2_ASAP7_75t_L g582 ( 
.A1(n_550),
.A2(n_553),
.A3(n_535),
.B(n_525),
.Y(n_582)
);

NAND3xp33_ASAP7_75t_L g583 ( 
.A(n_498),
.B(n_500),
.C(n_502),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_520),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_534),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_496),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_534),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_541),
.B(n_547),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_542),
.B(n_559),
.Y(n_589)
);

OA21x2_ASAP7_75t_L g590 ( 
.A1(n_537),
.A2(n_552),
.B(n_508),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_523),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_558),
.B(n_513),
.Y(n_592)
);

OR2x2_ASAP7_75t_L g593 ( 
.A(n_521),
.B(n_554),
.Y(n_593)
);

OR2x2_ASAP7_75t_L g594 ( 
.A(n_510),
.B(n_507),
.Y(n_594)
);

CKINVDCx6p67_ASAP7_75t_R g595 ( 
.A(n_505),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_L g596 ( 
.A1(n_552),
.A2(n_508),
.B(n_504),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_504),
.B(n_532),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_518),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_509),
.Y(n_599)
);

OAI21x1_ASAP7_75t_L g600 ( 
.A1(n_508),
.A2(n_495),
.B(n_493),
.Y(n_600)
);

BUFx2_ASAP7_75t_R g601 ( 
.A(n_549),
.Y(n_601)
);

BUFx8_ASAP7_75t_SL g602 ( 
.A(n_531),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_492),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_492),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_557),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_517),
.B(n_527),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_557),
.Y(n_607)
);

OR2x6_ASAP7_75t_L g608 ( 
.A(n_504),
.B(n_473),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_491),
.B(n_544),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_515),
.B(n_538),
.Y(n_610)
);

CKINVDCx6p67_ASAP7_75t_R g611 ( 
.A(n_554),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_R g612 ( 
.A(n_510),
.B(n_290),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_491),
.B(n_544),
.Y(n_613)
);

AO31x2_ASAP7_75t_L g614 ( 
.A1(n_545),
.A2(n_501),
.A3(n_516),
.B(n_494),
.Y(n_614)
);

INVx1_ASAP7_75t_SL g615 ( 
.A(n_513),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_522),
.A2(n_555),
.B1(n_473),
.B2(n_490),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_608),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_609),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_616),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g620 ( 
.A(n_576),
.B(n_574),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_605),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_573),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_566),
.Y(n_623)
);

INVx4_ASAP7_75t_L g624 ( 
.A(n_566),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_613),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_613),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_561),
.B(n_570),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_582),
.Y(n_628)
);

INVx4_ASAP7_75t_L g629 ( 
.A(n_608),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_582),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_606),
.B(n_574),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_597),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_569),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_569),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_563),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_570),
.B(n_606),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_562),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_564),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_568),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_578),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_603),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_565),
.B(n_610),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_560),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_604),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_596),
.B(n_581),
.Y(n_645)
);

OAI22xp33_ASAP7_75t_L g646 ( 
.A1(n_592),
.A2(n_581),
.B1(n_588),
.B2(n_591),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_572),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_622),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_621),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_636),
.B(n_590),
.Y(n_650)
);

NAND4xp25_ASAP7_75t_L g651 ( 
.A(n_631),
.B(n_583),
.C(n_585),
.D(n_587),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_622),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_618),
.Y(n_653)
);

OAI221xp5_ASAP7_75t_L g654 ( 
.A1(n_627),
.A2(n_583),
.B1(n_599),
.B2(n_584),
.C(n_615),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_636),
.B(n_567),
.Y(n_655)
);

OAI221xp5_ASAP7_75t_L g656 ( 
.A1(n_620),
.A2(n_615),
.B1(n_594),
.B2(n_593),
.C(n_580),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_643),
.Y(n_657)
);

OR2x2_ASAP7_75t_L g658 ( 
.A(n_645),
.B(n_600),
.Y(n_658)
);

NOR2x1_ASAP7_75t_SL g659 ( 
.A(n_624),
.B(n_586),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_635),
.B(n_614),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_621),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_625),
.B(n_614),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_626),
.B(n_614),
.Y(n_663)
);

INVx5_ASAP7_75t_L g664 ( 
.A(n_624),
.Y(n_664)
);

OAI211xp5_ASAP7_75t_L g665 ( 
.A1(n_617),
.A2(n_612),
.B(n_598),
.C(n_607),
.Y(n_665)
);

OR2x2_ASAP7_75t_L g666 ( 
.A(n_645),
.B(n_575),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_SL g667 ( 
.A1(n_624),
.A2(n_589),
.B(n_579),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_619),
.B(n_571),
.Y(n_668)
);

OR2x6_ASAP7_75t_L g669 ( 
.A(n_629),
.B(n_577),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_621),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_642),
.B(n_607),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_650),
.B(n_628),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_657),
.Y(n_673)
);

OR2x2_ASAP7_75t_L g674 ( 
.A(n_650),
.B(n_632),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_666),
.B(n_637),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_655),
.B(n_630),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_662),
.B(n_663),
.Y(n_677)
);

HB1xp67_ASAP7_75t_SL g678 ( 
.A(n_649),
.Y(n_678)
);

INVxp33_ASAP7_75t_L g679 ( 
.A(n_671),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_653),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_660),
.B(n_629),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_660),
.B(n_629),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_677),
.B(n_648),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_677),
.B(n_668),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_681),
.B(n_682),
.Y(n_685)
);

AND2x2_ASAP7_75t_SL g686 ( 
.A(n_681),
.B(n_617),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_673),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_678),
.Y(n_688)
);

AND2x4_ASAP7_75t_L g689 ( 
.A(n_681),
.B(n_652),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_675),
.B(n_652),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_680),
.Y(n_691)
);

OR2x6_ASAP7_75t_L g692 ( 
.A(n_682),
.B(n_667),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_674),
.B(n_658),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_682),
.B(n_664),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_672),
.B(n_668),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_672),
.B(n_662),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_680),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_684),
.B(n_696),
.Y(n_698)
);

INVxp67_ASAP7_75t_L g699 ( 
.A(n_693),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_687),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_696),
.B(n_695),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_695),
.B(n_676),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_683),
.B(n_656),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_691),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_687),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_684),
.B(n_676),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_697),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_688),
.B(n_664),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_703),
.A2(n_689),
.B1(n_686),
.B2(n_692),
.Y(n_709)
);

INVxp67_ASAP7_75t_L g710 ( 
.A(n_703),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_699),
.B(n_611),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_708),
.A2(n_692),
.B(n_686),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_708),
.Y(n_713)
);

OAI32xp33_ASAP7_75t_L g714 ( 
.A1(n_701),
.A2(n_649),
.A3(n_661),
.B1(n_670),
.B2(n_679),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_702),
.B(n_674),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_698),
.B(n_690),
.Y(n_716)
);

NAND2x1p5_ASAP7_75t_L g717 ( 
.A(n_700),
.B(n_649),
.Y(n_717)
);

O2A1O1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_710),
.A2(n_646),
.B(n_654),
.C(n_651),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_SL g719 ( 
.A1(n_712),
.A2(n_685),
.B1(n_694),
.B2(n_692),
.Y(n_719)
);

AOI21xp33_ASAP7_75t_L g720 ( 
.A1(n_711),
.A2(n_665),
.B(n_642),
.Y(n_720)
);

AOI32xp33_ASAP7_75t_L g721 ( 
.A1(n_713),
.A2(n_685),
.A3(n_694),
.B1(n_706),
.B2(n_689),
.Y(n_721)
);

OAI22xp33_ASAP7_75t_L g722 ( 
.A1(n_719),
.A2(n_709),
.B1(n_692),
.B2(n_717),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_720),
.A2(n_689),
.B1(n_716),
.B2(n_704),
.Y(n_723)
);

OAI211xp5_ASAP7_75t_SL g724 ( 
.A1(n_721),
.A2(n_667),
.B(n_715),
.C(n_623),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_723),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_722),
.B(n_595),
.Y(n_726)
);

NOR2xp67_ASAP7_75t_L g727 ( 
.A(n_726),
.B(n_724),
.Y(n_727)
);

OAI211xp5_ASAP7_75t_SL g728 ( 
.A1(n_725),
.A2(n_718),
.B(n_612),
.C(n_601),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_728),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_727),
.A2(n_685),
.B1(n_601),
.B2(n_694),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_730),
.Y(n_731)
);

XNOR2x1_ASAP7_75t_L g732 ( 
.A(n_729),
.B(n_602),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_731),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_732),
.B(n_705),
.Y(n_734)
);

OAI21x1_ASAP7_75t_SL g735 ( 
.A1(n_732),
.A2(n_602),
.B(n_659),
.Y(n_735)
);

XNOR2xp5_ASAP7_75t_L g736 ( 
.A(n_733),
.B(n_651),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_734),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_735),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_733),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_734),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_740),
.Y(n_741)
);

NOR2xp67_ASAP7_75t_L g742 ( 
.A(n_738),
.B(n_633),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_739),
.A2(n_714),
.B(n_634),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_740),
.A2(n_669),
.B1(n_700),
.B2(n_664),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_737),
.A2(n_669),
.B1(n_664),
.B2(n_633),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_736),
.B(n_707),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_740),
.Y(n_747)
);

AOI221xp5_ASAP7_75t_L g748 ( 
.A1(n_741),
.A2(n_640),
.B1(n_641),
.B2(n_644),
.C(n_638),
.Y(n_748)
);

OA21x2_ASAP7_75t_L g749 ( 
.A1(n_747),
.A2(n_639),
.B(n_640),
.Y(n_749)
);

OAI21xp5_ASAP7_75t_SL g750 ( 
.A1(n_746),
.A2(n_745),
.B(n_743),
.Y(n_750)
);

OAI21x1_ASAP7_75t_SL g751 ( 
.A1(n_742),
.A2(n_659),
.B(n_647),
.Y(n_751)
);

OAI21xp5_ASAP7_75t_L g752 ( 
.A1(n_750),
.A2(n_744),
.B(n_633),
.Y(n_752)
);

OAI21xp5_ASAP7_75t_L g753 ( 
.A1(n_749),
.A2(n_634),
.B(n_633),
.Y(n_753)
);

BUFx24_ASAP7_75t_SL g754 ( 
.A(n_752),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_754),
.A2(n_751),
.B1(n_753),
.B2(n_748),
.Y(n_755)
);


endmodule