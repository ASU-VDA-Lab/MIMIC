module fake_jpeg_3689_n_187 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_187);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_3),
.B(n_0),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_44),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_31),
.Y(n_51)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_20),
.Y(n_39)
);

CKINVDCx6p67_ASAP7_75t_R g70 ( 
.A(n_39),
.Y(n_70)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_1),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_43),
.B(n_2),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_48),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_18),
.B(n_15),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_49),
.Y(n_54)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_28),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_51),
.B(n_58),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_48),
.A2(n_31),
.B1(n_32),
.B2(n_30),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_56),
.B1(n_62),
.B2(n_64),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_31),
.B1(n_32),
.B2(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_19),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_40),
.B(n_18),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_73),
.Y(n_94)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_36),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_17),
.C(n_26),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_24),
.C(n_33),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_27),
.B1(n_23),
.B2(n_17),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_67),
.B(n_71),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_43),
.B(n_34),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_34),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

AND2x6_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_12),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_84),
.Y(n_102)
);

HAxp5_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_19),
.CON(n_78),
.SN(n_78)
);

NOR2x1_ASAP7_75t_R g115 ( 
.A(n_78),
.B(n_99),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_68),
.A2(n_24),
.B1(n_33),
.B2(n_23),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_88),
.B1(n_89),
.B2(n_74),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_91),
.Y(n_104)
);

INVxp33_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_58),
.Y(n_84)
);

AND2x6_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_8),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_95),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_55),
.A2(n_24),
.B1(n_23),
.B2(n_5),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_55),
.A2(n_23),
.B1(n_4),
.B2(n_5),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_2),
.C(n_4),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_55),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_93),
.B(n_70),
.Y(n_101)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_98),
.Y(n_118)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_70),
.B(n_51),
.Y(n_99)
);

BUFx4f_ASAP7_75t_SL g100 ( 
.A(n_97),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_100),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g124 ( 
.A1(n_101),
.A2(n_79),
.B(n_81),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_94),
.B(n_65),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_103),
.B(n_113),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_83),
.Y(n_123)
);

OAI32xp33_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_70),
.A3(n_54),
.B1(n_53),
.B2(n_65),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_81),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_78),
.A2(n_69),
.B(n_65),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_88),
.B1(n_92),
.B2(n_83),
.Y(n_121)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_99),
.A2(n_75),
.B1(n_66),
.B2(n_69),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_112),
.A2(n_66),
.B1(n_81),
.B2(n_61),
.Y(n_130)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_76),
.A2(n_61),
.B(n_66),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_119),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_90),
.B(n_77),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_117),
.B(n_8),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_99),
.A2(n_81),
.B(n_89),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_121),
.A2(n_130),
.B1(n_131),
.B2(n_110),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_127),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_91),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_126),
.B(n_134),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_85),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_108),
.Y(n_132)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_114),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_114),
.B(n_13),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_135),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_61),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_137),
.C(n_115),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_5),
.C(n_6),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_137),
.Y(n_161)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_109),
.C(n_119),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_150),
.C(n_133),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_122),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_151),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_120),
.Y(n_148)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_116),
.C(n_118),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_120),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_154),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_144),
.B(n_125),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_160),
.C(n_161),
.Y(n_163)
);

XNOR2x2_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_146),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_141),
.A2(n_133),
.B1(n_128),
.B2(n_112),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_157),
.A2(n_101),
.B1(n_107),
.B2(n_148),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_136),
.C(n_128),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_138),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_140),
.C(n_142),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_113),
.C(n_106),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_SL g166 ( 
.A1(n_158),
.A2(n_141),
.B(n_130),
.C(n_106),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_166),
.A2(n_168),
.B(n_100),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_169),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_158),
.A2(n_143),
.B1(n_139),
.B2(n_118),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_120),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_156),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_6),
.B1(n_7),
.B2(n_176),
.Y(n_179)
);

A2O1A1O1Ixp25_ASAP7_75t_L g172 ( 
.A1(n_163),
.A2(n_154),
.B(n_160),
.C(n_153),
.D(n_155),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_172),
.A2(n_175),
.B(n_7),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_173),
.A2(n_176),
.B(n_166),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_170),
.A2(n_111),
.B(n_100),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_174),
.A2(n_166),
.B1(n_165),
.B2(n_100),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_178),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_179),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_180),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_177),
.C(n_7),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_184),
.A2(n_185),
.B(n_181),
.Y(n_186)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_183),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_181),
.Y(n_187)
);


endmodule