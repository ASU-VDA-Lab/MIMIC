module fake_jpeg_28752_n_99 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_99);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_99;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_25),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_0),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_43),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_32),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_62),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_48),
.A2(n_40),
.B1(n_37),
.B2(n_34),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_55),
.A2(n_59),
.B1(n_1),
.B2(n_2),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_58),
.B(n_60),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_49),
.A2(n_41),
.B1(n_38),
.B2(n_33),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_51),
.B(n_44),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_43),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_59),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_61),
.A2(n_42),
.B1(n_39),
.B2(n_43),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_66),
.A2(n_67),
.B1(n_74),
.B2(n_1),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_55),
.A2(n_13),
.B1(n_28),
.B2(n_26),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_72),
.Y(n_77)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_10),
.C(n_21),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_73),
.C(n_7),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_62),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_29),
.C(n_20),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_18),
.B1(n_17),
.B2(n_14),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_84),
.B1(n_8),
.B2(n_77),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_2),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_75),
.B(n_3),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_80),
.A2(n_81),
.B(n_83),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_75),
.B(n_3),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_4),
.B(n_6),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_4),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_65),
.A2(n_11),
.B1(n_7),
.B2(n_8),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_82),
.C(n_86),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_89),
.Y(n_93)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_92),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_94),
.A2(n_91),
.B(n_93),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_95),
.B(n_88),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_87),
.Y(n_99)
);


endmodule