module fake_jpeg_28961_n_50 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_50);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_50;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_44;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_14),
.B(n_15),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_19),
.Y(n_26)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_1),
.C(n_2),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_18),
.A2(n_23),
.B(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_5),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_9),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_20)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_12),
.B1(n_13),
.B2(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_8),
.Y(n_21)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_22),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_9),
.A2(n_3),
.B(n_4),
.C(n_12),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_24),
.A2(n_21),
.B1(n_22),
.B2(n_17),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_18),
.B(n_23),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_24),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_33),
.B1(n_34),
.B2(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_28),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_10),
.B1(n_11),
.B2(n_27),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_10),
.B1(n_11),
.B2(n_27),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_36),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_29),
.C(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_38),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_37),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_42),
.Y(n_43)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_31),
.B1(n_24),
.B2(n_32),
.Y(n_44)
);

AO21x1_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_39),
.B(n_25),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_42),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_45),
.B(n_39),
.Y(n_46)
);

AOI322xp5_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_47),
.A3(n_25),
.B1(n_45),
.B2(n_43),
.C1(n_11),
.C2(n_26),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_43),
.C(n_45),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_26),
.C(n_25),
.Y(n_50)
);


endmodule