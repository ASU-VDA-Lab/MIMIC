module fake_ariane_252_n_1207 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1207);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1207;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_1127;
wire n_1072;
wire n_695;
wire n_913;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_1137;
wire n_646;
wire n_1174;
wire n_197;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_1118;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_183;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_1123;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_1169;
wire n_789;
wire n_788;
wire n_908;
wire n_850;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_205;
wire n_1029;
wire n_341;
wire n_1187;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_760;
wire n_522;
wire n_319;
wire n_591;
wire n_906;
wire n_690;
wire n_416;
wire n_1180;
wire n_969;
wire n_283;
wire n_1109;
wire n_919;
wire n_525;
wire n_187;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_1095;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_819;
wire n_717;
wire n_189;
wire n_286;
wire n_586;
wire n_443;
wire n_952;
wire n_864;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_1154;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1130;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_940;
wire n_756;
wire n_466;
wire n_1016;
wire n_346;
wire n_1138;
wire n_214;
wire n_1149;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_1196;
wire n_607;
wire n_670;
wire n_897;
wire n_956;
wire n_949;
wire n_410;
wire n_1181;
wire n_379;
wire n_515;
wire n_807;
wire n_445;
wire n_1131;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_1177;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_1167;
wire n_1170;
wire n_1151;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_905;
wire n_279;
wire n_958;
wire n_702;
wire n_945;
wire n_790;
wire n_857;
wire n_898;
wire n_207;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_194;
wire n_1064;
wire n_633;
wire n_900;
wire n_1133;
wire n_883;
wire n_338;
wire n_1163;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_186;
wire n_801;
wire n_1184;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_1173;
wire n_311;
wire n_239;
wire n_402;
wire n_1068;
wire n_1052;
wire n_272;
wire n_829;
wire n_1198;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_1018;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_989;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_1125;
wire n_625;
wire n_405;
wire n_557;
wire n_1201;
wire n_1107;
wire n_858;
wire n_242;
wire n_645;
wire n_1185;
wire n_320;
wire n_331;
wire n_309;
wire n_559;
wire n_1134;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_1141;
wire n_350;
wire n_291;
wire n_822;
wire n_1143;
wire n_381;
wire n_344;
wire n_840;
wire n_426;
wire n_481;
wire n_433;
wire n_600;
wire n_721;
wire n_795;
wire n_1053;
wire n_1084;
wire n_398;
wire n_210;
wire n_1090;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_928;
wire n_839;
wire n_1099;
wire n_218;
wire n_1153;
wire n_271;
wire n_507;
wire n_465;
wire n_486;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_1145;
wire n_971;
wire n_240;
wire n_369;
wire n_1192;
wire n_224;
wire n_894;
wire n_787;
wire n_1105;
wire n_547;
wire n_1195;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_1172;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_1160;
wire n_874;
wire n_188;
wire n_323;
wire n_550;
wire n_1023;
wire n_997;
wire n_635;
wire n_707;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_1116;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_1085;
wire n_1152;
wire n_432;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_1197;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_1165;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_920;
wire n_899;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_238;
wire n_365;
wire n_455;
wire n_654;
wire n_429;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_192;
wire n_1128;
wire n_887;
wire n_729;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1122;
wire n_1049;
wire n_1205;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_1132;
wire n_390;
wire n_1156;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_1120;
wire n_440;
wire n_1202;
wire n_627;
wire n_1039;
wire n_1188;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_1150;
wire n_233;
wire n_728;
wire n_957;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_321;
wire n_911;
wire n_221;
wire n_1136;
wire n_361;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_1119;
wire n_734;
wire n_491;
wire n_810;
wire n_181;
wire n_723;
wire n_1142;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_1140;
wire n_570;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_1121;
wire n_490;
wire n_262;
wire n_209;
wire n_743;
wire n_1194;
wire n_907;
wire n_225;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_1019;
wire n_735;
wire n_575;
wire n_546;
wire n_464;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_1159;
wire n_910;
wire n_290;
wire n_527;
wire n_772;
wire n_741;
wire n_847;
wire n_747;
wire n_939;
wire n_1135;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_217;
wire n_1114;
wire n_676;
wire n_708;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_1038;
wire n_572;
wire n_343;
wire n_1199;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_1108;
wire n_355;
wire n_851;
wire n_212;
wire n_444;
wire n_609;
wire n_1164;
wire n_1043;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_1193;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_1179;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_1081;
wire n_1166;
wire n_182;
wire n_696;
wire n_1040;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_1158;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_872;
wire n_774;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_1168;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_1157;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_252;
wire n_629;
wire n_664;
wire n_215;
wire n_1075;
wire n_454;
wire n_992;
wire n_966;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_1182;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_692;
wire n_216;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_991;
wire n_834;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_179;
wire n_812;
wire n_1126;
wire n_395;
wire n_621;
wire n_1178;
wire n_195;
wire n_606;
wire n_951;
wire n_1026;
wire n_938;
wire n_213;
wire n_862;
wire n_895;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_1206;
wire n_203;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1146;
wire n_1100;
wire n_1171;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_1203;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_998;
wire n_999;
wire n_967;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1175;
wire n_1044;
wire n_1148;
wire n_751;
wire n_1027;
wire n_615;
wire n_1070;
wire n_204;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1139;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_1101;
wire n_975;
wire n_1102;
wire n_1129;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_1189;
wire n_1124;
wire n_250;
wire n_932;
wire n_1183;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_944;
wire n_749;
wire n_1204;
wire n_994;
wire n_289;
wire n_548;
wire n_815;
wire n_542;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_184;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_1161;
wire n_431;
wire n_1176;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1155;
wire n_1191;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_191;
wire n_489;
wire n_480;
wire n_1011;
wire n_642;
wire n_211;
wire n_978;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_1147;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g179 ( 
.A(n_70),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_101),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_105),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_81),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_99),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_111),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_127),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_67),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_78),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_177),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_74),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_59),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_141),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_6),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_29),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g195 ( 
.A(n_145),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_21),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_17),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_16),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_77),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_62),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_48),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_16),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_154),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_158),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_11),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_117),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_122),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_115),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_75),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_149),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_162),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_28),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_68),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_125),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_131),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_71),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_118),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_172),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_47),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_9),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_169),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_175),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_93),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_116),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_129),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_43),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_53),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_159),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_144),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_164),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_124),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_90),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_4),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_7),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_182),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_182),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_188),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_196),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_199),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_188),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_206),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_234),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_234),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_192),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_235),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_194),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_194),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_194),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_183),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_194),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_203),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_203),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_183),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_214),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_222),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_179),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_236),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_223),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_180),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_181),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_184),
.Y(n_265)
);

BUFx10_ASAP7_75t_L g266 ( 
.A(n_186),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_244),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_262),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_250),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_240),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_241),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_265),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_237),
.Y(n_277)
);

INVxp67_ASAP7_75t_SL g278 ( 
.A(n_260),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_237),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_255),
.Y(n_281)
);

INVxp67_ASAP7_75t_SL g282 ( 
.A(n_256),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_247),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_238),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_248),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_263),
.Y(n_286)
);

INVxp67_ASAP7_75t_SL g287 ( 
.A(n_258),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_238),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_246),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_239),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_252),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_252),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_257),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_257),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_239),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_259),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_264),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_264),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_245),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_242),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_266),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_259),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_266),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_254),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_242),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_240),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_240),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_244),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_244),
.Y(n_309)
);

BUFx5_ASAP7_75t_L g310 ( 
.A(n_249),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_261),
.Y(n_311)
);

BUFx10_ASAP7_75t_L g312 ( 
.A(n_264),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_255),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_244),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_269),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_272),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_273),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_311),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_274),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_268),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_267),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_299),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_271),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_279),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_278),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_283),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_283),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_285),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_310),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_276),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_306),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_277),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_268),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_286),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_304),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_270),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_307),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_270),
.Y(n_338)
);

INVxp33_ASAP7_75t_L g339 ( 
.A(n_296),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_280),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_312),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_288),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_290),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_275),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_295),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_304),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_310),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_284),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_287),
.Y(n_349)
);

INVxp33_ASAP7_75t_SL g350 ( 
.A(n_284),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_310),
.Y(n_351)
);

INVxp33_ASAP7_75t_SL g352 ( 
.A(n_300),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_275),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_312),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_300),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_315),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_321),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_330),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_322),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_330),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_321),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_318),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_335),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_332),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_323),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_323),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_332),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_328),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_328),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_348),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_318),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_340),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_355),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_325),
.B(n_302),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_340),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_326),
.Y(n_376)
);

NOR2xp67_ASAP7_75t_L g377 ( 
.A(n_341),
.B(n_314),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_348),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_327),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_327),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_342),
.Y(n_381)
);

NOR2xp67_ASAP7_75t_L g382 ( 
.A(n_341),
.B(n_308),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_324),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_320),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_342),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_345),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_324),
.Y(n_387)
);

CKINVDCx14_ASAP7_75t_R g388 ( 
.A(n_345),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_350),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_316),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_343),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_352),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_333),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_354),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_354),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_346),
.Y(n_396)
);

BUFx8_ASAP7_75t_L g397 ( 
.A(n_384),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_368),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_362),
.B(n_371),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_373),
.A2(n_291),
.B1(n_293),
.B2(n_292),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_369),
.B(n_334),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_376),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_383),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_386),
.B(n_339),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_376),
.Y(n_405)
);

NAND2xp33_ASAP7_75t_L g406 ( 
.A(n_394),
.B(n_329),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_379),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_379),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_387),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_390),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_356),
.Y(n_411)
);

AND2x6_ASAP7_75t_L g412 ( 
.A(n_357),
.B(n_325),
.Y(n_412)
);

AND2x2_ASAP7_75t_SL g413 ( 
.A(n_395),
.B(n_190),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_391),
.B(n_294),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_361),
.Y(n_415)
);

INVx6_ASAP7_75t_L g416 ( 
.A(n_388),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_366),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_380),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_370),
.A2(n_378),
.B1(n_381),
.B2(n_359),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_396),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_370),
.A2(n_281),
.B1(n_313),
.B2(n_299),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_396),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_364),
.Y(n_423)
);

INVx4_ASAP7_75t_L g424 ( 
.A(n_393),
.Y(n_424)
);

INVx2_ASAP7_75t_SL g425 ( 
.A(n_359),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_360),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_386),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_367),
.Y(n_428)
);

AND2x6_ASAP7_75t_L g429 ( 
.A(n_382),
.B(n_347),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_372),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_393),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_377),
.B(n_351),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_375),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_360),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_385),
.B(n_312),
.Y(n_435)
);

NOR2x1_ASAP7_75t_L g436 ( 
.A(n_381),
.B(n_289),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_358),
.B(n_282),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_389),
.B(n_297),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_378),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_363),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_392),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_363),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_368),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_365),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_368),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_374),
.B(n_298),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_364),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_368),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_365),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_368),
.A2(n_319),
.B1(n_331),
.B2(n_317),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_374),
.A2(n_349),
.B1(n_305),
.B2(n_303),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_381),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_365),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_368),
.B(n_337),
.Y(n_454)
);

INVxp33_ASAP7_75t_L g455 ( 
.A(n_382),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_359),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_368),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_365),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_356),
.Y(n_459)
);

BUFx8_ASAP7_75t_L g460 ( 
.A(n_384),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_359),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_362),
.B(n_308),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_365),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_368),
.Y(n_464)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_394),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_362),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_368),
.Y(n_467)
);

AOI22x1_ASAP7_75t_SL g468 ( 
.A1(n_359),
.A2(n_313),
.B1(n_281),
.B2(n_309),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_407),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_407),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_438),
.B(n_437),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_446),
.A2(n_301),
.B1(n_197),
.B2(n_336),
.Y(n_472)
);

XOR2x2_ASAP7_75t_L g473 ( 
.A(n_421),
.B(n_309),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_408),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_408),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_402),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_466),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_454),
.B(n_336),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_449),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_449),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_402),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_402),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_466),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_454),
.B(n_336),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_454),
.B(n_338),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_453),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_402),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_446),
.B(n_344),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_425),
.Y(n_489)
);

BUFx8_ASAP7_75t_L g490 ( 
.A(n_411),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_414),
.B(n_353),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_447),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_405),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_458),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_414),
.B(n_401),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_456),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_458),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_399),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_444),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_463),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_415),
.B(n_185),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_412),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_463),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_417),
.B(n_187),
.Y(n_504)
);

AND2x2_ASAP7_75t_SL g505 ( 
.A(n_413),
.B(n_190),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_447),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_492),
.Y(n_507)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_496),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_506),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_R g510 ( 
.A(n_490),
.B(n_456),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_469),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_R g512 ( 
.A(n_490),
.B(n_461),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_490),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_470),
.Y(n_514)
);

AND3x2_ASAP7_75t_L g515 ( 
.A(n_471),
.B(n_459),
.C(n_435),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_490),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_502),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_470),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_477),
.Y(n_519)
);

INVxp67_ASAP7_75t_SL g520 ( 
.A(n_483),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_479),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_469),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_498),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_473),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_R g525 ( 
.A(n_505),
.B(n_461),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_473),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_489),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_505),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_479),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_495),
.B(n_438),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_484),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_505),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_484),
.B(n_413),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_485),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_481),
.Y(n_535)
);

AND2x6_ASAP7_75t_L g536 ( 
.A(n_502),
.B(n_444),
.Y(n_536)
);

INVxp67_ASAP7_75t_SL g537 ( 
.A(n_481),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_481),
.Y(n_538)
);

NOR2xp67_ASAP7_75t_L g539 ( 
.A(n_476),
.B(n_424),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_R g540 ( 
.A(n_476),
.B(n_440),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_481),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_481),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_481),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_478),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_493),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_493),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_530),
.B(n_410),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_514),
.Y(n_548)
);

BUFx10_ASAP7_75t_L g549 ( 
.A(n_509),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_519),
.B(n_491),
.Y(n_550)
);

INVxp67_ASAP7_75t_SL g551 ( 
.A(n_537),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_524),
.A2(n_526),
.B1(n_528),
.B2(n_532),
.Y(n_552)
);

BUFx6f_ASAP7_75t_SL g553 ( 
.A(n_544),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_534),
.B(n_485),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_518),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_521),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_529),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_533),
.B(n_426),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_520),
.B(n_501),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_523),
.B(n_501),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_544),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_508),
.B(n_501),
.Y(n_562)
);

INVx4_ASAP7_75t_L g563 ( 
.A(n_509),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_528),
.B(n_502),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_515),
.B(n_501),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_527),
.B(n_426),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_536),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_525),
.B(n_488),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_511),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_531),
.B(n_442),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_531),
.B(n_504),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_535),
.B(n_493),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_536),
.Y(n_573)
);

NAND3xp33_ASAP7_75t_L g574 ( 
.A(n_539),
.B(n_472),
.C(n_422),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_511),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_542),
.B(n_493),
.Y(n_576)
);

AND2x6_ASAP7_75t_L g577 ( 
.A(n_517),
.B(n_493),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_522),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_522),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_543),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_507),
.Y(n_581)
);

INVx4_ASAP7_75t_L g582 ( 
.A(n_513),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_545),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_546),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_541),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_540),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_517),
.B(n_420),
.Y(n_587)
);

OR2x6_ASAP7_75t_L g588 ( 
.A(n_517),
.B(n_493),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_541),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_538),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_538),
.B(n_499),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_538),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_538),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_516),
.B(n_439),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_536),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_536),
.Y(n_596)
);

AND3x2_ASAP7_75t_L g597 ( 
.A(n_536),
.B(n_504),
.C(n_439),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_536),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_510),
.B(n_504),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_512),
.Y(n_600)
);

INVx5_ASAP7_75t_L g601 ( 
.A(n_536),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_530),
.B(n_499),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_509),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_530),
.B(n_442),
.Y(n_604)
);

BUFx10_ASAP7_75t_L g605 ( 
.A(n_509),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_514),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_511),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_511),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_530),
.B(n_504),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_514),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_514),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_514),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_514),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_514),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_530),
.B(n_427),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_530),
.A2(n_472),
.B1(n_417),
.B2(n_442),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_514),
.Y(n_617)
);

INVx8_ASAP7_75t_L g618 ( 
.A(n_536),
.Y(n_618)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_520),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_540),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_530),
.B(n_434),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_514),
.Y(n_622)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_520),
.Y(n_623)
);

INVxp67_ASAP7_75t_SL g624 ( 
.A(n_537),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_514),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_530),
.B(n_499),
.Y(n_626)
);

INVx4_ASAP7_75t_L g627 ( 
.A(n_509),
.Y(n_627)
);

BUFx10_ASAP7_75t_L g628 ( 
.A(n_509),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_507),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_507),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_610),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_612),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_620),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_548),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_555),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_561),
.Y(n_636)
);

INVxp33_ASAP7_75t_SL g637 ( 
.A(n_581),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_619),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_556),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_557),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_615),
.B(n_441),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_606),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_SL g643 ( 
.A1(n_615),
.A2(n_419),
.B1(n_440),
.B2(n_452),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_547),
.B(n_442),
.Y(n_644)
);

AND2x6_ASAP7_75t_L g645 ( 
.A(n_567),
.B(n_499),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_561),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_613),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_611),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_586),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_609),
.B(n_433),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_625),
.Y(n_651)
);

CKINVDCx6p67_ASAP7_75t_R g652 ( 
.A(n_603),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_614),
.Y(n_653)
);

AND2x2_ASAP7_75t_SL g654 ( 
.A(n_565),
.B(n_599),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_621),
.B(n_441),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_619),
.B(n_404),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_617),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_622),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_601),
.B(n_476),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_623),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_618),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_618),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_623),
.B(n_621),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_568),
.B(n_433),
.Y(n_664)
);

INVx4_ASAP7_75t_L g665 ( 
.A(n_582),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_559),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_550),
.B(n_423),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_575),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_560),
.B(n_452),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_578),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_604),
.B(n_423),
.Y(n_671)
);

BUFx4f_ASAP7_75t_L g672 ( 
.A(n_618),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_566),
.B(n_433),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_558),
.B(n_478),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_579),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_569),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_554),
.B(n_562),
.Y(n_677)
);

INVx4_ASAP7_75t_L g678 ( 
.A(n_582),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_569),
.Y(n_679)
);

AND2x6_ASAP7_75t_L g680 ( 
.A(n_567),
.B(n_499),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_570),
.B(n_478),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_566),
.B(n_433),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_607),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_601),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_568),
.B(n_465),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_629),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_552),
.B(n_465),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_549),
.Y(n_688)
);

AND2x6_ASAP7_75t_L g689 ( 
.A(n_573),
.B(n_499),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_571),
.B(n_478),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_607),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_608),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_608),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_585),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_589),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_602),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_602),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_577),
.Y(n_698)
);

INVx8_ASAP7_75t_L g699 ( 
.A(n_630),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_587),
.B(n_428),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_563),
.B(n_428),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_587),
.B(n_430),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_549),
.Y(n_703)
);

INVx5_ASAP7_75t_L g704 ( 
.A(n_601),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_601),
.B(n_476),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_580),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_584),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_577),
.Y(n_708)
);

CKINVDCx8_ASAP7_75t_R g709 ( 
.A(n_594),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_563),
.B(n_430),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_626),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_605),
.Y(n_712)
);

OR2x2_ASAP7_75t_L g713 ( 
.A(n_626),
.B(n_431),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_583),
.B(n_480),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_551),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_668),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_668),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_638),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_684),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_641),
.B(n_655),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_634),
.Y(n_721)
);

INVx4_ASAP7_75t_L g722 ( 
.A(n_704),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_684),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_635),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_663),
.B(n_551),
.Y(n_725)
);

NAND3xp33_ASAP7_75t_L g726 ( 
.A(n_696),
.B(n_574),
.C(n_616),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_698),
.B(n_573),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_679),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_691),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_677),
.B(n_624),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_639),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_666),
.B(n_624),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_664),
.B(n_600),
.Y(n_733)
);

BUFx10_ASAP7_75t_L g734 ( 
.A(n_673),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_684),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_643),
.A2(n_616),
.B1(n_418),
.B2(n_412),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_706),
.B(n_572),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_682),
.B(n_594),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_706),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_675),
.Y(n_740)
);

INVx2_ASAP7_75t_SL g741 ( 
.A(n_706),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_676),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_683),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_660),
.B(n_644),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_700),
.B(n_572),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_702),
.B(n_576),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_692),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_674),
.B(n_627),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_693),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_661),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_698),
.B(n_598),
.Y(n_751)
);

AO22x2_ASAP7_75t_L g752 ( 
.A1(n_653),
.A2(n_564),
.B1(n_596),
.B2(n_595),
.Y(n_752)
);

OR2x2_ASAP7_75t_L g753 ( 
.A(n_640),
.B(n_590),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_642),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_685),
.B(n_576),
.Y(n_755)
);

OR2x2_ASAP7_75t_SL g756 ( 
.A(n_669),
.B(n_416),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_670),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_648),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_651),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_631),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_632),
.Y(n_761)
);

OAI221xp5_ASAP7_75t_L g762 ( 
.A1(n_667),
.A2(n_436),
.B1(n_400),
.B2(n_451),
.C(n_455),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_707),
.B(n_627),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_657),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_647),
.Y(n_765)
);

BUFx2_ASAP7_75t_L g766 ( 
.A(n_707),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_661),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_707),
.B(n_592),
.Y(n_768)
);

BUFx2_ASAP7_75t_L g769 ( 
.A(n_633),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_656),
.B(n_592),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_708),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_709),
.B(n_455),
.Y(n_772)
);

INVx4_ASAP7_75t_L g773 ( 
.A(n_704),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_658),
.Y(n_774)
);

INVx8_ASAP7_75t_L g775 ( 
.A(n_704),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_694),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_695),
.B(n_593),
.Y(n_777)
);

INVx4_ASAP7_75t_L g778 ( 
.A(n_708),
.Y(n_778)
);

OR2x2_ASAP7_75t_L g779 ( 
.A(n_715),
.B(n_593),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_715),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_697),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_671),
.B(n_577),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_711),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_714),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_713),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_636),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_681),
.B(n_588),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_633),
.B(n_650),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_636),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_646),
.B(n_577),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_716),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_726),
.A2(n_654),
.B1(n_564),
.B2(n_597),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_720),
.B(n_665),
.Y(n_793)
);

NAND2xp33_ASAP7_75t_L g794 ( 
.A(n_750),
.B(n_712),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_720),
.B(n_665),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_734),
.B(n_738),
.Y(n_796)
);

INVx2_ASAP7_75t_SL g797 ( 
.A(n_763),
.Y(n_797)
);

INVxp67_ASAP7_75t_L g798 ( 
.A(n_769),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_734),
.B(n_678),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_771),
.B(n_646),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_739),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_736),
.A2(n_597),
.B1(n_690),
.B2(n_475),
.Y(n_802)
);

NAND3xp33_ASAP7_75t_L g803 ( 
.A(n_781),
.B(n_710),
.C(n_701),
.Y(n_803)
);

CKINVDCx11_ASAP7_75t_R g804 ( 
.A(n_734),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_736),
.A2(n_475),
.B1(n_486),
.B2(n_474),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_748),
.B(n_652),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_718),
.B(n_688),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_785),
.B(n_649),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_716),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_R g810 ( 
.A(n_750),
.B(n_686),
.Y(n_810)
);

NAND2xp33_ASAP7_75t_L g811 ( 
.A(n_750),
.B(n_699),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_725),
.B(n_678),
.Y(n_812)
);

NOR2x1p5_ASAP7_75t_L g813 ( 
.A(n_771),
.B(n_649),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_730),
.B(n_645),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_719),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_762),
.A2(n_486),
.B1(n_494),
.B2(n_474),
.Y(n_816)
);

AO22x1_ASAP7_75t_L g817 ( 
.A1(n_784),
.A2(n_460),
.B1(n_397),
.B2(n_645),
.Y(n_817)
);

NOR2xp67_ASAP7_75t_L g818 ( 
.A(n_778),
.B(n_649),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_783),
.Y(n_819)
);

AND2x4_ASAP7_75t_SL g820 ( 
.A(n_750),
.B(n_605),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_732),
.B(n_645),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_717),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_772),
.B(n_637),
.Y(n_823)
);

BUFx3_ASAP7_75t_L g824 ( 
.A(n_766),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_772),
.B(n_703),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_744),
.B(n_645),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_780),
.B(n_680),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_767),
.B(n_788),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_739),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_767),
.B(n_661),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_776),
.B(n_680),
.Y(n_831)
);

AO22x1_ASAP7_75t_L g832 ( 
.A1(n_733),
.A2(n_460),
.B1(n_397),
.B2(n_680),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_717),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_733),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_776),
.B(n_680),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_767),
.B(n_662),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_752),
.A2(n_553),
.B1(n_687),
.B2(n_672),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_778),
.Y(n_838)
);

OR2x6_ASAP7_75t_L g839 ( 
.A(n_775),
.B(n_662),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_721),
.B(n_724),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_785),
.Y(n_841)
);

INVx2_ASAP7_75t_SL g842 ( 
.A(n_741),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_752),
.A2(n_497),
.B1(n_500),
.B2(n_494),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_757),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_767),
.B(n_662),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_731),
.B(n_689),
.Y(n_846)
);

INVx8_ASAP7_75t_L g847 ( 
.A(n_775),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_754),
.B(n_689),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_752),
.A2(n_500),
.B1(n_503),
.B2(n_497),
.Y(n_849)
);

BUFx8_ASAP7_75t_L g850 ( 
.A(n_741),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_758),
.B(n_689),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_759),
.B(n_689),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_757),
.B(n_577),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_770),
.B(n_591),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_760),
.Y(n_855)
);

INVxp67_ASAP7_75t_L g856 ( 
.A(n_768),
.Y(n_856)
);

AND2x6_ASAP7_75t_SL g857 ( 
.A(n_788),
.B(n_699),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_787),
.B(n_628),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_771),
.B(n_628),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_778),
.B(n_751),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_760),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_SL g862 ( 
.A(n_722),
.B(n_672),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_751),
.B(n_659),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_789),
.B(n_659),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_782),
.B(n_705),
.Y(n_865)
);

NAND2xp33_ASAP7_75t_L g866 ( 
.A(n_790),
.B(n_431),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_745),
.B(n_416),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_761),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_746),
.B(n_416),
.Y(n_869)
);

AO22x1_ASAP7_75t_L g870 ( 
.A1(n_764),
.A2(n_460),
.B1(n_397),
.B2(n_705),
.Y(n_870)
);

O2A1O1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_737),
.A2(n_755),
.B(n_198),
.C(n_200),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_810),
.B(n_719),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_807),
.Y(n_873)
);

OR2x2_ASAP7_75t_L g874 ( 
.A(n_854),
.B(n_779),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_857),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_L g876 ( 
.A1(n_834),
.A2(n_755),
.B1(n_756),
.B2(n_737),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_803),
.B(n_804),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_840),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_797),
.B(n_789),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_854),
.B(n_786),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_840),
.Y(n_881)
);

INVx4_ASAP7_75t_L g882 ( 
.A(n_820),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_800),
.B(n_719),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_791),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_819),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_798),
.B(n_777),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_844),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_812),
.B(n_753),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_814),
.B(n_727),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_826),
.B(n_727),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_796),
.B(n_468),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_821),
.B(n_727),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_846),
.B(n_742),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_809),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_815),
.Y(n_895)
);

INVxp67_ASAP7_75t_SL g896 ( 
.A(n_827),
.Y(n_896)
);

INVx1_ASAP7_75t_SL g897 ( 
.A(n_806),
.Y(n_897)
);

INVxp67_ASAP7_75t_L g898 ( 
.A(n_827),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_816),
.A2(n_418),
.B1(n_403),
.B2(n_409),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_R g900 ( 
.A(n_794),
.B(n_811),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_846),
.B(n_848),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_822),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_848),
.B(n_742),
.Y(n_903)
);

INVx1_ASAP7_75t_SL g904 ( 
.A(n_858),
.Y(n_904)
);

INVx4_ASAP7_75t_L g905 ( 
.A(n_847),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_802),
.A2(n_418),
.B1(n_443),
.B2(n_398),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_815),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_793),
.B(n_431),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_851),
.B(n_743),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_833),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_855),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_800),
.B(n_719),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_866),
.A2(n_591),
.B(n_775),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_792),
.A2(n_418),
.B1(n_448),
.B2(n_445),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_860),
.B(n_723),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_841),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_851),
.Y(n_917)
);

NOR2xp67_ASAP7_75t_L g918 ( 
.A(n_837),
.B(n_838),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_860),
.B(n_723),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_852),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_818),
.B(n_723),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_861),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_852),
.B(n_831),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_868),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_831),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_835),
.B(n_743),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_835),
.B(n_747),
.Y(n_927)
);

OR2x6_ASAP7_75t_L g928 ( 
.A(n_817),
.B(n_775),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_878),
.B(n_808),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_876),
.A2(n_871),
.B(n_849),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_877),
.A2(n_843),
.B(n_795),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_901),
.A2(n_828),
.B(n_799),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_881),
.B(n_880),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_928),
.A2(n_832),
.B(n_865),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_900),
.B(n_859),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_917),
.B(n_801),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_920),
.B(n_829),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_904),
.B(n_824),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_918),
.B(n_863),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_L g940 ( 
.A1(n_898),
.A2(n_823),
.B(n_825),
.Y(n_940)
);

BUFx4f_ASAP7_75t_L g941 ( 
.A(n_928),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_898),
.B(n_842),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_925),
.B(n_856),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_873),
.B(n_879),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_928),
.A2(n_870),
.B(n_853),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_875),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_877),
.A2(n_869),
.B(n_867),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_923),
.A2(n_853),
.B(n_836),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_897),
.B(n_431),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_889),
.B(n_813),
.Y(n_950)
);

OAI21x1_ASAP7_75t_L g951 ( 
.A1(n_926),
.A2(n_838),
.B(n_749),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_896),
.B(n_864),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_882),
.B(n_863),
.Y(n_953)
);

O2A1O1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_891),
.A2(n_845),
.B(n_830),
.C(n_201),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_884),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_891),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_882),
.B(n_850),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_885),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_872),
.A2(n_862),
.B(n_839),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_874),
.B(n_815),
.Y(n_960)
);

AOI21x1_ASAP7_75t_L g961 ( 
.A1(n_927),
.A2(n_839),
.B(n_751),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_896),
.A2(n_862),
.B(n_839),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_893),
.B(n_850),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_883),
.A2(n_847),
.B(n_773),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_895),
.B(n_723),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_912),
.A2(n_847),
.B(n_773),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_921),
.A2(n_773),
.B(n_722),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_892),
.A2(n_805),
.B1(n_735),
.B2(n_722),
.Y(n_968)
);

NOR3xp33_ASAP7_75t_L g969 ( 
.A(n_908),
.B(n_465),
.C(n_424),
.Y(n_969)
);

BUFx3_ASAP7_75t_L g970 ( 
.A(n_886),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_903),
.B(n_747),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_890),
.A2(n_735),
.B1(n_588),
.B2(n_598),
.Y(n_972)
);

AO21x1_ASAP7_75t_L g973 ( 
.A1(n_909),
.A2(n_406),
.B(n_749),
.Y(n_973)
);

INVx4_ASAP7_75t_L g974 ( 
.A(n_905),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_915),
.A2(n_735),
.B(n_588),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_914),
.A2(n_193),
.B(n_208),
.C(n_205),
.Y(n_976)
);

AO21x1_ASAP7_75t_L g977 ( 
.A1(n_908),
.A2(n_406),
.B(n_424),
.Y(n_977)
);

AOI22xp33_ASAP7_75t_L g978 ( 
.A1(n_914),
.A2(n_906),
.B1(n_899),
.B2(n_887),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_894),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_905),
.B(n_888),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_919),
.A2(n_735),
.B(n_761),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_906),
.A2(n_553),
.B1(n_774),
.B2(n_765),
.Y(n_982)
);

AND2x4_ASAP7_75t_SL g983 ( 
.A(n_895),
.B(n_765),
.Y(n_983)
);

AOI21xp33_ASAP7_75t_L g984 ( 
.A1(n_916),
.A2(n_774),
.B(n_210),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_913),
.A2(n_740),
.B(n_729),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_913),
.A2(n_740),
.B(n_729),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_895),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_907),
.B(n_728),
.Y(n_988)
);

AOI21x1_ASAP7_75t_L g989 ( 
.A1(n_902),
.A2(n_728),
.B(n_432),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_907),
.B(n_462),
.Y(n_990)
);

OR2x2_ASAP7_75t_L g991 ( 
.A(n_910),
.B(n_0),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_907),
.A2(n_432),
.B(n_211),
.Y(n_992)
);

INVx4_ASAP7_75t_L g993 ( 
.A(n_911),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_922),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_958),
.B(n_924),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_950),
.B(n_899),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_941),
.A2(n_212),
.B(n_209),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_946),
.B(n_0),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_944),
.B(n_1),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_941),
.B(n_482),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_939),
.A2(n_216),
.B(n_215),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_970),
.B(n_1),
.Y(n_1002)
);

NAND2xp33_ASAP7_75t_L g1003 ( 
.A(n_956),
.B(n_429),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_930),
.A2(n_219),
.B(n_217),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_957),
.B(n_2),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_933),
.B(n_2),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_943),
.B(n_3),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_971),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_930),
.A2(n_225),
.B(n_224),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_987),
.Y(n_1010)
);

BUFx2_ASAP7_75t_L g1011 ( 
.A(n_974),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_952),
.B(n_932),
.Y(n_1012)
);

OAI21xp33_ASAP7_75t_L g1013 ( 
.A1(n_942),
.A2(n_227),
.B(n_233),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_934),
.A2(n_487),
.B(n_482),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_974),
.B(n_3),
.Y(n_1015)
);

OAI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_1004),
.A2(n_931),
.B(n_962),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_1011),
.B(n_938),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_1009),
.A2(n_935),
.B(n_931),
.Y(n_1018)
);

NOR3xp33_ASAP7_75t_L g1019 ( 
.A(n_1013),
.B(n_954),
.C(n_969),
.Y(n_1019)
);

AOI21x1_ASAP7_75t_SL g1020 ( 
.A1(n_1012),
.A2(n_1007),
.B(n_1006),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_1002),
.A2(n_940),
.B(n_953),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_1005),
.A2(n_973),
.B(n_977),
.Y(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_1015),
.A2(n_976),
.B(n_991),
.C(n_984),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_998),
.B(n_980),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_1010),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_1010),
.Y(n_1026)
);

AOI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_996),
.A2(n_978),
.B1(n_949),
.B2(n_990),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_1001),
.A2(n_945),
.B(n_947),
.C(n_948),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_SL g1029 ( 
.A(n_999),
.B(n_959),
.Y(n_1029)
);

OR2x6_ASAP7_75t_L g1030 ( 
.A(n_997),
.B(n_947),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_1008),
.A2(n_975),
.B(n_986),
.C(n_985),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_L g1032 ( 
.A1(n_995),
.A2(n_951),
.B(n_961),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_995),
.Y(n_1033)
);

HB1xp67_ASAP7_75t_L g1034 ( 
.A(n_1000),
.Y(n_1034)
);

AO32x1_ASAP7_75t_L g1035 ( 
.A1(n_1003),
.A2(n_993),
.A3(n_968),
.B1(n_972),
.B2(n_983),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_SL g1036 ( 
.A1(n_1014),
.A2(n_963),
.B1(n_987),
.B2(n_936),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_1012),
.B(n_987),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1012),
.B(n_993),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_1010),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_1004),
.A2(n_992),
.B(n_960),
.C(n_937),
.Y(n_1040)
);

OR2x2_ASAP7_75t_L g1041 ( 
.A(n_1033),
.B(n_929),
.Y(n_1041)
);

OR2x2_ASAP7_75t_L g1042 ( 
.A(n_1038),
.B(n_981),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_1029),
.B(n_964),
.Y(n_1043)
);

NAND2x1p5_ASAP7_75t_L g1044 ( 
.A(n_1017),
.B(n_965),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_1030),
.A2(n_967),
.B(n_966),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_1017),
.B(n_988),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_1030),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1047),
.B(n_1018),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_1044),
.A2(n_1026),
.B(n_1025),
.Y(n_1049)
);

AO21x2_ASAP7_75t_L g1050 ( 
.A1(n_1048),
.A2(n_1028),
.B(n_1043),
.Y(n_1050)
);

AO21x2_ASAP7_75t_L g1051 ( 
.A1(n_1049),
.A2(n_1037),
.B(n_1016),
.Y(n_1051)
);

INVx2_ASAP7_75t_SL g1052 ( 
.A(n_1049),
.Y(n_1052)
);

NAND2x1_ASAP7_75t_L g1053 ( 
.A(n_1052),
.B(n_1046),
.Y(n_1053)
);

OAI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_1051),
.A2(n_1022),
.B1(n_1027),
.B2(n_1045),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_1050),
.B(n_1024),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_1055),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1053),
.Y(n_1057)
);

AO31x2_ASAP7_75t_L g1058 ( 
.A1(n_1057),
.A2(n_1054),
.A3(n_1050),
.B(n_1051),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_1057),
.A2(n_1020),
.B(n_1042),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_1059),
.B(n_1056),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1058),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_1060),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_1061),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_1062),
.A2(n_1039),
.B1(n_1019),
.B2(n_1058),
.Y(n_1064)
);

OAI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_1063),
.A2(n_1041),
.B1(n_1021),
.B2(n_1034),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_1064),
.A2(n_1063),
.B1(n_1036),
.B2(n_1032),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_1065),
.A2(n_1031),
.B1(n_1040),
.B2(n_1023),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1067),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1066),
.B(n_1035),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1067),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1068),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1070),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_1069),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_1073),
.B(n_1035),
.Y(n_1074)
);

OAI221xp5_ASAP7_75t_SL g1075 ( 
.A1(n_1071),
.A2(n_1035),
.B1(n_457),
.B2(n_467),
.C(n_464),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_1074),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_1075),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1076),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_1077),
.B(n_1072),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_1078),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_1079),
.B(n_955),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1080),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_1081),
.B(n_979),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_1082),
.B(n_1083),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1082),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_1084),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1085),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1085),
.Y(n_1088)
);

OR2x2_ASAP7_75t_L g1089 ( 
.A(n_1086),
.B(n_4),
.Y(n_1089)
);

OR2x2_ASAP7_75t_L g1090 ( 
.A(n_1087),
.B(n_5),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1088),
.B(n_5),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_1089),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_1090),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1093),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1092),
.Y(n_1095)
);

NAND2x1p5_ASAP7_75t_L g1096 ( 
.A(n_1094),
.B(n_1091),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1095),
.Y(n_1097)
);

OAI211xp5_ASAP7_75t_SL g1098 ( 
.A1(n_1097),
.A2(n_195),
.B(n_191),
.C(n_202),
.Y(n_1098)
);

INVx1_ASAP7_75t_SL g1099 ( 
.A(n_1096),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_1099),
.A2(n_221),
.B(n_204),
.C(n_207),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1098),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_1101),
.A2(n_189),
.B1(n_195),
.B2(n_213),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1100),
.B(n_6),
.Y(n_1103)
);

AOI21xp33_ASAP7_75t_L g1104 ( 
.A1(n_1102),
.A2(n_220),
.B(n_218),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_1103),
.B(n_7),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1103),
.B(n_8),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_1106),
.B(n_1105),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_1104),
.B(n_195),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1104),
.A2(n_228),
.B(n_226),
.Y(n_1109)
);

AOI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1107),
.A2(n_195),
.B1(n_232),
.B2(n_230),
.Y(n_1110)
);

AOI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_1108),
.A2(n_195),
.B1(n_231),
.B2(n_189),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1111),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_1110),
.Y(n_1113)
);

AOI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1113),
.A2(n_1109),
.B1(n_195),
.B2(n_189),
.Y(n_1114)
);

INVx1_ASAP7_75t_SL g1115 ( 
.A(n_1112),
.Y(n_1115)
);

OAI211xp5_ASAP7_75t_L g1116 ( 
.A1(n_1115),
.A2(n_189),
.B(n_9),
.C(n_10),
.Y(n_1116)
);

INVx1_ASAP7_75t_SL g1117 ( 
.A(n_1114),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_1117),
.B(n_195),
.Y(n_1118)
);

NOR2x1_ASAP7_75t_L g1119 ( 
.A(n_1116),
.B(n_310),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1118),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1119),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1120),
.A2(n_450),
.B(n_310),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_1121),
.B(n_8),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1121),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1124),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1123),
.B(n_10),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_1122),
.B(n_11),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1125),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1126),
.Y(n_1129)
);

INVxp67_ASAP7_75t_SL g1130 ( 
.A(n_1128),
.Y(n_1130)
);

NAND4xp75_ASAP7_75t_L g1131 ( 
.A(n_1129),
.B(n_1127),
.C(n_13),
.D(n_14),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_SL g1132 ( 
.A1(n_1130),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1131),
.A2(n_12),
.B1(n_15),
.B2(n_17),
.Y(n_1133)
);

OR3x2_ASAP7_75t_L g1134 ( 
.A(n_1133),
.B(n_15),
.C(n_18),
.Y(n_1134)
);

OAI211xp5_ASAP7_75t_L g1135 ( 
.A1(n_1132),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_1135)
);

OAI211xp5_ASAP7_75t_SL g1136 ( 
.A1(n_1134),
.A2(n_19),
.B(n_20),
.C(n_21),
.Y(n_1136)
);

NOR2x1_ASAP7_75t_L g1137 ( 
.A(n_1135),
.B(n_22),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1137),
.A2(n_1136),
.B(n_22),
.Y(n_1138)
);

AND2x4_ASAP7_75t_L g1139 ( 
.A(n_1137),
.B(n_23),
.Y(n_1139)
);

XOR2x1_ASAP7_75t_L g1140 ( 
.A(n_1139),
.B(n_23),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_R g1141 ( 
.A(n_1138),
.B(n_24),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1139),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1140),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1141),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1142),
.Y(n_1145)
);

AO22x2_ASAP7_75t_L g1146 ( 
.A1(n_1145),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1144),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1147),
.Y(n_1148)
);

OAI221xp5_ASAP7_75t_L g1149 ( 
.A1(n_1146),
.A2(n_1143),
.B1(n_26),
.B2(n_27),
.C(n_28),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1148),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1149),
.Y(n_1151)
);

AO22x2_ASAP7_75t_L g1152 ( 
.A1(n_1150),
.A2(n_25),
.B1(n_27),
.B2(n_29),
.Y(n_1152)
);

AOI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1151),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_1153)
);

OAI22x1_ASAP7_75t_L g1154 ( 
.A1(n_1153),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_1154)
);

OAI22x1_ASAP7_75t_L g1155 ( 
.A1(n_1152),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_1155)
);

OR2x2_ASAP7_75t_L g1156 ( 
.A(n_1154),
.B(n_33),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_1155),
.Y(n_1157)
);

CKINVDCx20_ASAP7_75t_R g1158 ( 
.A(n_1154),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1157),
.Y(n_1159)
);

NAND3xp33_ASAP7_75t_L g1160 ( 
.A(n_1158),
.B(n_36),
.C(n_37),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1156),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1157),
.A2(n_41),
.B(n_42),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1159),
.A2(n_44),
.B(n_45),
.Y(n_1163)
);

AO21x2_ASAP7_75t_L g1164 ( 
.A1(n_1160),
.A2(n_46),
.B(n_49),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1162),
.A2(n_50),
.B(n_51),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1161),
.B(n_52),
.Y(n_1166)
);

AO22x2_ASAP7_75t_L g1167 ( 
.A1(n_1163),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_1167)
);

OAI222xp33_ASAP7_75t_L g1168 ( 
.A1(n_1164),
.A2(n_1166),
.B1(n_1165),
.B2(n_60),
.C1(n_61),
.C2(n_63),
.Y(n_1168)
);

AOI222xp33_ASAP7_75t_L g1169 ( 
.A1(n_1163),
.A2(n_57),
.B1(n_58),
.B2(n_64),
.C1(n_65),
.C2(n_66),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1164),
.A2(n_69),
.B(n_72),
.Y(n_1170)
);

NAND3xp33_ASAP7_75t_L g1171 ( 
.A(n_1163),
.B(n_73),
.C(n_76),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1164),
.Y(n_1172)
);

AOI221xp5_ASAP7_75t_L g1173 ( 
.A1(n_1163),
.A2(n_79),
.B1(n_80),
.B2(n_82),
.C(n_83),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1164),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1164),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_1175)
);

AOI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1164),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_1176)
);

OAI222xp33_ASAP7_75t_L g1177 ( 
.A1(n_1163),
.A2(n_91),
.B1(n_92),
.B2(n_94),
.C1(n_95),
.C2(n_96),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1164),
.A2(n_97),
.B(n_98),
.Y(n_1178)
);

AOI32xp33_ASAP7_75t_L g1179 ( 
.A1(n_1175),
.A2(n_100),
.A3(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_1179)
);

AO221x1_ASAP7_75t_L g1180 ( 
.A1(n_1171),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.C(n_109),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_SL g1181 ( 
.A1(n_1176),
.A2(n_110),
.B(n_112),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1169),
.A2(n_113),
.B1(n_114),
.B2(n_119),
.Y(n_1182)
);

AOI221xp5_ASAP7_75t_L g1183 ( 
.A1(n_1173),
.A2(n_120),
.B1(n_121),
.B2(n_123),
.C(n_126),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1174),
.B(n_128),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1177),
.A2(n_130),
.B(n_132),
.Y(n_1185)
);

AOI21xp33_ASAP7_75t_SL g1186 ( 
.A1(n_1168),
.A2(n_133),
.B(n_134),
.Y(n_1186)
);

AOI221xp5_ASAP7_75t_L g1187 ( 
.A1(n_1170),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.C(n_138),
.Y(n_1187)
);

AOI221xp5_ASAP7_75t_L g1188 ( 
.A1(n_1180),
.A2(n_1178),
.B1(n_1167),
.B2(n_1172),
.C(n_143),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_1181),
.Y(n_1189)
);

NOR3xp33_ASAP7_75t_SL g1190 ( 
.A(n_1187),
.B(n_1167),
.C(n_140),
.Y(n_1190)
);

INVx1_ASAP7_75t_SL g1191 ( 
.A(n_1184),
.Y(n_1191)
);

NOR2xp67_ASAP7_75t_L g1192 ( 
.A(n_1186),
.B(n_139),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1182),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1183),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_SL g1195 ( 
.A1(n_1191),
.A2(n_1185),
.B1(n_1179),
.B2(n_147),
.Y(n_1195)
);

NOR3xp33_ASAP7_75t_L g1196 ( 
.A(n_1194),
.B(n_142),
.C(n_146),
.Y(n_1196)
);

AOI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1193),
.A2(n_148),
.B(n_150),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1192),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1196),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1199),
.A2(n_1195),
.B1(n_1198),
.B2(n_1197),
.Y(n_1200)
);

AOI21xp33_ASAP7_75t_SL g1201 ( 
.A1(n_1200),
.A2(n_1189),
.B(n_1190),
.Y(n_1201)
);

OAI21xp33_ASAP7_75t_L g1202 ( 
.A1(n_1201),
.A2(n_1188),
.B(n_982),
.Y(n_1202)
);

OAI221xp5_ASAP7_75t_R g1203 ( 
.A1(n_1202),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.C(n_161),
.Y(n_1203)
);

AOI221xp5_ASAP7_75t_L g1204 ( 
.A1(n_1203),
.A2(n_163),
.B1(n_165),
.B2(n_166),
.C(n_167),
.Y(n_1204)
);

AOI21xp33_ASAP7_75t_SL g1205 ( 
.A1(n_1204),
.A2(n_168),
.B(n_173),
.Y(n_1205)
);

AOI211xp5_ASAP7_75t_L g1206 ( 
.A1(n_1205),
.A2(n_994),
.B(n_176),
.C(n_178),
.Y(n_1206)
);

AOI211xp5_ASAP7_75t_L g1207 ( 
.A1(n_1206),
.A2(n_174),
.B(n_989),
.C(n_482),
.Y(n_1207)
);


endmodule