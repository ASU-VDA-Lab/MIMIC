module fake_jpeg_5767_n_284 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_284);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_32),
.B1(n_24),
.B2(n_26),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_22),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_38),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_21),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_40),
.Y(n_49)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_41),
.B(n_44),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_43),
.Y(n_81)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NAND3xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_17),
.C(n_19),
.Y(n_45)
);

NAND3xp33_ASAP7_75t_SL g65 ( 
.A(n_45),
.B(n_36),
.C(n_29),
.Y(n_65)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_51),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_17),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_52),
.Y(n_60)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_22),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_38),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_56),
.Y(n_66)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_59),
.Y(n_88)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_53),
.A2(n_32),
.B1(n_24),
.B2(n_40),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_55),
.A2(n_32),
.B1(n_24),
.B2(n_40),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_64),
.Y(n_91)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_67),
.Y(n_96)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_72),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_41),
.A2(n_39),
.B1(n_19),
.B2(n_29),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_71),
.A2(n_23),
.B1(n_31),
.B2(n_30),
.Y(n_99)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_33),
.B1(n_38),
.B2(n_37),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_74),
.A2(n_33),
.B1(n_22),
.B2(n_27),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_75),
.B(n_25),
.Y(n_94)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_76),
.Y(n_111)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_79),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_46),
.A2(n_39),
.B1(n_44),
.B2(n_38),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_25),
.B1(n_30),
.B2(n_33),
.Y(n_102)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_82),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_27),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_31),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_85),
.B(n_86),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_56),
.B(n_23),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_89),
.A2(n_100),
.B(n_86),
.Y(n_120)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_95),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_33),
.B1(n_37),
.B2(n_27),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_105),
.B1(n_111),
.B2(n_73),
.Y(n_114)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_60),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_70),
.A2(n_58),
.B1(n_59),
.B2(n_74),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_102),
.B1(n_64),
.B2(n_81),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_99),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_75),
.A2(n_33),
.B(n_37),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_37),
.B1(n_21),
.B2(n_20),
.Y(n_105)
);

HB1xp67_ASAP7_75t_SL g106 ( 
.A(n_74),
.Y(n_106)
);

NOR2xp67_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_105),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_28),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_110),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_28),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_69),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_114),
.A2(n_122),
.B1(n_123),
.B2(n_111),
.Y(n_165)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_116),
.B(n_119),
.Y(n_158)
);

MAJx2_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_74),
.C(n_67),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_130),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_118),
.A2(n_126),
.B(n_85),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_120),
.A2(n_94),
.B1(n_99),
.B2(n_88),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_60),
.Y(n_121)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_105),
.A2(n_70),
.B1(n_77),
.B2(n_79),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_66),
.B(n_63),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_77),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_66),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_141),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_132),
.B(n_140),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_95),
.C(n_113),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_108),
.Y(n_147)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_135),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_139),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_72),
.Y(n_137)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_137),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_91),
.B(n_21),
.Y(n_138)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_91),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_89),
.B(n_28),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_120),
.A2(n_107),
.B(n_110),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_142),
.A2(n_169),
.B(n_171),
.Y(n_192)
);

AND2x4_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_102),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_146),
.A2(n_148),
.B(n_153),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_133),
.C(n_129),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_97),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_134),
.A2(n_90),
.B1(n_87),
.B2(n_96),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_149),
.A2(n_170),
.B1(n_122),
.B2(n_123),
.Y(n_175)
);

AND2x6_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_96),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_129),
.Y(n_178)
);

NAND2xp33_ASAP7_75t_SL g153 ( 
.A(n_117),
.B(n_88),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_141),
.Y(n_181)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_159),
.Y(n_186)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_18),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_131),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_164),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_116),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_165),
.A2(n_20),
.B1(n_18),
.B2(n_127),
.Y(n_187)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_168),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_101),
.Y(n_167)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_124),
.A2(n_103),
.B1(n_101),
.B2(n_21),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_117),
.A2(n_20),
.B(n_18),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_165),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_180),
.C(n_185),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_146),
.A2(n_124),
.B1(n_141),
.B2(n_125),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_177),
.A2(n_196),
.B(n_154),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_181),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_161),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_182),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_139),
.C(n_114),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_143),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_190),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_125),
.C(n_136),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_187),
.A2(n_170),
.B1(n_157),
.B2(n_150),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_127),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_189),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_142),
.B(n_20),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_146),
.A2(n_151),
.B1(n_144),
.B2(n_160),
.Y(n_191)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_191),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_156),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_195),
.Y(n_215)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_18),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_146),
.B(n_147),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_144),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_198),
.A2(n_200),
.B1(n_1),
.B2(n_2),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_183),
.A2(n_153),
.B1(n_152),
.B2(n_144),
.Y(n_199)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

INVx11_ASAP7_75t_L g200 ( 
.A(n_186),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_191),
.B(n_184),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_208),
.C(n_216),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_148),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_211),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_181),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_184),
.B(n_148),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_212),
.A2(n_159),
.B1(n_2),
.B2(n_3),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_174),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_217),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_180),
.A2(n_192),
.B(n_185),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_173),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_178),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_221),
.Y(n_240)
);

NAND2xp33_ASAP7_75t_R g220 ( 
.A(n_201),
.B(n_188),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_220),
.A2(n_228),
.B(n_231),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_176),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_223),
.C(n_226),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_189),
.C(n_177),
.Y(n_223)
);

OA21x2_ASAP7_75t_L g224 ( 
.A1(n_204),
.A2(n_172),
.B(n_175),
.Y(n_224)
);

OA21x2_ASAP7_75t_L g243 ( 
.A1(n_224),
.A2(n_211),
.B(n_206),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_149),
.C(n_196),
.Y(n_226)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_227),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_1),
.Y(n_228)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_229),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_4),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_4),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_233),
.A2(n_207),
.B(n_215),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_203),
.B(n_4),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_234),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_230),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_237),
.A2(n_239),
.B(n_241),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_232),
.A2(n_205),
.B1(n_199),
.B2(n_210),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_242),
.A2(n_244),
.B1(n_5),
.B2(n_6),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_5),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_224),
.A2(n_200),
.B1(n_214),
.B2(n_8),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_225),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_247),
.B(n_218),
.Y(n_249)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_237),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_248),
.B(n_251),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_8),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_235),
.A2(n_224),
.B1(n_223),
.B2(n_219),
.Y(n_250)
);

O2A1O1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_250),
.A2(n_246),
.B(n_9),
.C(n_10),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_245),
.B(n_233),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_243),
.B(n_218),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_258),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_253),
.A2(n_255),
.B1(n_256),
.B2(n_11),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_239),
.A2(n_243),
.B1(n_238),
.B2(n_247),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_6),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_257),
.B(n_10),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_240),
.C(n_236),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_260),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_263),
.Y(n_270)
);

OAI321xp33_ASAP7_75t_L g262 ( 
.A1(n_255),
.A2(n_15),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C(n_11),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_262),
.A2(n_265),
.B(n_13),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_11),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_12),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_13),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_258),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_269),
.B(n_273),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_272),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_14),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_266),
.Y(n_274)
);

NOR2x1_ASAP7_75t_SL g277 ( 
.A(n_274),
.B(n_15),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_252),
.Y(n_275)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_275),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_277),
.B(n_270),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_279),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_280),
.C(n_275),
.Y(n_282)
);

NOR3xp33_ASAP7_75t_SL g283 ( 
.A(n_282),
.B(n_276),
.C(n_268),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_278),
.Y(n_284)
);


endmodule