module fake_ibex_1134_n_885 (n_151, n_147, n_85, n_128, n_84, n_64, n_3, n_73, n_152, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_120, n_93, n_155, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_885);

input n_151;
input n_147;
input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_120;
input n_93;
input n_155;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_885;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_372;
wire n_341;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_583;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_317;
wire n_280;
wire n_375;
wire n_340;
wire n_708;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_170;
wire n_270;
wire n_383;
wire n_346;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_711;
wire n_228;
wire n_671;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_798;
wire n_732;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_636;
wire n_594;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_844;
wire n_245;
wire n_648;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_589;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_839;
wire n_768;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_869;
wire n_718;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_882;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_567;
wire n_548;
wire n_516;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_397;
wire n_366;
wire n_803;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_843;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_817;
wire n_744;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_288;
wire n_320;
wire n_247;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_385;
wire n_233;
wire n_414;
wire n_342;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_874;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_149),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_130),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_70),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_18),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_69),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_151),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_92),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_51),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_111),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_100),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_93),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_39),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_7),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_50),
.Y(n_176)
);

BUFx10_ASAP7_75t_L g177 ( 
.A(n_42),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_74),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_66),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_53),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_76),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_123),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_0),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_105),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_6),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_63),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_22),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_119),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_3),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_1),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_56),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_95),
.B(n_109),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_59),
.Y(n_195)
);

BUFx10_ASAP7_75t_L g196 ( 
.A(n_48),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_29),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_79),
.Y(n_198)
);

INVxp33_ASAP7_75t_SL g199 ( 
.A(n_148),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_13),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_32),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_8),
.Y(n_202)
);

INVxp67_ASAP7_75t_SL g203 ( 
.A(n_152),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_96),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_118),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_127),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_131),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_21),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_120),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_161),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_11),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_85),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_136),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_65),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_81),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_82),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_30),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_140),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_60),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_86),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_37),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_94),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_57),
.Y(n_224)
);

INVxp67_ASAP7_75t_SL g225 ( 
.A(n_83),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_43),
.Y(n_226)
);

BUFx8_ASAP7_75t_SL g227 ( 
.A(n_155),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_55),
.Y(n_228)
);

INVxp33_ASAP7_75t_SL g229 ( 
.A(n_23),
.Y(n_229)
);

NOR2xp67_ASAP7_75t_L g230 ( 
.A(n_9),
.B(n_31),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_4),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_84),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_135),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_110),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_124),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_116),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_117),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_73),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_98),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_67),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_102),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_77),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_1),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_17),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_13),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_22),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_122),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_141),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_28),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_36),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_5),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_91),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_33),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_24),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_61),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_104),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_87),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_44),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_125),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_253),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_170),
.Y(n_261)
);

NOR2x1_ASAP7_75t_L g262 ( 
.A(n_201),
.B(n_38),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_207),
.B(n_2),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_2),
.Y(n_264)
);

NOR2x1_ASAP7_75t_L g265 ( 
.A(n_183),
.B(n_40),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_227),
.B(n_41),
.Y(n_266)
);

AND2x6_ASAP7_75t_L g267 ( 
.A(n_168),
.B(n_194),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_183),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_168),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_202),
.Y(n_270)
);

XNOR2x2_ASAP7_75t_L g271 ( 
.A(n_165),
.B(n_5),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_166),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_187),
.A2(n_191),
.B1(n_229),
.B2(n_175),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_187),
.B(n_8),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_177),
.B(n_9),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_177),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_177),
.Y(n_277)
);

AND2x4_ASAP7_75t_L g278 ( 
.A(n_212),
.B(n_10),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_212),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_179),
.B(n_10),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_249),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_170),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_227),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_191),
.B(n_12),
.Y(n_284)
);

OA21x2_ASAP7_75t_L g285 ( 
.A1(n_174),
.A2(n_80),
.B(n_158),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_196),
.B(n_12),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_249),
.Y(n_287)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_254),
.Y(n_288)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_196),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_254),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_185),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_174),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_170),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_170),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_208),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_218),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_204),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_204),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_172),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_196),
.B(n_14),
.Y(n_300)
);

AND2x6_ASAP7_75t_L g301 ( 
.A(n_194),
.B(n_195),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_172),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_219),
.Y(n_303)
);

AND2x4_ASAP7_75t_L g304 ( 
.A(n_195),
.B(n_14),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_164),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_171),
.Y(n_306)
);

NOR2x1_ASAP7_75t_L g307 ( 
.A(n_173),
.B(n_45),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_229),
.B(n_15),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_172),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_219),
.B(n_15),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_222),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_222),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_206),
.B(n_16),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_206),
.B(n_16),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_172),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_200),
.Y(n_316)
);

OAI21x1_ASAP7_75t_L g317 ( 
.A1(n_228),
.A2(n_89),
.B(n_157),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_226),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_226),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_197),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_176),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_211),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_228),
.Y(n_323)
);

OAI22x1_ASAP7_75t_L g324 ( 
.A1(n_190),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_235),
.B(n_19),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_236),
.Y(n_326)
);

NAND2xp33_ASAP7_75t_L g327 ( 
.A(n_200),
.B(n_46),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_188),
.B(n_47),
.Y(n_328)
);

AND2x6_ASAP7_75t_L g329 ( 
.A(n_236),
.B(n_49),
.Y(n_329)
);

OA21x2_ASAP7_75t_L g330 ( 
.A1(n_235),
.A2(n_97),
.B(n_156),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_200),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_211),
.B(n_20),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_317),
.A2(n_240),
.B(n_238),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g334 ( 
.A(n_260),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_278),
.Y(n_335)
);

AOI21x1_ASAP7_75t_L g336 ( 
.A1(n_285),
.A2(n_240),
.B(n_238),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_278),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_261),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_289),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_261),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_261),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_282),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_282),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_288),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_320),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_282),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_283),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_275),
.Y(n_348)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_329),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_282),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_293),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_293),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_293),
.Y(n_353)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_329),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_294),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_304),
.B(n_305),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_273),
.A2(n_162),
.B1(n_163),
.B2(n_186),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_294),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_294),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_304),
.B(n_241),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_288),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_264),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_L g363 ( 
.A1(n_263),
.A2(n_199),
.B1(n_246),
.B2(n_200),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_269),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_272),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_306),
.B(n_241),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_269),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_276),
.B(n_231),
.Y(n_368)
);

INVx5_ASAP7_75t_L g369 ( 
.A(n_329),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_294),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_277),
.B(n_178),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_321),
.B(n_180),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_322),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_299),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_299),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_299),
.Y(n_376)
);

NOR2xp67_ASAP7_75t_L g377 ( 
.A(n_268),
.B(n_181),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_326),
.Y(n_378)
);

INVx5_ASAP7_75t_L g379 ( 
.A(n_329),
.Y(n_379)
);

NAND2xp33_ASAP7_75t_L g380 ( 
.A(n_329),
.B(n_267),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_268),
.B(n_189),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_272),
.Y(n_382)
);

BUFx6f_ASAP7_75t_SL g383 ( 
.A(n_267),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_326),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_299),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_281),
.B(n_286),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_291),
.B(n_245),
.Y(n_387)
);

INVxp33_ASAP7_75t_SL g388 ( 
.A(n_283),
.Y(n_388)
);

OAI22xp33_ASAP7_75t_L g389 ( 
.A1(n_266),
.A2(n_244),
.B1(n_163),
.B2(n_186),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_295),
.B(n_192),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_313),
.A2(n_162),
.B1(n_198),
.B2(n_251),
.Y(n_391)
);

INVxp33_ASAP7_75t_L g392 ( 
.A(n_300),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_292),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_302),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_302),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_296),
.B(n_167),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_297),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_302),
.Y(n_398)
);

AND2x4_ASAP7_75t_L g399 ( 
.A(n_270),
.B(n_230),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_309),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_307),
.B(n_242),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_309),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_309),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_309),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_315),
.Y(n_405)
);

AND2x2_ASAP7_75t_SL g406 ( 
.A(n_314),
.B(n_193),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_297),
.Y(n_407)
);

BUFx8_ASAP7_75t_SL g408 ( 
.A(n_274),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_315),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_332),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_315),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_315),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_284),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_298),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_318),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_L g416 ( 
.A1(n_308),
.A2(n_280),
.B1(n_301),
.B2(n_267),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_298),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_318),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_318),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_318),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_319),
.Y(n_421)
);

AND3x2_ASAP7_75t_L g422 ( 
.A(n_308),
.B(n_225),
.C(n_203),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_303),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_319),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_271),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_328),
.B(n_198),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_319),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_316),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_311),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_279),
.B(n_169),
.Y(n_430)
);

INVx11_ASAP7_75t_L g431 ( 
.A(n_267),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_312),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_362),
.B(n_280),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_364),
.Y(n_434)
);

OAI221xp5_ASAP7_75t_L g435 ( 
.A1(n_344),
.A2(n_287),
.B1(n_290),
.B2(n_325),
.C(n_310),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_380),
.A2(n_327),
.B(n_310),
.Y(n_436)
);

O2A1O1Ixp5_ASAP7_75t_L g437 ( 
.A1(n_333),
.A2(n_312),
.B(n_323),
.C(n_250),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_386),
.B(n_301),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_349),
.B(n_182),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_349),
.B(n_184),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_336),
.A2(n_330),
.B(n_285),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_406),
.A2(n_324),
.B1(n_244),
.B2(n_262),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_368),
.B(n_205),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_406),
.A2(n_323),
.B1(n_331),
.B2(n_246),
.Y(n_444)
);

OAI22xp33_ASAP7_75t_L g445 ( 
.A1(n_425),
.A2(n_331),
.B1(n_224),
.B2(n_223),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_364),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_361),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_413),
.B(n_213),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_396),
.B(n_214),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_387),
.B(n_217),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_354),
.B(n_220),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_348),
.B(n_265),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_334),
.B(n_232),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_371),
.B(n_233),
.Y(n_454)
);

NAND3xp33_ASAP7_75t_L g455 ( 
.A(n_363),
.B(n_327),
.C(n_330),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_430),
.B(n_239),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_367),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_L g458 ( 
.A1(n_335),
.A2(n_330),
.B1(n_237),
.B2(n_234),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_337),
.B(n_248),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_422),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_392),
.B(n_256),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_356),
.B(n_377),
.Y(n_462)
);

INVx8_ASAP7_75t_L g463 ( 
.A(n_383),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_426),
.A2(n_247),
.B1(n_210),
.B2(n_258),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_360),
.A2(n_209),
.B(n_216),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_365),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_367),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_378),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_378),
.B(n_215),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_384),
.B(n_221),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_384),
.B(n_252),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_384),
.B(n_255),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_382),
.Y(n_473)
);

OR2x6_ASAP7_75t_L g474 ( 
.A(n_357),
.B(n_257),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_345),
.B(n_259),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_360),
.A2(n_259),
.B(n_316),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_381),
.B(n_226),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_372),
.B(n_20),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_393),
.Y(n_479)
);

BUFx4f_ASAP7_75t_L g480 ( 
.A(n_373),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_369),
.B(n_52),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_369),
.B(n_379),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_390),
.B(n_23),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_407),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_379),
.B(n_54),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_416),
.B(n_58),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_L g487 ( 
.A1(n_397),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_487)
);

NOR2x1p5_ASAP7_75t_L g488 ( 
.A(n_347),
.B(n_27),
.Y(n_488)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_417),
.Y(n_489)
);

BUFx6f_ASAP7_75t_SL g490 ( 
.A(n_399),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_339),
.B(n_62),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_366),
.B(n_29),
.Y(n_492)
);

AND2x4_ASAP7_75t_SL g493 ( 
.A(n_410),
.B(n_30),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_401),
.A2(n_106),
.B(n_153),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_391),
.B(n_31),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_429),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_414),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_432),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_399),
.B(n_389),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_414),
.Y(n_500)
);

OAI22xp33_ASAP7_75t_L g501 ( 
.A1(n_425),
.A2(n_34),
.B1(n_35),
.B2(n_64),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_489),
.B(n_410),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_437),
.A2(n_423),
.B(n_428),
.Y(n_503)
);

OA22x2_ASAP7_75t_L g504 ( 
.A1(n_474),
.A2(n_347),
.B1(n_408),
.B2(n_388),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_463),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_447),
.A2(n_431),
.B1(n_427),
.B2(n_424),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_433),
.B(n_68),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_480),
.Y(n_508)
);

NAND2x1p5_ASAP7_75t_L g509 ( 
.A(n_480),
.B(n_341),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_452),
.B(n_498),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_434),
.Y(n_511)
);

AOI21xp33_ASAP7_75t_L g512 ( 
.A1(n_453),
.A2(n_71),
.B(n_72),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_493),
.B(n_75),
.Y(n_513)
);

A2O1A1Ixp33_ASAP7_75t_L g514 ( 
.A1(n_437),
.A2(n_421),
.B(n_420),
.C(n_419),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_500),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_441),
.A2(n_418),
.B(n_415),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_448),
.B(n_475),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_438),
.B(n_450),
.Y(n_518)
);

NOR2x1p5_ASAP7_75t_L g519 ( 
.A(n_461),
.B(n_78),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_466),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_463),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_497),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_499),
.A2(n_418),
.B1(n_415),
.B2(n_412),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_473),
.Y(n_524)
);

AO32x1_ASAP7_75t_L g525 ( 
.A1(n_444),
.A2(n_412),
.A3(n_411),
.B1(n_409),
.B2(n_338),
.Y(n_525)
);

NOR2x1p5_ASAP7_75t_L g526 ( 
.A(n_488),
.B(n_88),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_435),
.A2(n_359),
.B1(n_404),
.B2(n_403),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_462),
.B(n_90),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_458),
.A2(n_359),
.B(n_404),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_482),
.A2(n_358),
.B(n_403),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_479),
.B(n_99),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g532 ( 
.A1(n_458),
.A2(n_355),
.B(n_402),
.Y(n_532)
);

NOR2x1_ASAP7_75t_L g533 ( 
.A(n_445),
.B(n_355),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_455),
.A2(n_358),
.B(n_402),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_497),
.Y(n_535)
);

AO21x1_ASAP7_75t_L g536 ( 
.A1(n_436),
.A2(n_400),
.B(n_398),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_496),
.B(n_101),
.Y(n_537)
);

NAND3xp33_ASAP7_75t_SL g538 ( 
.A(n_442),
.B(n_400),
.C(n_398),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_469),
.Y(n_539)
);

OA22x2_ASAP7_75t_L g540 ( 
.A1(n_460),
.A2(n_395),
.B1(n_394),
.B2(n_385),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_436),
.A2(n_352),
.B(n_394),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_463),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_446),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_490),
.Y(n_544)
);

O2A1O1Ixp33_ASAP7_75t_L g545 ( 
.A1(n_445),
.A2(n_376),
.B(n_375),
.C(n_374),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_435),
.A2(n_351),
.B1(n_376),
.B2(n_375),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_443),
.B(n_103),
.Y(n_547)
);

NAND3xp33_ASAP7_75t_L g548 ( 
.A(n_478),
.B(n_346),
.C(n_370),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_470),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_484),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g551 ( 
.A1(n_487),
.A2(n_340),
.B1(n_353),
.B2(n_351),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_490),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_459),
.A2(n_350),
.B(n_342),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_457),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_454),
.B(n_107),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_449),
.B(n_108),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_465),
.B(n_112),
.Y(n_557)
);

NAND3xp33_ASAP7_75t_SL g558 ( 
.A(n_487),
.B(n_113),
.C(n_114),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_471),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_465),
.B(n_115),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_456),
.B(n_121),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_439),
.A2(n_440),
.B(n_451),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_467),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_464),
.B(n_405),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_472),
.A2(n_405),
.B1(n_343),
.B2(n_341),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_483),
.B(n_126),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_468),
.A2(n_128),
.B(n_129),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_L g568 ( 
.A1(n_477),
.A2(n_132),
.B(n_133),
.Y(n_568)
);

AO32x2_ASAP7_75t_L g569 ( 
.A1(n_476),
.A2(n_134),
.A3(n_137),
.B1(n_139),
.B2(n_142),
.Y(n_569)
);

NAND3xp33_ASAP7_75t_L g570 ( 
.A(n_476),
.B(n_143),
.C(n_144),
.Y(n_570)
);

AOI221xp5_ASAP7_75t_L g571 ( 
.A1(n_501),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.C(n_150),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_505),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_L g573 ( 
.A1(n_539),
.A2(n_491),
.B(n_492),
.Y(n_573)
);

OA21x2_ASAP7_75t_L g574 ( 
.A1(n_534),
.A2(n_536),
.B(n_541),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_502),
.B(n_501),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_520),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_L g577 ( 
.A1(n_549),
.A2(n_491),
.B(n_494),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_505),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_524),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_517),
.B(n_481),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_559),
.B(n_485),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_521),
.B(n_542),
.Y(n_582)
);

AO31x2_ASAP7_75t_L g583 ( 
.A1(n_527),
.A2(n_523),
.A3(n_514),
.B(n_565),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_521),
.B(n_542),
.Y(n_584)
);

CKINVDCx14_ASAP7_75t_R g585 ( 
.A(n_552),
.Y(n_585)
);

AO31x2_ASAP7_75t_L g586 ( 
.A1(n_557),
.A2(n_560),
.A3(n_566),
.B(n_551),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_508),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_L g588 ( 
.A1(n_503),
.A2(n_545),
.B(n_529),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_521),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_542),
.B(n_510),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_515),
.Y(n_591)
);

A2O1A1Ixp33_ASAP7_75t_L g592 ( 
.A1(n_556),
.A2(n_561),
.B(n_555),
.C(n_571),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_544),
.B(n_504),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_544),
.Y(n_594)
);

BUFx12f_ASAP7_75t_L g595 ( 
.A(n_526),
.Y(n_595)
);

AND2x4_ASAP7_75t_L g596 ( 
.A(n_513),
.B(n_519),
.Y(n_596)
);

AO32x2_ASAP7_75t_L g597 ( 
.A1(n_525),
.A2(n_506),
.A3(n_569),
.B1(n_558),
.B2(n_540),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_533),
.Y(n_598)
);

OR2x6_ASAP7_75t_L g599 ( 
.A(n_509),
.B(n_562),
.Y(n_599)
);

AND2x6_ASAP7_75t_L g600 ( 
.A(n_522),
.B(n_535),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_550),
.B(n_543),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_522),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_511),
.B(n_554),
.Y(n_603)
);

O2A1O1Ixp33_ASAP7_75t_L g604 ( 
.A1(n_564),
.A2(n_512),
.B(n_547),
.C(n_528),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_532),
.A2(n_531),
.B(n_537),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_563),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_L g607 ( 
.A1(n_548),
.A2(n_546),
.B(n_553),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_546),
.Y(n_608)
);

NOR3xp33_ASAP7_75t_L g609 ( 
.A(n_570),
.B(n_568),
.C(n_567),
.Y(n_609)
);

OAI21xp5_ASAP7_75t_L g610 ( 
.A1(n_570),
.A2(n_530),
.B(n_525),
.Y(n_610)
);

CKINVDCx11_ASAP7_75t_R g611 ( 
.A(n_569),
.Y(n_611)
);

AO21x1_ASAP7_75t_L g612 ( 
.A1(n_512),
.A2(n_486),
.B(n_507),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_502),
.A2(n_357),
.B1(n_410),
.B2(n_389),
.Y(n_613)
);

OAI21x1_ASAP7_75t_L g614 ( 
.A1(n_516),
.A2(n_441),
.B(n_534),
.Y(n_614)
);

AO31x2_ASAP7_75t_L g615 ( 
.A1(n_536),
.A2(n_527),
.A3(n_523),
.B(n_514),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_505),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_502),
.B(n_334),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_518),
.A2(n_380),
.B(n_354),
.Y(n_618)
);

OAI21x1_ASAP7_75t_L g619 ( 
.A1(n_516),
.A2(n_441),
.B(n_534),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_520),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_502),
.B(n_334),
.Y(n_621)
);

A2O1A1Ixp33_ASAP7_75t_L g622 ( 
.A1(n_539),
.A2(n_559),
.B(n_549),
.C(n_433),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_505),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_518),
.A2(n_380),
.B(n_354),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_L g625 ( 
.A1(n_539),
.A2(n_437),
.B(n_455),
.Y(n_625)
);

A2O1A1Ixp33_ASAP7_75t_L g626 ( 
.A1(n_539),
.A2(n_559),
.B(n_549),
.C(n_433),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_502),
.B(n_334),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_L g628 ( 
.A1(n_539),
.A2(n_437),
.B(n_455),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_505),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_502),
.B(n_334),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_502),
.B(n_334),
.Y(n_631)
);

OAI21x1_ASAP7_75t_L g632 ( 
.A1(n_516),
.A2(n_441),
.B(n_534),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_520),
.Y(n_633)
);

NAND3x1_ASAP7_75t_L g634 ( 
.A(n_502),
.B(n_442),
.C(n_495),
.Y(n_634)
);

NOR2xp67_ASAP7_75t_L g635 ( 
.A(n_508),
.B(n_357),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_518),
.A2(n_380),
.B(n_354),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_520),
.Y(n_637)
);

NOR4xp25_ASAP7_75t_L g638 ( 
.A(n_538),
.B(n_501),
.C(n_487),
.D(n_499),
.Y(n_638)
);

AO31x2_ASAP7_75t_L g639 ( 
.A1(n_536),
.A2(n_527),
.A3(n_523),
.B(n_514),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_SL g640 ( 
.A(n_508),
.B(n_357),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_520),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_505),
.B(n_521),
.Y(n_642)
);

OAI21xp5_ASAP7_75t_SL g643 ( 
.A1(n_502),
.A2(n_389),
.B(n_357),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_502),
.A2(n_357),
.B1(n_410),
.B2(n_389),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_502),
.B(n_334),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_502),
.B(n_334),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_520),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_L g648 ( 
.A1(n_539),
.A2(n_437),
.B(n_455),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_502),
.B(n_334),
.Y(n_649)
);

OAI21x1_ASAP7_75t_L g650 ( 
.A1(n_516),
.A2(n_441),
.B(n_534),
.Y(n_650)
);

OAI22x1_ASAP7_75t_L g651 ( 
.A1(n_526),
.A2(n_391),
.B1(n_442),
.B2(n_488),
.Y(n_651)
);

AO21x2_ASAP7_75t_L g652 ( 
.A1(n_536),
.A2(n_441),
.B(n_333),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_520),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_585),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_652),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_579),
.Y(n_656)
);

INVx5_ASAP7_75t_L g657 ( 
.A(n_578),
.Y(n_657)
);

OA21x2_ASAP7_75t_L g658 ( 
.A1(n_610),
.A2(n_632),
.B(n_650),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_578),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_620),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_637),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_643),
.B(n_575),
.Y(n_662)
);

INVx6_ASAP7_75t_L g663 ( 
.A(n_578),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_627),
.B(n_617),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_576),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_633),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_621),
.B(n_630),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_574),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_631),
.B(n_645),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_629),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_584),
.Y(n_671)
);

INVxp67_ASAP7_75t_L g672 ( 
.A(n_646),
.Y(n_672)
);

AO21x2_ASAP7_75t_L g673 ( 
.A1(n_588),
.A2(n_628),
.B(n_625),
.Y(n_673)
);

AO21x2_ASAP7_75t_L g674 ( 
.A1(n_648),
.A2(n_605),
.B(n_609),
.Y(n_674)
);

NAND3xp33_ASAP7_75t_L g675 ( 
.A(n_640),
.B(n_613),
.C(n_644),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_649),
.B(n_635),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_595),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_641),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_604),
.A2(n_592),
.B(n_577),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_647),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_591),
.B(n_590),
.Y(n_681)
);

NAND2x1p5_ASAP7_75t_L g682 ( 
.A(n_584),
.B(n_642),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_653),
.Y(n_683)
);

OA21x2_ASAP7_75t_L g684 ( 
.A1(n_612),
.A2(n_608),
.B(n_598),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_618),
.A2(n_636),
.B(n_624),
.Y(n_685)
);

NOR2x1_ASAP7_75t_SL g686 ( 
.A(n_616),
.B(n_582),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_603),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_642),
.B(n_590),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_634),
.B(n_638),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_572),
.B(n_623),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_601),
.Y(n_691)
);

OA21x2_ASAP7_75t_L g692 ( 
.A1(n_573),
.A2(n_581),
.B(n_580),
.Y(n_692)
);

CKINVDCx11_ASAP7_75t_R g693 ( 
.A(n_587),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_651),
.B(n_596),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_589),
.Y(n_695)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_594),
.Y(n_696)
);

INVx1_ASAP7_75t_SL g697 ( 
.A(n_593),
.Y(n_697)
);

OAI21x1_ASAP7_75t_L g698 ( 
.A1(n_606),
.A2(n_602),
.B(n_615),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_599),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_615),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_600),
.B(n_583),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_611),
.A2(n_600),
.B1(n_597),
.B2(n_639),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_583),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_597),
.B(n_586),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_585),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_575),
.B(n_627),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_579),
.Y(n_707)
);

OR2x6_ASAP7_75t_L g708 ( 
.A(n_595),
.B(n_505),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_579),
.Y(n_709)
);

AO21x2_ASAP7_75t_L g710 ( 
.A1(n_610),
.A2(n_588),
.B(n_607),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_575),
.B(n_627),
.Y(n_711)
);

OA21x2_ASAP7_75t_L g712 ( 
.A1(n_610),
.A2(n_619),
.B(n_614),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_584),
.Y(n_713)
);

NOR2xp67_ASAP7_75t_L g714 ( 
.A(n_595),
.B(n_508),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_622),
.B(n_626),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_579),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_575),
.B(n_627),
.Y(n_717)
);

OR2x2_ASAP7_75t_L g718 ( 
.A(n_689),
.B(n_683),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_680),
.Y(n_719)
);

BUFx2_ASAP7_75t_L g720 ( 
.A(n_701),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_668),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_667),
.B(n_669),
.Y(n_722)
);

OAI21xp5_ASAP7_75t_L g723 ( 
.A1(n_679),
.A2(n_676),
.B(n_675),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_680),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_683),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_664),
.B(n_662),
.Y(n_726)
);

BUFx2_ASAP7_75t_L g727 ( 
.A(n_701),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_701),
.B(n_699),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_655),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_665),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_662),
.B(n_715),
.Y(n_731)
);

INVx1_ASAP7_75t_SL g732 ( 
.A(n_696),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_666),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_694),
.B(n_672),
.Y(n_734)
);

HB1xp67_ASAP7_75t_L g735 ( 
.A(n_681),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_715),
.B(n_687),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_657),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_678),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_672),
.Y(n_739)
);

HB1xp67_ASAP7_75t_L g740 ( 
.A(n_656),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_684),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_684),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_657),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_717),
.B(n_706),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_715),
.A2(n_676),
.B1(n_711),
.B2(n_697),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_684),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_693),
.Y(n_747)
);

INVx1_ASAP7_75t_SL g748 ( 
.A(n_693),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_698),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_657),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_659),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_660),
.B(n_709),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_661),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_705),
.Y(n_754)
);

NOR2x1_ASAP7_75t_SL g755 ( 
.A(n_657),
.B(n_670),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_692),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_707),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_716),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_670),
.Y(n_759)
);

INVx1_ASAP7_75t_SL g760 ( 
.A(n_654),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_700),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_703),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_761),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_731),
.B(n_704),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_731),
.B(n_719),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_725),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_759),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_725),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_724),
.B(n_736),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_718),
.B(n_710),
.Y(n_770)
);

OR2x2_ASAP7_75t_L g771 ( 
.A(n_718),
.B(n_710),
.Y(n_771)
);

BUFx2_ASAP7_75t_L g772 ( 
.A(n_720),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_721),
.B(n_673),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_722),
.B(n_705),
.Y(n_774)
);

BUFx2_ASAP7_75t_L g775 ( 
.A(n_720),
.Y(n_775)
);

OR2x2_ASAP7_75t_L g776 ( 
.A(n_726),
.B(n_762),
.Y(n_776)
);

OAI221xp5_ASAP7_75t_L g777 ( 
.A1(n_723),
.A2(n_691),
.B1(n_702),
.B2(n_714),
.C(n_685),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_756),
.B(n_658),
.Y(n_778)
);

HB1xp67_ASAP7_75t_L g779 ( 
.A(n_751),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_729),
.Y(n_780)
);

BUFx2_ASAP7_75t_L g781 ( 
.A(n_727),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_728),
.B(n_712),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_752),
.B(n_712),
.Y(n_783)
);

OR2x2_ASAP7_75t_L g784 ( 
.A(n_728),
.B(n_712),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_730),
.B(n_674),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_747),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_779),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_780),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_765),
.B(n_730),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_774),
.B(n_748),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_782),
.B(n_741),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_763),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_765),
.B(n_733),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_763),
.Y(n_794)
);

BUFx2_ASAP7_75t_L g795 ( 
.A(n_772),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_764),
.B(n_741),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_782),
.B(n_742),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_764),
.B(n_746),
.Y(n_798)
);

INVx1_ASAP7_75t_SL g799 ( 
.A(n_772),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_779),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_770),
.B(n_746),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_776),
.B(n_769),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_784),
.B(n_749),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_783),
.B(n_769),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_787),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_804),
.B(n_783),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_796),
.B(n_776),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_792),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_804),
.B(n_773),
.Y(n_809)
);

NOR2x1_ASAP7_75t_L g810 ( 
.A(n_790),
.B(n_750),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_794),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_796),
.B(n_773),
.Y(n_812)
);

INVx6_ASAP7_75t_L g813 ( 
.A(n_803),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_798),
.B(n_773),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_798),
.B(n_766),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_802),
.B(n_766),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_791),
.B(n_778),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_788),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_791),
.B(n_778),
.Y(n_819)
);

OR2x2_ASAP7_75t_L g820 ( 
.A(n_801),
.B(n_770),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_801),
.B(n_771),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_791),
.B(n_778),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_805),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_818),
.Y(n_824)
);

NAND3xp33_ASAP7_75t_L g825 ( 
.A(n_810),
.B(n_771),
.C(n_800),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_806),
.B(n_799),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_806),
.B(n_791),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_808),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_SL g829 ( 
.A1(n_813),
.A2(n_795),
.B1(n_775),
.B2(n_781),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_808),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_817),
.B(n_797),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_815),
.B(n_789),
.Y(n_832)
);

OR2x2_ASAP7_75t_L g833 ( 
.A(n_807),
.B(n_800),
.Y(n_833)
);

NAND4xp25_ASAP7_75t_L g834 ( 
.A(n_816),
.B(n_745),
.C(n_734),
.D(n_777),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_818),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_811),
.Y(n_836)
);

AOI31xp33_ASAP7_75t_L g837 ( 
.A1(n_825),
.A2(n_829),
.A3(n_760),
.B(n_823),
.Y(n_837)
);

AOI322xp5_ASAP7_75t_L g838 ( 
.A1(n_827),
.A2(n_809),
.A3(n_814),
.B1(n_812),
.B2(n_819),
.C1(n_817),
.C2(n_822),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_828),
.Y(n_839)
);

NOR3xp33_ASAP7_75t_L g840 ( 
.A(n_834),
.B(n_732),
.C(n_777),
.Y(n_840)
);

OR2x2_ASAP7_75t_L g841 ( 
.A(n_832),
.B(n_820),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_824),
.Y(n_842)
);

OAI31xp33_ASAP7_75t_L g843 ( 
.A1(n_831),
.A2(n_795),
.A3(n_739),
.B(n_820),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_830),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_836),
.Y(n_845)
);

NAND3xp33_ASAP7_75t_L g846 ( 
.A(n_829),
.B(n_821),
.C(n_785),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_833),
.Y(n_847)
);

A2O1A1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_831),
.A2(n_822),
.B(n_819),
.C(n_793),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_838),
.B(n_809),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_848),
.A2(n_831),
.B1(n_813),
.B2(n_827),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_843),
.B(n_812),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_848),
.A2(n_837),
.B1(n_846),
.B2(n_813),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_847),
.B(n_814),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_839),
.Y(n_854)
);

OAI22xp33_ASAP7_75t_L g855 ( 
.A1(n_850),
.A2(n_813),
.B1(n_841),
.B2(n_821),
.Y(n_855)
);

A2O1A1Ixp33_ASAP7_75t_L g856 ( 
.A1(n_852),
.A2(n_840),
.B(n_826),
.C(n_844),
.Y(n_856)
);

NAND3xp33_ASAP7_75t_L g857 ( 
.A(n_849),
.B(n_840),
.C(n_845),
.Y(n_857)
);

OAI211xp5_ASAP7_75t_L g858 ( 
.A1(n_856),
.A2(n_851),
.B(n_677),
.C(n_786),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_857),
.B(n_854),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_859),
.B(n_855),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_858),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_861),
.Y(n_862)
);

OR2x2_ASAP7_75t_L g863 ( 
.A(n_860),
.B(n_853),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_862),
.Y(n_864)
);

XNOR2xp5_ASAP7_75t_L g865 ( 
.A(n_863),
.B(n_754),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_865),
.B(n_842),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_864),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_865),
.B(n_824),
.Y(n_868)
);

NOR4xp25_ASAP7_75t_L g869 ( 
.A(n_867),
.B(n_677),
.C(n_708),
.D(n_738),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_866),
.A2(n_708),
.B(n_744),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_SL g871 ( 
.A1(n_868),
.A2(n_708),
.B1(n_750),
.B2(n_743),
.Y(n_871)
);

OA21x2_ASAP7_75t_L g872 ( 
.A1(n_866),
.A2(n_695),
.B(n_733),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_866),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_873),
.A2(n_743),
.B1(n_737),
.B2(n_750),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_871),
.A2(n_737),
.B1(n_835),
.B2(n_738),
.Y(n_875)
);

NAND3x1_ASAP7_75t_L g876 ( 
.A(n_870),
.B(n_752),
.C(n_758),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_869),
.A2(n_690),
.B(n_753),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_872),
.A2(n_835),
.B1(n_768),
.B2(n_767),
.Y(n_878)
);

OAI21x1_ASAP7_75t_L g879 ( 
.A1(n_873),
.A2(n_682),
.B(n_758),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_877),
.A2(n_740),
.B(n_686),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_879),
.A2(n_755),
.B(n_671),
.Y(n_881)
);

AOI222xp33_ASAP7_75t_L g882 ( 
.A1(n_875),
.A2(n_878),
.B1(n_876),
.B2(n_874),
.C1(n_757),
.C2(n_735),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_882),
.B(n_880),
.Y(n_883)
);

OR2x6_ASAP7_75t_L g884 ( 
.A(n_883),
.B(n_881),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_884),
.A2(n_663),
.B1(n_713),
.B2(n_688),
.Y(n_885)
);


endmodule