module real_jpeg_17618_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AND2x4_ASAP7_75t_L g15 ( 
.A(n_0),
.B(n_16),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_0),
.B(n_45),
.Y(n_44)
);

AND2x4_ASAP7_75t_SL g52 ( 
.A(n_0),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_0),
.B(n_42),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_0),
.B(n_75),
.Y(n_74)
);

AND2x4_ASAP7_75t_L g97 ( 
.A(n_0),
.B(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_1),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_4),
.B(n_21),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_4),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_4),
.B(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g13 ( 
.A(n_6),
.B(n_14),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_6),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_6),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_6),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_6),
.B(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_7),
.Y(n_99)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_85),
.Y(n_9)
);

AOI21xp5_ASAP7_75t_L g10 ( 
.A1(n_11),
.A2(n_66),
.B(n_84),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_31),
.Y(n_11)
);

NOR2xp67_ASAP7_75t_L g84 ( 
.A(n_12),
.B(n_31),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_SL g12 ( 
.A1(n_13),
.A2(n_15),
.B(n_19),
.C(n_30),
.Y(n_12)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_15),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_13),
.A2(n_15),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_13),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_13),
.A2(n_81),
.B1(n_109),
.B2(n_111),
.Y(n_108)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_15),
.Y(n_82)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_18),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_19),
.B(n_80),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_20),
.Y(n_28)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

INVxp33_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NOR2x1_ASAP7_75t_R g72 ( 
.A(n_24),
.B(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_49),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_32),
.B(n_59),
.C(n_64),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_37),
.B1(n_47),
.B2(n_48),
.Y(n_32)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_39),
.B(n_43),
.C(n_47),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_59),
.B1(n_64),
.B2(n_65),
.Y(n_49)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_58),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_52),
.A2(n_74),
.B(n_110),
.Y(n_109)
);

NAND2x1p5_ASAP7_75t_L g110 ( 
.A(n_52),
.B(n_74),
.Y(n_110)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_54),
.B(n_60),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_54),
.A2(n_59),
.B(n_60),
.Y(n_69)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_79),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_78),
.B(n_83),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_72),
.B(n_77),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_70),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_113),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NOR2xp67_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_112),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_112),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_106),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_104),
.B2(n_105),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_95),
.B1(n_96),
.B2(n_103),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_92),
.Y(n_103)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_109),
.Y(n_111)
);


endmodule