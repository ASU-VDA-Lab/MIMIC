module fake_jpeg_18104_n_161 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_161);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_161;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_45),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_16),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_9),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_4),
.Y(n_68)
);

BUFx24_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_7),
.B(n_2),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx4f_ASAP7_75t_SL g73 ( 
.A(n_41),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_11),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_13),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_79),
.Y(n_88)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_0),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_57),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_83),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_78),
.A2(n_75),
.B1(n_68),
.B2(n_63),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_89),
.A2(n_77),
.B1(n_69),
.B2(n_67),
.Y(n_96)
);

AOI21xp33_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_70),
.B(n_66),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_90),
.B(n_74),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_67),
.B1(n_75),
.B2(n_55),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_93),
.A2(n_51),
.B1(n_68),
.B2(n_50),
.Y(n_101)
);

FAx1_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_69),
.CI(n_64),
.CON(n_95),
.SN(n_95)
);

AOI21xp33_ASAP7_75t_L g107 ( 
.A1(n_95),
.A2(n_98),
.B(n_99),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_101),
.B1(n_106),
.B2(n_91),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_87),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_48),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_82),
.B(n_51),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_105),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_85),
.A2(n_49),
.B1(n_73),
.B2(n_61),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_100),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_109),
.B(n_110),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_106),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_98),
.A2(n_92),
.B1(n_85),
.B2(n_86),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_116),
.B1(n_120),
.B2(n_5),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_113),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_118),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_92),
.B1(n_84),
.B2(n_72),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_65),
.Y(n_118)
);

OAI32xp33_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_73),
.A3(n_58),
.B1(n_71),
.B2(n_56),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_121),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_97),
.A2(n_72),
.B1(n_23),
.B2(n_24),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_0),
.Y(n_121)
);

FAx1_ASAP7_75t_SL g123 ( 
.A(n_107),
.B(n_62),
.CI(n_53),
.CON(n_123),
.SN(n_123)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_124),
.Y(n_137)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_52),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_129),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_127),
.A2(n_133),
.B1(n_116),
.B2(n_112),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_120),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_119),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_130),
.A2(n_134),
.B(n_10),
.Y(n_136)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_132),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_25),
.C(n_43),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_112),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_134)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_122),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_139)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_141),
.B(n_142),
.Y(n_146)
);

OAI22x1_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_125),
.B1(n_133),
.B2(n_123),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_126),
.A2(n_30),
.B(n_17),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_145),
.A2(n_142),
.B1(n_138),
.B2(n_137),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_148),
.B(n_149),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_140),
.C(n_143),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_140),
.C(n_147),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_132),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_144),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_144),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_134),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_33),
.C(n_18),
.Y(n_157)
);

NAND3xp33_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_35),
.C(n_21),
.Y(n_158)
);

AO22x1_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_36),
.B1(n_22),
.B2(n_26),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_27),
.B(n_38),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_160),
.B(n_46),
.Y(n_161)
);


endmodule