module fake_ariane_3057_n_2180 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2180);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2180;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2116;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_851;
wire n_444;
wire n_355;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2168;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1769;
wire n_1632;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_2016;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2143;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_2173;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_928;
wire n_253;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g219 ( 
.A(n_172),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_167),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_9),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_50),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_178),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_155),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_137),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_154),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_139),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_152),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_78),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_49),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_210),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_74),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_101),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_22),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_83),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_186),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_4),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_73),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_34),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_74),
.Y(n_240)
);

BUFx5_ASAP7_75t_L g241 ( 
.A(n_53),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_148),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_41),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_13),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_176),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_14),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_19),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_142),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_6),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_109),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_121),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_153),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_128),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_204),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_134),
.Y(n_255)
);

BUFx5_ASAP7_75t_L g256 ( 
.A(n_47),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_3),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_15),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_0),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_27),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_183),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_76),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_34),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_59),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_174),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_36),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_151),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_119),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_161),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_12),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_27),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_67),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_111),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_45),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_70),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_40),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_38),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_84),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_48),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_28),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_170),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_146),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_72),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_19),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_37),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_188),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_107),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_24),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_182),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_55),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_2),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_118),
.Y(n_292)
);

BUFx8_ASAP7_75t_SL g293 ( 
.A(n_98),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_81),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_3),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_23),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_66),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_94),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_129),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_145),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_215),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_91),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_42),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_76),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_217),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_32),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_25),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_163),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_212),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_166),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_140),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_201),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_124),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_45),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_190),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_43),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_22),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_12),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_196),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_56),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_115),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_30),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_132),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_103),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_189),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_90),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_73),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_16),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_162),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_47),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_15),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_112),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_149),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_102),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_86),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_14),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_20),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_58),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g339 ( 
.A(n_10),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_58),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_184),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_164),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_136),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_13),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_122),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_65),
.Y(n_346)
);

INVx2_ASAP7_75t_SL g347 ( 
.A(n_71),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_33),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_41),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_31),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_20),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_9),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_198),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_216),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_67),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_179),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_100),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_2),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_193),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_92),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_56),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_33),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_191),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_48),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_80),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_70),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_53),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_59),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_150),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_123),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_52),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_141),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_63),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_40),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_159),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_72),
.Y(n_376)
);

INVxp33_ASAP7_75t_SL g377 ( 
.A(n_116),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_23),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_75),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_105),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_6),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_17),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_29),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_65),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_99),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_88),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_205),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_87),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_62),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_165),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_31),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_95),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_57),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_173),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_218),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_187),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_43),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_80),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_89),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_209),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_213),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_177),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_50),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_69),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_175),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_8),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_71),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_106),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_171),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_44),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_25),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_62),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_52),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_211),
.Y(n_414)
);

CKINVDCx14_ASAP7_75t_R g415 ( 
.A(n_10),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_5),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_16),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_125),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_54),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_54),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_36),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_55),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_42),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_120),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_68),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_126),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_97),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_108),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_79),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_0),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_293),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_339),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_251),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_241),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_415),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_241),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_241),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_289),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_241),
.Y(n_439)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_393),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_312),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_313),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_241),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_387),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_241),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_241),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_395),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_241),
.Y(n_448)
);

INVxp67_ASAP7_75t_SL g449 ( 
.A(n_393),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_241),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_256),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_256),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_409),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_256),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_275),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_270),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_270),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_275),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_419),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_256),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_392),
.B(n_1),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_256),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_256),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_256),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_256),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_250),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_256),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_221),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_419),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_234),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_393),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_316),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_283),
.Y(n_473)
);

INVxp33_ASAP7_75t_SL g474 ( 
.A(n_283),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_219),
.Y(n_475)
);

INVxp67_ASAP7_75t_SL g476 ( 
.A(n_271),
.Y(n_476)
);

INVxp33_ASAP7_75t_SL g477 ( 
.A(n_366),
.Y(n_477)
);

INVxp67_ASAP7_75t_SL g478 ( 
.A(n_271),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_222),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_368),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_383),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_219),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_235),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_235),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_236),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_230),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_236),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_366),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_237),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_245),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_238),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_245),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_239),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_392),
.B(n_1),
.Y(n_494)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_307),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_240),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_403),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_421),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_250),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_302),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_265),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_265),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_399),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_282),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_282),
.Y(n_505)
);

INVxp67_ASAP7_75t_SL g506 ( 
.A(n_307),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_229),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_247),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_286),
.B(n_4),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_286),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_229),
.Y(n_511)
);

NOR2xp67_ASAP7_75t_L g512 ( 
.A(n_262),
.B(n_5),
.Y(n_512)
);

INVxp67_ASAP7_75t_SL g513 ( 
.A(n_407),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_300),
.B(n_7),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_300),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_257),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_258),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_259),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_260),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_362),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_315),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_263),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_315),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_321),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_243),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_264),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_302),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_266),
.Y(n_528)
);

CKINVDCx16_ASAP7_75t_R g529 ( 
.A(n_375),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_321),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_272),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_326),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_274),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_326),
.B(n_7),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_329),
.Y(n_535)
);

INVxp33_ASAP7_75t_L g536 ( 
.A(n_243),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_407),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_329),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_362),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_277),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_280),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_341),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_341),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_342),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_362),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_434),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_475),
.B(n_417),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_434),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_436),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_436),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_503),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_437),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_437),
.Y(n_553)
);

INVx5_ASAP7_75t_L g554 ( 
.A(n_520),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_475),
.B(n_417),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_439),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_439),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_443),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_482),
.B(n_244),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_440),
.B(n_342),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_545),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_443),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_482),
.B(n_262),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_545),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_537),
.Y(n_565)
);

INVx6_ASAP7_75t_L g566 ( 
.A(n_503),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_455),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_449),
.B(n_353),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_471),
.B(n_353),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_445),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_445),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_473),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_446),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_446),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_448),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_520),
.Y(n_576)
);

OAI21x1_ASAP7_75t_L g577 ( 
.A1(n_448),
.A2(n_356),
.B(n_354),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_483),
.B(n_244),
.Y(n_578)
);

INVx5_ASAP7_75t_L g579 ( 
.A(n_539),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_483),
.B(n_288),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_450),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_471),
.B(n_354),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_450),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_451),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_451),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_452),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_452),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_454),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_454),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_460),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_460),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_462),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_462),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_539),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_463),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_484),
.B(n_288),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_463),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_484),
.B(n_347),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_485),
.B(n_246),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_464),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_464),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_465),
.Y(n_602)
);

AND2x6_ASAP7_75t_L g603 ( 
.A(n_544),
.B(n_356),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_465),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_485),
.B(n_246),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_467),
.Y(n_606)
);

BUFx8_ASAP7_75t_L g607 ( 
.A(n_456),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_487),
.B(n_359),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_467),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_487),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_490),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_490),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_492),
.Y(n_613)
);

NAND2xp33_ASAP7_75t_L g614 ( 
.A(n_509),
.B(n_362),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_476),
.B(n_377),
.Y(n_615)
);

AND2x6_ASAP7_75t_L g616 ( 
.A(n_492),
.B(n_356),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_501),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_501),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_502),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_502),
.B(n_359),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_504),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_504),
.B(n_249),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_505),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_505),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_510),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_510),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_474),
.A2(n_328),
.B1(n_330),
.B2(n_232),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_515),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_515),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_521),
.B(n_347),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_521),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_523),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_523),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_524),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_524),
.B(n_363),
.Y(n_635)
);

OR2x6_ASAP7_75t_L g636 ( 
.A(n_563),
.B(n_461),
.Y(n_636)
);

BUFx10_ASAP7_75t_L g637 ( 
.A(n_615),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_566),
.Y(n_638)
);

BUFx10_ASAP7_75t_L g639 ( 
.A(n_615),
.Y(n_639)
);

INVxp33_ASAP7_75t_L g640 ( 
.A(n_567),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_546),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_551),
.B(n_624),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_603),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_627),
.A2(n_477),
.B1(n_494),
.B2(n_456),
.Y(n_644)
);

INVx1_ASAP7_75t_SL g645 ( 
.A(n_567),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_546),
.Y(n_646)
);

OR2x6_ASAP7_75t_L g647 ( 
.A(n_563),
.B(n_512),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_546),
.Y(n_648)
);

AND2x6_ASAP7_75t_L g649 ( 
.A(n_599),
.B(n_363),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_551),
.B(n_466),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_551),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_610),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_572),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_603),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_624),
.B(n_466),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_610),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_566),
.B(n_529),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_546),
.Y(n_658)
);

AO22x2_ASAP7_75t_L g659 ( 
.A1(n_627),
.A2(n_457),
.B1(n_534),
.B2(n_514),
.Y(n_659)
);

OR2x6_ASAP7_75t_L g660 ( 
.A(n_563),
.B(n_507),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_617),
.B(n_529),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_548),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_611),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_566),
.Y(n_664)
);

BUFx6f_ASAP7_75t_SL g665 ( 
.A(n_563),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_617),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_565),
.A2(n_486),
.B1(n_489),
.B2(n_479),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_585),
.Y(n_668)
);

BUFx10_ASAP7_75t_L g669 ( 
.A(n_566),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_548),
.Y(n_670)
);

INVx5_ASAP7_75t_L g671 ( 
.A(n_603),
.Y(n_671)
);

OR2x6_ASAP7_75t_L g672 ( 
.A(n_563),
.B(n_511),
.Y(n_672)
);

INVx5_ASAP7_75t_L g673 ( 
.A(n_603),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_611),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_617),
.B(n_618),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_612),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_598),
.A2(n_488),
.B1(n_536),
.B2(n_532),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_566),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_548),
.Y(n_679)
);

INVx4_ASAP7_75t_L g680 ( 
.A(n_603),
.Y(n_680)
);

OR2x6_ASAP7_75t_L g681 ( 
.A(n_598),
.B(n_525),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_585),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_548),
.Y(n_683)
);

INVx4_ASAP7_75t_L g684 ( 
.A(n_603),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_624),
.B(n_530),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_566),
.B(n_491),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_549),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_565),
.A2(n_496),
.B1(n_508),
.B2(n_493),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_549),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_572),
.B(n_458),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_549),
.Y(n_691)
);

OAI22xp5_ASAP7_75t_L g692 ( 
.A1(n_560),
.A2(n_469),
.B1(n_459),
.B2(n_285),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_L g693 ( 
.A1(n_560),
.A2(n_290),
.B1(n_294),
.B2(n_284),
.Y(n_693)
);

INVx5_ASAP7_75t_L g694 ( 
.A(n_603),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_585),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_549),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_612),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_552),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_585),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_552),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_598),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_624),
.B(n_530),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_619),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_619),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_553),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_617),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_624),
.B(n_532),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_568),
.B(n_535),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_628),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_568),
.B(n_433),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_628),
.B(n_535),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_598),
.B(n_478),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_552),
.Y(n_713)
);

AND2x2_ASAP7_75t_SL g714 ( 
.A(n_614),
.B(n_223),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_631),
.B(n_538),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_617),
.B(n_516),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_631),
.B(n_517),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_634),
.B(n_538),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_617),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_559),
.B(n_495),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_552),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_634),
.Y(n_722)
);

OAI22xp33_ASAP7_75t_SL g723 ( 
.A1(n_608),
.A2(n_444),
.B1(n_447),
.B2(n_438),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_588),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_617),
.B(n_518),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_598),
.B(n_542),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_613),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_588),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_613),
.Y(n_729)
);

AO21x2_ASAP7_75t_L g730 ( 
.A1(n_577),
.A2(n_372),
.B(n_370),
.Y(n_730)
);

AND2x6_ASAP7_75t_L g731 ( 
.A(n_599),
.B(n_370),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_588),
.Y(n_732)
);

NAND2xp33_ASAP7_75t_L g733 ( 
.A(n_603),
.B(n_362),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_630),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_559),
.B(n_506),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_559),
.B(n_513),
.Y(n_736)
);

BUFx2_ASAP7_75t_L g737 ( 
.A(n_607),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_613),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_621),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_630),
.B(n_542),
.Y(n_740)
);

OR2x6_ASAP7_75t_L g741 ( 
.A(n_630),
.B(n_543),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_621),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_588),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_621),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_630),
.A2(n_296),
.B1(n_297),
.B2(n_295),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_621),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_630),
.B(n_543),
.Y(n_747)
);

INVx5_ASAP7_75t_L g748 ( 
.A(n_603),
.Y(n_748)
);

OR2x6_ASAP7_75t_L g749 ( 
.A(n_599),
.B(n_544),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_623),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_623),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_623),
.Y(n_752)
);

AND2x6_ASAP7_75t_L g753 ( 
.A(n_605),
.B(n_372),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_623),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_617),
.B(n_519),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_608),
.A2(n_314),
.B1(n_317),
.B2(n_306),
.Y(n_756)
);

INVx4_ASAP7_75t_SL g757 ( 
.A(n_603),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_625),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_553),
.B(n_522),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_556),
.B(n_526),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_547),
.A2(n_276),
.B1(n_279),
.B2(n_249),
.Y(n_761)
);

INVx5_ASAP7_75t_L g762 ( 
.A(n_616),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_618),
.B(n_528),
.Y(n_763)
);

NAND2x1p5_ASAP7_75t_L g764 ( 
.A(n_578),
.B(n_269),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_556),
.B(n_531),
.Y(n_765)
);

INVx1_ASAP7_75t_SL g766 ( 
.A(n_555),
.Y(n_766)
);

BUFx2_ASAP7_75t_L g767 ( 
.A(n_607),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_607),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_625),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_625),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_562),
.B(n_533),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_625),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_618),
.B(n_540),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_591),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_591),
.Y(n_775)
);

INVx6_ASAP7_75t_L g776 ( 
.A(n_547),
.Y(n_776)
);

NOR3xp33_ASAP7_75t_L g777 ( 
.A(n_569),
.B(n_541),
.C(n_384),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_591),
.Y(n_778)
);

AND2x6_ASAP7_75t_L g779 ( 
.A(n_605),
.B(n_380),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_591),
.Y(n_780)
);

BUFx10_ASAP7_75t_L g781 ( 
.A(n_547),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_600),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_618),
.Y(n_783)
);

INVx1_ASAP7_75t_SL g784 ( 
.A(n_555),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_562),
.B(n_360),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_618),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_571),
.B(n_432),
.Y(n_787)
);

NAND2xp33_ASAP7_75t_L g788 ( 
.A(n_616),
.B(n_420),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_600),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_618),
.B(n_380),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_607),
.Y(n_791)
);

BUFx3_ASAP7_75t_L g792 ( 
.A(n_571),
.Y(n_792)
);

OAI21xp5_ASAP7_75t_L g793 ( 
.A1(n_641),
.A2(n_577),
.B(n_574),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_765),
.B(n_557),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_653),
.B(n_499),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_643),
.B(n_557),
.Y(n_796)
);

NAND2xp33_ASAP7_75t_L g797 ( 
.A(n_649),
.B(n_616),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_645),
.B(n_766),
.Y(n_798)
);

AO21x2_ASAP7_75t_L g799 ( 
.A1(n_716),
.A2(n_755),
.B(n_725),
.Y(n_799)
);

INVxp67_ASAP7_75t_L g800 ( 
.A(n_787),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_717),
.B(n_557),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_638),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_708),
.B(n_557),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_701),
.B(n_557),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_640),
.B(n_500),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_SL g806 ( 
.A1(n_659),
.A2(n_607),
.B1(n_527),
.B2(n_442),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_705),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_782),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_705),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_643),
.B(n_597),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_784),
.B(n_555),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_701),
.B(n_597),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_643),
.B(n_597),
.Y(n_813)
);

NAND2x1_ASAP7_75t_L g814 ( 
.A(n_654),
.B(n_616),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_734),
.B(n_597),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_654),
.B(n_597),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_734),
.B(n_712),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_712),
.B(n_547),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_792),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_792),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_712),
.B(n_547),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_759),
.B(n_605),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_654),
.B(n_573),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_782),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_760),
.B(n_622),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_652),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_771),
.B(n_622),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_640),
.B(n_441),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_680),
.B(n_573),
.Y(n_829)
);

OAI21xp5_ASAP7_75t_L g830 ( 
.A1(n_641),
.A2(n_577),
.B(n_575),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_655),
.B(n_622),
.Y(n_831)
);

A2O1A1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_726),
.A2(n_635),
.B(n_620),
.C(n_582),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_649),
.B(n_574),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_710),
.B(n_453),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_710),
.B(n_435),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_695),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_789),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_649),
.A2(n_616),
.B1(n_614),
.B2(n_602),
.Y(n_838)
);

NAND3xp33_ASAP7_75t_L g839 ( 
.A(n_644),
.B(n_431),
.C(n_618),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_649),
.B(n_575),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_690),
.B(n_578),
.Y(n_841)
);

NAND2xp33_ASAP7_75t_L g842 ( 
.A(n_649),
.B(n_616),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_720),
.B(n_578),
.Y(n_843)
);

INVx2_ASAP7_75t_SL g844 ( 
.A(n_720),
.Y(n_844)
);

AND2x2_ASAP7_75t_SL g845 ( 
.A(n_737),
.B(n_620),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_656),
.Y(n_846)
);

INVxp67_ASAP7_75t_L g847 ( 
.A(n_735),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_680),
.B(n_581),
.Y(n_848)
);

INVx4_ASAP7_75t_L g849 ( 
.A(n_680),
.Y(n_849)
);

INVx8_ASAP7_75t_L g850 ( 
.A(n_649),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_663),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_684),
.B(n_637),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_637),
.B(n_468),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_731),
.B(n_581),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_637),
.B(n_470),
.Y(n_855)
);

NAND2xp33_ASAP7_75t_L g856 ( 
.A(n_731),
.B(n_616),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_674),
.Y(n_857)
);

NOR2xp67_ASAP7_75t_L g858 ( 
.A(n_667),
.B(n_635),
.Y(n_858)
);

OR2x2_ASAP7_75t_L g859 ( 
.A(n_677),
.B(n_580),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_789),
.Y(n_860)
);

INVx8_ASAP7_75t_L g861 ( 
.A(n_731),
.Y(n_861)
);

AO22x2_ASAP7_75t_L g862 ( 
.A1(n_659),
.A2(n_661),
.B1(n_745),
.B2(n_777),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_684),
.B(n_584),
.Y(n_863)
);

NOR3xp33_ASAP7_75t_L g864 ( 
.A(n_692),
.B(n_406),
.C(n_348),
.Y(n_864)
);

NAND3xp33_ASAP7_75t_L g865 ( 
.A(n_688),
.B(n_626),
.C(n_618),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_731),
.B(n_584),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_676),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_639),
.B(n_472),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_731),
.B(n_586),
.Y(n_869)
);

BUFx6f_ASAP7_75t_SL g870 ( 
.A(n_639),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_697),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_684),
.B(n_586),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_731),
.B(n_753),
.Y(n_873)
);

NOR3xp33_ASAP7_75t_L g874 ( 
.A(n_693),
.B(n_279),
.C(n_276),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_753),
.B(n_587),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_668),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_735),
.B(n_580),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_753),
.B(n_589),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_753),
.B(n_590),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_639),
.B(n_590),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_642),
.A2(n_593),
.B(n_592),
.Y(n_881)
);

NAND3xp33_ASAP7_75t_L g882 ( 
.A(n_650),
.B(n_629),
.C(n_626),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_764),
.B(n_480),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_646),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_779),
.B(n_592),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_749),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_779),
.B(n_785),
.Y(n_887)
);

NAND2xp33_ASAP7_75t_L g888 ( 
.A(n_779),
.B(n_616),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_671),
.B(n_593),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_779),
.B(n_595),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_779),
.A2(n_616),
.B1(n_580),
.B2(n_596),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_736),
.Y(n_892)
);

A2O1A1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_740),
.A2(n_582),
.B(n_569),
.C(n_596),
.Y(n_893)
);

OAI22xp5_ASAP7_75t_SL g894 ( 
.A1(n_768),
.A2(n_497),
.B1(n_498),
.B2(n_481),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_648),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_779),
.B(n_595),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_L g897 ( 
.A1(n_665),
.A2(n_616),
.B1(n_596),
.B2(n_606),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_648),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_716),
.A2(n_606),
.B(n_601),
.Y(n_899)
);

OAI22xp33_ASAP7_75t_L g900 ( 
.A1(n_749),
.A2(n_303),
.B1(n_304),
.B2(n_291),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_741),
.B(n_601),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_741),
.B(n_609),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_741),
.B(n_609),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_736),
.B(n_626),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_658),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_764),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_658),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_741),
.B(n_626),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_703),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_749),
.B(n_626),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_749),
.B(n_651),
.Y(n_911)
);

OAI22x1_ASAP7_75t_R g912 ( 
.A1(n_768),
.A2(n_327),
.B1(n_331),
.B2(n_318),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_662),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_651),
.B(n_626),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_704),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_686),
.B(n_626),
.Y(n_916)
);

AOI22xp33_ASAP7_75t_L g917 ( 
.A1(n_659),
.A2(n_600),
.B1(n_604),
.B2(n_602),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_709),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_722),
.B(n_626),
.Y(n_919)
);

AND2x2_ASAP7_75t_SL g920 ( 
.A(n_767),
.B(n_223),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_747),
.B(n_629),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_662),
.Y(n_922)
);

INVx4_ASAP7_75t_L g923 ( 
.A(n_757),
.Y(n_923)
);

INVx8_ASAP7_75t_L g924 ( 
.A(n_665),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_670),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_660),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_668),
.Y(n_927)
);

INVxp33_ASAP7_75t_L g928 ( 
.A(n_791),
.Y(n_928)
);

INVx5_ASAP7_75t_L g929 ( 
.A(n_669),
.Y(n_929)
);

INVx4_ASAP7_75t_L g930 ( 
.A(n_757),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_657),
.B(n_629),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_670),
.A2(n_604),
.B(n_602),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_661),
.B(n_604),
.Y(n_933)
);

OAI22x1_ASAP7_75t_SL g934 ( 
.A1(n_723),
.A2(n_340),
.B1(n_364),
.B2(n_365),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_SL g935 ( 
.A(n_665),
.B(n_390),
.Y(n_935)
);

NAND2xp33_ASAP7_75t_SL g936 ( 
.A(n_711),
.B(n_629),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_671),
.B(n_629),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_636),
.B(n_629),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_776),
.B(n_337),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_671),
.B(n_629),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_636),
.B(n_629),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_727),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_671),
.B(n_632),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_679),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_SL g945 ( 
.A(n_660),
.B(n_400),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_756),
.Y(n_946)
);

INVxp67_ASAP7_75t_L g947 ( 
.A(n_647),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_668),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_776),
.B(n_344),
.Y(n_949)
);

OAI221xp5_ASAP7_75t_L g950 ( 
.A1(n_761),
.A2(n_378),
.B1(n_382),
.B2(n_291),
.C(n_303),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_671),
.B(n_632),
.Y(n_951)
);

INVx2_ASAP7_75t_SL g952 ( 
.A(n_660),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_776),
.B(n_349),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_673),
.B(n_632),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_L g955 ( 
.A1(n_714),
.A2(n_633),
.B1(n_632),
.B2(n_420),
.Y(n_955)
);

INVx1_ASAP7_75t_SL g956 ( 
.A(n_660),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_729),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_636),
.A2(n_310),
.B1(n_633),
.B2(n_632),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_636),
.B(n_632),
.Y(n_959)
);

NOR2xp67_ASAP7_75t_L g960 ( 
.A(n_715),
.B(n_718),
.Y(n_960)
);

AOI221xp5_ASAP7_75t_L g961 ( 
.A1(n_685),
.A2(n_346),
.B1(n_304),
.B2(n_430),
.C(n_429),
.Y(n_961)
);

NAND2xp33_ASAP7_75t_L g962 ( 
.A(n_666),
.B(n_632),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_794),
.A2(n_755),
.B(n_725),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_826),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_800),
.B(n_672),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_801),
.A2(n_773),
.B(n_763),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_798),
.B(n_672),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_796),
.A2(n_773),
.B(n_763),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_822),
.B(n_672),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_841),
.B(n_672),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_832),
.A2(n_675),
.B(n_679),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_832),
.A2(n_675),
.B(n_683),
.Y(n_972)
);

OAI321xp33_ASAP7_75t_L g973 ( 
.A1(n_900),
.A2(n_382),
.A3(n_430),
.B1(n_429),
.B2(n_422),
.C(n_320),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_825),
.B(n_681),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_835),
.B(n_681),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_926),
.B(n_781),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_827),
.B(n_681),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_952),
.B(n_681),
.Y(n_978)
);

OAI21x1_ASAP7_75t_L g979 ( 
.A1(n_793),
.A2(n_830),
.B(n_932),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_796),
.A2(n_687),
.B(n_683),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_810),
.A2(n_689),
.B(n_687),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_843),
.B(n_647),
.Y(n_982)
);

O2A1O1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_831),
.A2(n_707),
.B(n_702),
.C(n_739),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_893),
.A2(n_744),
.B(n_746),
.C(n_742),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_916),
.A2(n_682),
.B(n_695),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_946),
.A2(n_647),
.B1(n_781),
.B2(n_714),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_810),
.A2(n_682),
.B(n_699),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_877),
.B(n_647),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_858),
.A2(n_682),
.B(n_751),
.C(n_750),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_813),
.A2(n_699),
.B(n_691),
.Y(n_990)
);

O2A1O1Ixp33_ASAP7_75t_SL g991 ( 
.A1(n_852),
.A2(n_752),
.B(n_758),
.C(n_754),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_923),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_844),
.B(n_781),
.Y(n_993)
);

AOI21x1_ASAP7_75t_L g994 ( 
.A1(n_931),
.A2(n_738),
.B(n_769),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_892),
.B(n_696),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_847),
.B(n_696),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_924),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_834),
.B(n_770),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_846),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_816),
.A2(n_700),
.B(n_698),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_851),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_945),
.B(n_673),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_817),
.A2(n_772),
.B1(n_706),
.B2(n_700),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_923),
.Y(n_1004)
);

AO21x1_ASAP7_75t_L g1005 ( 
.A1(n_936),
.A2(n_786),
.B(n_783),
.Y(n_1005)
);

CKINVDCx8_ASAP7_75t_R g1006 ( 
.A(n_828),
.Y(n_1006)
);

AOI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_956),
.A2(n_706),
.B1(n_790),
.B2(n_788),
.Y(n_1007)
);

OAI21xp33_ASAP7_75t_L g1008 ( 
.A1(n_874),
.A2(n_355),
.B(n_351),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_805),
.B(n_698),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_899),
.A2(n_721),
.B(n_713),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_904),
.B(n_713),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_906),
.B(n_886),
.Y(n_1012)
);

OAI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_893),
.A2(n_724),
.B(n_721),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_929),
.B(n_673),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_SL g1015 ( 
.A1(n_852),
.A2(n_706),
.B(n_790),
.C(n_728),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_811),
.B(n_724),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_947),
.B(n_757),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_L g1018 ( 
.A1(n_881),
.A2(n_732),
.B(n_728),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_929),
.A2(n_774),
.B(n_743),
.Y(n_1019)
);

CKINVDCx10_ASAP7_75t_R g1020 ( 
.A(n_870),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_929),
.A2(n_775),
.B(n_774),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_929),
.B(n_673),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_853),
.B(n_775),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_901),
.A2(n_780),
.B1(n_778),
.B2(n_664),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_924),
.Y(n_1025)
);

BUFx12f_ASAP7_75t_L g1026 ( 
.A(n_795),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_894),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_859),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_803),
.A2(n_780),
.B(n_778),
.Y(n_1029)
);

HB1xp67_ASAP7_75t_L g1030 ( 
.A(n_818),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_924),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_821),
.B(n_632),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_923),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_823),
.A2(n_664),
.B(n_666),
.Y(n_1034)
);

BUFx4f_ASAP7_75t_L g1035 ( 
.A(n_924),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_823),
.A2(n_848),
.B(n_829),
.Y(n_1036)
);

NAND3xp33_ASAP7_75t_L g1037 ( 
.A(n_855),
.B(n_788),
.C(n_733),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_960),
.B(n_857),
.Y(n_1038)
);

AOI22xp33_ASAP7_75t_L g1039 ( 
.A1(n_920),
.A2(n_862),
.B1(n_864),
.B2(n_806),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_880),
.A2(n_871),
.B(n_909),
.C(n_867),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_883),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_804),
.A2(n_733),
.B(n_694),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_845),
.Y(n_1043)
);

OAI21xp33_ASAP7_75t_L g1044 ( 
.A1(n_939),
.A2(n_361),
.B(n_358),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_829),
.A2(n_719),
.B(n_666),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_812),
.A2(n_694),
.B(n_673),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_887),
.A2(n_408),
.B(n_401),
.C(n_414),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_848),
.A2(n_719),
.B(n_666),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_863),
.A2(n_719),
.B(n_730),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_915),
.B(n_633),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_863),
.A2(n_719),
.B(n_730),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_868),
.B(n_638),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_928),
.B(n_320),
.Y(n_1053)
);

INVx1_ASAP7_75t_SL g1054 ( 
.A(n_920),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_911),
.B(n_694),
.Y(n_1055)
);

OAI321xp33_ASAP7_75t_L g1056 ( 
.A1(n_950),
.A2(n_352),
.A3(n_422),
.B1(n_378),
.B2(n_350),
.C(n_346),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_815),
.A2(n_748),
.B(n_694),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_902),
.A2(n_414),
.B(n_408),
.C(n_401),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_918),
.B(n_633),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_942),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_845),
.B(n_633),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_949),
.B(n_633),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_903),
.A2(n_336),
.B(n_322),
.C(n_352),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_910),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_957),
.Y(n_1065)
);

OR2x2_ASAP7_75t_L g1066 ( 
.A(n_928),
.B(n_633),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_802),
.Y(n_1067)
);

OR2x6_ASAP7_75t_L g1068 ( 
.A(n_850),
.B(n_678),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_953),
.B(n_807),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_802),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_891),
.A2(n_322),
.B(n_350),
.C(n_338),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_809),
.B(n_633),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_921),
.A2(n_914),
.B(n_919),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_833),
.A2(n_748),
.B(n_694),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_819),
.B(n_678),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_880),
.B(n_367),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_836),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_820),
.B(n_730),
.Y(n_1078)
);

A2O1A1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_840),
.A2(n_338),
.B(n_336),
.C(n_305),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_935),
.B(n_371),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_872),
.A2(n_558),
.B(n_550),
.Y(n_1081)
);

INVx2_ASAP7_75t_SL g1082 ( 
.A(n_912),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_872),
.A2(n_558),
.B(n_550),
.Y(n_1083)
);

O2A1O1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_854),
.A2(n_305),
.B(n_292),
.C(n_299),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_866),
.A2(n_558),
.B(n_550),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_869),
.A2(n_558),
.B(n_550),
.Y(n_1086)
);

AOI21x1_ASAP7_75t_L g1087 ( 
.A1(n_875),
.A2(n_564),
.B(n_561),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_873),
.A2(n_404),
.B1(n_398),
.B2(n_373),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_878),
.A2(n_558),
.B(n_550),
.Y(n_1089)
);

O2A1O1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_879),
.A2(n_402),
.B(n_576),
.C(n_564),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_870),
.B(n_374),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_876),
.B(n_748),
.Y(n_1092)
);

INVx4_ASAP7_75t_L g1093 ( 
.A(n_930),
.Y(n_1093)
);

O2A1O1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_885),
.A2(n_594),
.B(n_576),
.C(n_564),
.Y(n_1094)
);

NAND2xp33_ASAP7_75t_L g1095 ( 
.A(n_850),
.B(n_762),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_890),
.A2(n_896),
.B(n_962),
.Y(n_1096)
);

INVxp67_ASAP7_75t_L g1097 ( 
.A(n_839),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_876),
.B(n_762),
.Y(n_1098)
);

INVxp67_ASAP7_75t_L g1099 ( 
.A(n_961),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_876),
.B(n_762),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_930),
.B(n_836),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_849),
.B(n_762),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_927),
.B(n_762),
.Y(n_1103)
);

AO21x1_ASAP7_75t_L g1104 ( 
.A1(n_936),
.A2(n_576),
.B(n_561),
.Y(n_1104)
);

NAND2x1p5_ASAP7_75t_L g1105 ( 
.A(n_930),
.B(n_561),
.Y(n_1105)
);

INVxp67_ASAP7_75t_L g1106 ( 
.A(n_938),
.Y(n_1106)
);

BUFx2_ASAP7_75t_SL g1107 ( 
.A(n_849),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_802),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_927),
.B(n_948),
.Y(n_1109)
);

AOI21x1_ASAP7_75t_L g1110 ( 
.A1(n_941),
.A2(n_594),
.B(n_669),
.Y(n_1110)
);

INVx3_ASAP7_75t_L g1111 ( 
.A(n_802),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_927),
.B(n_550),
.Y(n_1112)
);

AND2x6_ASAP7_75t_L g1113 ( 
.A(n_897),
.B(n_399),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_962),
.A2(n_558),
.B(n_550),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_882),
.A2(n_558),
.B(n_550),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_948),
.B(n_558),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_959),
.A2(n_594),
.B(n_379),
.C(n_381),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_933),
.A2(n_865),
.B(n_797),
.C(n_842),
.Y(n_1118)
);

BUFx2_ASAP7_75t_L g1119 ( 
.A(n_908),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_850),
.Y(n_1120)
);

NOR2xp67_ASAP7_75t_L g1121 ( 
.A(n_917),
.B(n_220),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_948),
.B(n_570),
.Y(n_1122)
);

NAND3xp33_ASAP7_75t_L g1123 ( 
.A(n_958),
.B(n_389),
.C(n_376),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_797),
.A2(n_583),
.B(n_570),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_884),
.B(n_570),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_895),
.A2(n_397),
.B(n_391),
.Y(n_1126)
);

O2A1O1Ixp33_ASAP7_75t_SL g1127 ( 
.A1(n_814),
.A2(n_8),
.B(n_11),
.C(n_17),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_895),
.A2(n_411),
.B(n_410),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_898),
.B(n_570),
.Y(n_1129)
);

NOR2x1p5_ASAP7_75t_L g1130 ( 
.A(n_934),
.B(n_412),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_842),
.A2(n_570),
.B(n_583),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_850),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_SL g1133 ( 
.A1(n_889),
.A2(n_11),
.B(n_18),
.C(n_21),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_856),
.A2(n_570),
.B(n_583),
.Y(n_1134)
);

BUFx3_ASAP7_75t_L g1135 ( 
.A(n_861),
.Y(n_1135)
);

NAND2xp33_ASAP7_75t_L g1136 ( 
.A(n_861),
.B(n_570),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_861),
.Y(n_1137)
);

O2A1O1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_856),
.A2(n_413),
.B(n_416),
.C(n_423),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_888),
.A2(n_905),
.B(n_898),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_861),
.A2(n_425),
.B1(n_224),
.B2(n_323),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_808),
.A2(n_860),
.B1(n_824),
.B2(n_837),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_888),
.A2(n_583),
.B(n_570),
.Y(n_1142)
);

NOR2x1_ASAP7_75t_L g1143 ( 
.A(n_889),
.B(n_583),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_849),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_905),
.A2(n_583),
.B(n_669),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_907),
.A2(n_583),
.B(n_420),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_967),
.B(n_824),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_963),
.A2(n_799),
.B(n_955),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1099),
.B(n_907),
.Y(n_1149)
);

INVxp67_ASAP7_75t_L g1150 ( 
.A(n_1041),
.Y(n_1150)
);

BUFx12f_ASAP7_75t_L g1151 ( 
.A(n_1026),
.Y(n_1151)
);

O2A1O1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_969),
.A2(n_925),
.B(n_944),
.C(n_913),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_963),
.A2(n_799),
.B(n_913),
.Y(n_1153)
);

NAND2x1p5_ASAP7_75t_L g1154 ( 
.A(n_1132),
.B(n_937),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_966),
.A2(n_925),
.B(n_922),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_998),
.B(n_922),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_R g1157 ( 
.A(n_1020),
.B(n_838),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_974),
.A2(n_944),
.B1(n_837),
.B2(n_860),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_L g1159 ( 
.A(n_970),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1028),
.B(n_937),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_975),
.B(n_940),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_1035),
.Y(n_1162)
);

NAND3xp33_ASAP7_75t_L g1163 ( 
.A(n_965),
.B(n_420),
.C(n_951),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_SL g1164 ( 
.A1(n_1076),
.A2(n_954),
.B(n_951),
.C(n_943),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_1093),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_964),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1027),
.B(n_420),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_1006),
.B(n_940),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1030),
.B(n_943),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1018),
.A2(n_954),
.B(n_583),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_986),
.B(n_225),
.Y(n_1171)
);

OAI22xp33_ASAP7_75t_L g1172 ( 
.A1(n_977),
.A2(n_319),
.B1(n_227),
.B2(n_428),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_1093),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_SL g1174 ( 
.A1(n_983),
.A2(n_18),
.B(n_21),
.C(n_24),
.Y(n_1174)
);

OA22x2_ASAP7_75t_L g1175 ( 
.A1(n_1043),
.A2(n_394),
.B1(n_228),
.B2(n_231),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_997),
.Y(n_1176)
);

O2A1O1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1071),
.A2(n_26),
.B(n_28),
.C(n_29),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_978),
.B(n_1052),
.Y(n_1178)
);

INVx8_ASAP7_75t_L g1179 ( 
.A(n_997),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_997),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_999),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1069),
.A2(n_386),
.B1(n_233),
.B2(n_242),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1001),
.Y(n_1183)
);

A2O1A1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1023),
.A2(n_324),
.B(n_248),
.C(n_427),
.Y(n_1184)
);

NOR3xp33_ASAP7_75t_L g1185 ( 
.A(n_1008),
.B(n_418),
.C(n_252),
.Y(n_1185)
);

AO21x1_ASAP7_75t_L g1186 ( 
.A1(n_966),
.A2(n_335),
.B(n_325),
.Y(n_1186)
);

BUFx4_ASAP7_75t_SL g1187 ( 
.A(n_1037),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_982),
.A2(n_396),
.B1(n_253),
.B2(n_255),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1054),
.B(n_226),
.Y(n_1189)
);

INVx3_ASAP7_75t_L g1190 ( 
.A(n_1135),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1062),
.A2(n_254),
.B(n_325),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1009),
.B(n_26),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_978),
.B(n_261),
.Y(n_1193)
);

O2A1O1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1040),
.A2(n_30),
.B(n_32),
.C(n_35),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1038),
.A2(n_332),
.B(n_267),
.C(n_426),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_SL g1196 ( 
.A1(n_971),
.A2(n_35),
.B(n_37),
.C(n_38),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1060),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1065),
.Y(n_1198)
);

INVx4_ASAP7_75t_L g1199 ( 
.A(n_1025),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1118),
.A2(n_333),
.B(n_268),
.C(n_424),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1136),
.A2(n_325),
.B(n_254),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1053),
.B(n_1080),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1126),
.A2(n_273),
.B(n_278),
.C(n_405),
.Y(n_1203)
);

BUFx8_ASAP7_75t_SL g1204 ( 
.A(n_1025),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_996),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_1025),
.B(n_554),
.Y(n_1206)
);

AOI21x1_ASAP7_75t_L g1207 ( 
.A1(n_994),
.A2(n_1104),
.B(n_1005),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1124),
.A2(n_254),
.B(n_325),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_988),
.B(n_39),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1101),
.B(n_281),
.Y(n_1210)
);

NOR2xp67_ASAP7_75t_SL g1211 ( 
.A(n_1082),
.B(n_287),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1124),
.A2(n_335),
.B(n_325),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_995),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1064),
.B(n_39),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_1012),
.Y(n_1215)
);

O2A1O1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_973),
.A2(n_44),
.B(n_46),
.C(n_49),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_1101),
.B(n_298),
.Y(n_1217)
);

O2A1O1Ixp5_ASAP7_75t_L g1218 ( 
.A1(n_968),
.A2(n_46),
.B(n_51),
.C(n_57),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1016),
.B(n_1119),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1131),
.A2(n_254),
.B(n_335),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1107),
.A2(n_388),
.B1(n_301),
.B2(n_308),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1131),
.A2(n_254),
.B(n_335),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1106),
.B(n_51),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1134),
.A2(n_1142),
.B(n_1073),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1066),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1050),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_1031),
.Y(n_1227)
);

NOR2x1_ASAP7_75t_L g1228 ( 
.A(n_1111),
.B(n_335),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1097),
.B(n_309),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1012),
.B(n_60),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1039),
.B(n_60),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1044),
.B(n_311),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_979),
.A2(n_579),
.B(n_554),
.Y(n_1233)
);

INVx4_ASAP7_75t_L g1234 ( 
.A(n_1031),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1137),
.A2(n_334),
.B1(n_343),
.B2(n_345),
.Y(n_1235)
);

AOI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1091),
.A2(n_385),
.B1(n_369),
.B2(n_357),
.Y(n_1236)
);

O2A1O1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_989),
.A2(n_1063),
.B(n_1079),
.C(n_1128),
.Y(n_1237)
);

AOI32xp33_ASAP7_75t_L g1238 ( 
.A1(n_1056),
.A2(n_61),
.A3(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1077),
.B(n_61),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1134),
.A2(n_579),
.B(n_554),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1059),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_993),
.B(n_64),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1142),
.A2(n_579),
.B(n_554),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_1035),
.B(n_579),
.Y(n_1244)
);

O2A1O1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_1127),
.A2(n_68),
.B(n_69),
.C(n_75),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1031),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1072),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1017),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_1130),
.Y(n_1249)
);

NOR3xp33_ASAP7_75t_SL g1250 ( 
.A(n_1088),
.B(n_77),
.C(n_78),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_984),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1017),
.B(n_579),
.Y(n_1252)
);

INVx6_ASAP7_75t_L g1253 ( 
.A(n_1067),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1138),
.A2(n_579),
.B(n_554),
.C(n_81),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1011),
.B(n_1121),
.Y(n_1255)
);

NOR2xp67_ASAP7_75t_L g1256 ( 
.A(n_1111),
.B(n_579),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1067),
.Y(n_1257)
);

AOI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1087),
.A2(n_579),
.B(n_554),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1073),
.A2(n_554),
.B(n_79),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1125),
.Y(n_1260)
);

AO22x1_ASAP7_75t_L g1261 ( 
.A1(n_1113),
.A2(n_554),
.B1(n_82),
.B2(n_77),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_968),
.A2(n_985),
.B(n_1029),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1109),
.Y(n_1263)
);

BUFx12f_ASAP7_75t_L g1264 ( 
.A(n_1067),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1061),
.B(n_82),
.Y(n_1265)
);

INVx1_ASAP7_75t_SL g1266 ( 
.A(n_1070),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1140),
.B(n_1141),
.Y(n_1267)
);

O2A1O1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1058),
.A2(n_85),
.B(n_93),
.C(n_96),
.Y(n_1268)
);

A2O1A1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1036),
.A2(n_104),
.B(n_110),
.C(n_113),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1129),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_991),
.A2(n_114),
.B(n_117),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_976),
.B(n_127),
.Y(n_1272)
);

BUFx4f_ASAP7_75t_L g1273 ( 
.A(n_1070),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1115),
.A2(n_130),
.B(n_131),
.Y(n_1274)
);

INVx3_ASAP7_75t_L g1275 ( 
.A(n_992),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1115),
.A2(n_133),
.B(n_135),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_992),
.B(n_138),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1113),
.A2(n_143),
.B1(n_144),
.B2(n_147),
.Y(n_1278)
);

AO31x2_ASAP7_75t_L g1279 ( 
.A1(n_1078),
.A2(n_156),
.A3(n_157),
.B(n_158),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_1004),
.B(n_160),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1049),
.A2(n_168),
.B(n_169),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1075),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1070),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1108),
.Y(n_1284)
);

AOI22x1_ASAP7_75t_L g1285 ( 
.A1(n_987),
.A2(n_180),
.B1(n_181),
.B2(n_185),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1032),
.B(n_192),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1113),
.B(n_194),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1144),
.A2(n_195),
.B1(n_197),
.B2(n_199),
.Y(n_1288)
);

INVx4_ASAP7_75t_L g1289 ( 
.A(n_1068),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1113),
.B(n_200),
.Y(n_1290)
);

NAND3xp33_ASAP7_75t_SL g1291 ( 
.A(n_1084),
.B(n_202),
.C(n_203),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1123),
.B(n_206),
.Y(n_1292)
);

A2O1A1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1096),
.A2(n_207),
.B(n_208),
.C(n_214),
.Y(n_1293)
);

NAND2xp33_ASAP7_75t_SL g1294 ( 
.A(n_1144),
.B(n_1120),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_1108),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1033),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1068),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1112),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1113),
.B(n_1002),
.Y(n_1299)
);

NOR3xp33_ASAP7_75t_SL g1300 ( 
.A(n_1047),
.B(n_972),
.C(n_1122),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1116),
.Y(n_1301)
);

BUFx3_ASAP7_75t_L g1302 ( 
.A(n_1068),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1051),
.A2(n_980),
.B(n_981),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1143),
.Y(n_1304)
);

NAND2x1p5_ASAP7_75t_L g1305 ( 
.A(n_1120),
.B(n_1055),
.Y(n_1305)
);

INVx3_ASAP7_75t_L g1306 ( 
.A(n_1105),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1007),
.B(n_1013),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1105),
.Y(n_1308)
);

AOI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1231),
.A2(n_1003),
.B1(n_1024),
.B2(n_1133),
.Y(n_1309)
);

O2A1O1Ixp33_ASAP7_75t_L g1310 ( 
.A1(n_1192),
.A2(n_1117),
.B(n_1015),
.C(n_1010),
.Y(n_1310)
);

BUFx3_ASAP7_75t_L g1311 ( 
.A(n_1204),
.Y(n_1311)
);

OAI21xp33_ASAP7_75t_L g1312 ( 
.A1(n_1250),
.A2(n_980),
.B(n_981),
.Y(n_1312)
);

AO31x2_ASAP7_75t_L g1313 ( 
.A1(n_1186),
.A2(n_1146),
.A3(n_1139),
.B(n_1089),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1170),
.A2(n_1146),
.B(n_1110),
.Y(n_1314)
);

BUFx6f_ASAP7_75t_L g1315 ( 
.A(n_1264),
.Y(n_1315)
);

AOI221x1_ASAP7_75t_L g1316 ( 
.A1(n_1259),
.A2(n_1114),
.B1(n_1085),
.B2(n_1086),
.C(n_1089),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1153),
.A2(n_1155),
.B(n_1224),
.Y(n_1317)
);

AOI211x1_ASAP7_75t_L g1318 ( 
.A1(n_1209),
.A2(n_990),
.B(n_1081),
.C(n_1083),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1300),
.A2(n_1086),
.B(n_1085),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1151),
.Y(n_1320)
);

AO32x2_ASAP7_75t_L g1321 ( 
.A1(n_1158),
.A2(n_1090),
.A3(n_1094),
.B1(n_1139),
.B2(n_1114),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1155),
.A2(n_1145),
.B(n_1000),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1224),
.A2(n_1145),
.B(n_1095),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1286),
.A2(n_1021),
.B(n_1019),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1166),
.Y(n_1325)
);

INVx2_ASAP7_75t_SL g1326 ( 
.A(n_1295),
.Y(n_1326)
);

O2A1O1Ixp33_ASAP7_75t_SL g1327 ( 
.A1(n_1164),
.A2(n_1200),
.B(n_1203),
.C(n_1196),
.Y(n_1327)
);

INVx2_ASAP7_75t_SL g1328 ( 
.A(n_1179),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1303),
.A2(n_1081),
.B(n_1045),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1181),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1262),
.A2(n_1048),
.B(n_1034),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1150),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1183),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1159),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1197),
.Y(n_1335)
);

OAI22x1_ASAP7_75t_L g1336 ( 
.A1(n_1171),
.A2(n_1103),
.B1(n_1100),
.B2(n_1098),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1149),
.B(n_1092),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1307),
.A2(n_1042),
.B1(n_1046),
.B2(n_1057),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1198),
.Y(n_1339)
);

NAND3xp33_ASAP7_75t_SL g1340 ( 
.A(n_1194),
.B(n_1074),
.C(n_1022),
.Y(n_1340)
);

NOR2x1_ASAP7_75t_L g1341 ( 
.A(n_1283),
.B(n_1014),
.Y(n_1341)
);

OA21x2_ASAP7_75t_L g1342 ( 
.A1(n_1262),
.A2(n_1102),
.B(n_1303),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1168),
.B(n_1229),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1167),
.B(n_1215),
.Y(n_1344)
);

BUFx12f_ASAP7_75t_L g1345 ( 
.A(n_1249),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1156),
.B(n_1205),
.Y(n_1346)
);

NOR3xp33_ASAP7_75t_SL g1347 ( 
.A(n_1242),
.B(n_1239),
.C(n_1217),
.Y(n_1347)
);

A2O1A1Ixp33_ASAP7_75t_L g1348 ( 
.A1(n_1216),
.A2(n_1237),
.B(n_1194),
.C(n_1232),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1294),
.A2(n_1201),
.B(n_1148),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1161),
.B(n_1251),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1271),
.A2(n_1241),
.B(n_1226),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1233),
.A2(n_1258),
.B(n_1207),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1271),
.A2(n_1191),
.B(n_1281),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1147),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1189),
.B(n_1236),
.Y(n_1355)
);

BUFx6f_ASAP7_75t_L g1356 ( 
.A(n_1273),
.Y(n_1356)
);

INVx8_ASAP7_75t_L g1357 ( 
.A(n_1179),
.Y(n_1357)
);

OA21x2_ASAP7_75t_L g1358 ( 
.A1(n_1191),
.A2(n_1220),
.B(n_1208),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_1273),
.Y(n_1359)
);

NOR4xp25_ASAP7_75t_L g1360 ( 
.A(n_1216),
.B(n_1177),
.C(n_1245),
.D(n_1237),
.Y(n_1360)
);

O2A1O1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1174),
.A2(n_1177),
.B(n_1184),
.C(n_1245),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1193),
.B(n_1230),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1225),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1208),
.A2(n_1220),
.B(n_1222),
.Y(n_1364)
);

OA21x2_ASAP7_75t_L g1365 ( 
.A1(n_1212),
.A2(n_1222),
.B(n_1276),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1274),
.A2(n_1298),
.B(n_1301),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_L g1367 ( 
.A(n_1297),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1213),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1282),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1212),
.A2(n_1277),
.B(n_1280),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1214),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1223),
.A2(n_1265),
.B1(n_1267),
.B2(n_1178),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1152),
.A2(n_1293),
.B(n_1263),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1152),
.A2(n_1243),
.B(n_1240),
.Y(n_1374)
);

INVx3_ASAP7_75t_SL g1375 ( 
.A(n_1179),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1187),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1219),
.A2(n_1278),
.B1(n_1254),
.B2(n_1160),
.Y(n_1377)
);

AO21x1_ASAP7_75t_L g1378 ( 
.A1(n_1292),
.A2(n_1268),
.B(n_1255),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1299),
.A2(n_1247),
.B(n_1269),
.Y(n_1379)
);

AOI221x1_ASAP7_75t_L g1380 ( 
.A1(n_1291),
.A2(n_1163),
.B1(n_1288),
.B2(n_1185),
.C(n_1290),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1157),
.B(n_1248),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1291),
.A2(n_1260),
.B(n_1270),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1169),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1275),
.B(n_1296),
.Y(n_1384)
);

A2O1A1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1268),
.A2(n_1272),
.B(n_1218),
.C(n_1195),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1284),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1287),
.A2(n_1275),
.B(n_1296),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1165),
.A2(n_1173),
.B(n_1261),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1266),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1253),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1175),
.B(n_1246),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1218),
.A2(n_1240),
.B(n_1243),
.Y(n_1392)
);

NOR2xp67_ASAP7_75t_SL g1393 ( 
.A(n_1165),
.B(n_1173),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_1302),
.B(n_1162),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1175),
.B(n_1227),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1285),
.A2(n_1228),
.B(n_1305),
.Y(n_1396)
);

A2O1A1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1182),
.A2(n_1188),
.B(n_1210),
.C(n_1190),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1289),
.B(n_1297),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1305),
.A2(n_1306),
.B(n_1154),
.Y(n_1399)
);

AO31x2_ASAP7_75t_L g1400 ( 
.A1(n_1279),
.A2(n_1289),
.A3(n_1235),
.B(n_1221),
.Y(n_1400)
);

BUFx2_ASAP7_75t_L g1401 ( 
.A(n_1257),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1190),
.B(n_1252),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1253),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1306),
.A2(n_1154),
.B(n_1244),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_SL g1405 ( 
.A(n_1211),
.B(n_1297),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1176),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_SL g1407 ( 
.A(n_1257),
.B(n_1176),
.Y(n_1407)
);

BUFx8_ASAP7_75t_L g1408 ( 
.A(n_1176),
.Y(n_1408)
);

A2O1A1Ixp33_ASAP7_75t_L g1409 ( 
.A1(n_1256),
.A2(n_1252),
.B(n_1308),
.C(n_1206),
.Y(n_1409)
);

CKINVDCx20_ASAP7_75t_R g1410 ( 
.A(n_1180),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1257),
.B(n_1308),
.Y(n_1411)
);

NOR2xp67_ASAP7_75t_SL g1412 ( 
.A(n_1180),
.B(n_1199),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_SL g1413 ( 
.A(n_1180),
.B(n_1308),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1279),
.A2(n_1253),
.B(n_1199),
.Y(n_1414)
);

NAND2x1p5_ASAP7_75t_L g1415 ( 
.A(n_1234),
.B(n_1206),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1234),
.B(n_1172),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1279),
.A2(n_1136),
.B(n_1224),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1156),
.B(n_1205),
.Y(n_1418)
);

A2O1A1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1238),
.A2(n_998),
.B(n_975),
.C(n_1023),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1202),
.B(n_798),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1202),
.B(n_798),
.Y(n_1421)
);

AOI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1231),
.A2(n_975),
.B1(n_834),
.B2(n_855),
.Y(n_1422)
);

NAND3xp33_ASAP7_75t_L g1423 ( 
.A(n_1238),
.B(n_1194),
.C(n_998),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1170),
.A2(n_1153),
.B(n_1155),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1300),
.A2(n_1259),
.B(n_1153),
.Y(n_1425)
);

AOI221x1_ASAP7_75t_L g1426 ( 
.A1(n_1231),
.A2(n_862),
.B1(n_1259),
.B2(n_1148),
.C(n_1281),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1170),
.A2(n_1153),
.B(n_1155),
.Y(n_1427)
);

O2A1O1Ixp33_ASAP7_75t_SL g1428 ( 
.A1(n_1164),
.A2(n_852),
.B(n_880),
.C(n_1200),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_SL g1429 ( 
.A(n_1161),
.B(n_975),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_L g1430 ( 
.A(n_1264),
.Y(n_1430)
);

AOI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1231),
.A2(n_975),
.B1(n_834),
.B2(n_855),
.Y(n_1431)
);

OAI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1300),
.A2(n_1259),
.B(n_1153),
.Y(n_1432)
);

INVx8_ASAP7_75t_L g1433 ( 
.A(n_1179),
.Y(n_1433)
);

AO32x2_ASAP7_75t_L g1434 ( 
.A1(n_1158),
.A2(n_627),
.A3(n_1024),
.B1(n_1289),
.B2(n_1003),
.Y(n_1434)
);

BUFx6f_ASAP7_75t_L g1435 ( 
.A(n_1264),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1202),
.B(n_798),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1289),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1224),
.A2(n_1136),
.B(n_1286),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1202),
.B(n_798),
.Y(n_1439)
);

OR2x6_ASAP7_75t_L g1440 ( 
.A(n_1151),
.B(n_924),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1202),
.B(n_798),
.Y(n_1441)
);

OAI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1300),
.A2(n_1259),
.B(n_1153),
.Y(n_1442)
);

AO32x2_ASAP7_75t_L g1443 ( 
.A1(n_1158),
.A2(n_627),
.A3(n_1024),
.B1(n_1289),
.B2(n_1003),
.Y(n_1443)
);

OAI21xp5_ASAP7_75t_SL g1444 ( 
.A1(n_1238),
.A2(n_800),
.B(n_975),
.Y(n_1444)
);

BUFx10_ASAP7_75t_L g1445 ( 
.A(n_1193),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1224),
.A2(n_1136),
.B(n_1286),
.Y(n_1446)
);

NOR2x1_ASAP7_75t_SL g1447 ( 
.A(n_1289),
.B(n_1107),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1224),
.A2(n_1136),
.B(n_1286),
.Y(n_1448)
);

BUFx12f_ASAP7_75t_L g1449 ( 
.A(n_1151),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1224),
.A2(n_1136),
.B(n_1286),
.Y(n_1450)
);

O2A1O1Ixp33_ASAP7_75t_SL g1451 ( 
.A1(n_1164),
.A2(n_852),
.B(n_880),
.C(n_1200),
.Y(n_1451)
);

INVx3_ASAP7_75t_L g1452 ( 
.A(n_1289),
.Y(n_1452)
);

AND2x6_ASAP7_75t_L g1453 ( 
.A(n_1297),
.B(n_1302),
.Y(n_1453)
);

NOR2xp67_ASAP7_75t_L g1454 ( 
.A(n_1150),
.B(n_800),
.Y(n_1454)
);

OAI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1300),
.A2(n_1259),
.B(n_1153),
.Y(n_1455)
);

O2A1O1Ixp5_ASAP7_75t_SL g1456 ( 
.A1(n_1171),
.A2(n_475),
.B(n_483),
.C(n_482),
.Y(n_1456)
);

A2O1A1Ixp33_ASAP7_75t_L g1457 ( 
.A1(n_1238),
.A2(n_998),
.B(n_975),
.C(n_1023),
.Y(n_1457)
);

NOR4xp25_ASAP7_75t_L g1458 ( 
.A(n_1216),
.B(n_1194),
.C(n_1177),
.D(n_1238),
.Y(n_1458)
);

BUFx10_ASAP7_75t_L g1459 ( 
.A(n_1193),
.Y(n_1459)
);

INVx3_ASAP7_75t_L g1460 ( 
.A(n_1289),
.Y(n_1460)
);

BUFx4_ASAP7_75t_R g1461 ( 
.A(n_1204),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1156),
.B(n_1205),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1170),
.A2(n_1153),
.B(n_1155),
.Y(n_1463)
);

AOI31xp67_ASAP7_75t_L g1464 ( 
.A1(n_1304),
.A2(n_1247),
.A3(n_1301),
.B(n_1298),
.Y(n_1464)
);

AO21x1_ASAP7_75t_L g1465 ( 
.A1(n_1194),
.A2(n_1192),
.B(n_1216),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1156),
.B(n_1205),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1325),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1330),
.Y(n_1468)
);

INVx6_ASAP7_75t_L g1469 ( 
.A(n_1408),
.Y(n_1469)
);

OAI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1423),
.A2(n_1444),
.B1(n_1431),
.B2(n_1422),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1355),
.A2(n_1422),
.B1(n_1431),
.B2(n_1423),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1419),
.A2(n_1457),
.B1(n_1444),
.B2(n_1343),
.Y(n_1472)
);

AOI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1362),
.A2(n_1454),
.B1(n_1405),
.B2(n_1429),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1333),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1335),
.Y(n_1475)
);

INVx6_ASAP7_75t_L g1476 ( 
.A(n_1408),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_SL g1477 ( 
.A1(n_1376),
.A2(n_1458),
.B1(n_1360),
.B2(n_1326),
.Y(n_1477)
);

CKINVDCx11_ASAP7_75t_R g1478 ( 
.A(n_1449),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1465),
.A2(n_1420),
.B1(n_1441),
.B2(n_1372),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1421),
.A2(n_1436),
.B1(n_1439),
.B2(n_1371),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1339),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1378),
.A2(n_1354),
.B1(n_1369),
.B2(n_1466),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1410),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1363),
.Y(n_1484)
);

AOI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1348),
.A2(n_1347),
.B1(n_1458),
.B2(n_1381),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1385),
.A2(n_1397),
.B1(n_1332),
.B2(n_1350),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_SL g1487 ( 
.A1(n_1377),
.A2(n_1391),
.B1(n_1466),
.B2(n_1462),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1346),
.A2(n_1462),
.B1(n_1418),
.B2(n_1344),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1368),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1383),
.Y(n_1490)
);

AOI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1395),
.A2(n_1445),
.B1(n_1459),
.B2(n_1377),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1311),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1346),
.A2(n_1418),
.B1(n_1350),
.B2(n_1445),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1334),
.B(n_1459),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_L g1495 ( 
.A(n_1357),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1340),
.A2(n_1337),
.B1(n_1338),
.B2(n_1425),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1464),
.Y(n_1497)
);

INVx4_ASAP7_75t_L g1498 ( 
.A(n_1461),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1389),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1338),
.A2(n_1425),
.B1(n_1455),
.B2(n_1432),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1345),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_1315),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1386),
.Y(n_1503)
);

INVx6_ASAP7_75t_L g1504 ( 
.A(n_1357),
.Y(n_1504)
);

CKINVDCx14_ASAP7_75t_R g1505 ( 
.A(n_1315),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1402),
.B(n_1453),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1384),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1394),
.B(n_1440),
.Y(n_1508)
);

OAI21xp5_ASAP7_75t_SL g1509 ( 
.A1(n_1361),
.A2(n_1442),
.B(n_1432),
.Y(n_1509)
);

CKINVDCx6p67_ASAP7_75t_R g1510 ( 
.A(n_1375),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_1320),
.Y(n_1511)
);

BUFx2_ASAP7_75t_L g1512 ( 
.A(n_1401),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1411),
.Y(n_1513)
);

CKINVDCx11_ASAP7_75t_R g1514 ( 
.A(n_1315),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1411),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1398),
.Y(n_1516)
);

CKINVDCx20_ASAP7_75t_R g1517 ( 
.A(n_1430),
.Y(n_1517)
);

BUFx4f_ASAP7_75t_L g1518 ( 
.A(n_1356),
.Y(n_1518)
);

CKINVDCx11_ASAP7_75t_R g1519 ( 
.A(n_1430),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1309),
.A2(n_1442),
.B1(n_1455),
.B2(n_1416),
.Y(n_1520)
);

OAI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1426),
.A2(n_1309),
.B1(n_1416),
.B2(n_1380),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1390),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1398),
.Y(n_1523)
);

NAND2x1p5_ASAP7_75t_L g1524 ( 
.A(n_1367),
.B(n_1412),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1403),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1360),
.A2(n_1382),
.B1(n_1453),
.B2(n_1319),
.Y(n_1526)
);

NAND2x1p5_ASAP7_75t_L g1527 ( 
.A(n_1367),
.B(n_1356),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1367),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_SL g1529 ( 
.A1(n_1319),
.A2(n_1453),
.B1(n_1373),
.B2(n_1434),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1435),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_1435),
.Y(n_1531)
);

OAI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1440),
.A2(n_1415),
.B1(n_1460),
.B2(n_1452),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1399),
.Y(n_1533)
);

CKINVDCx6p67_ASAP7_75t_R g1534 ( 
.A(n_1440),
.Y(n_1534)
);

OAI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1415),
.A2(n_1437),
.B1(n_1460),
.B2(n_1452),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1414),
.Y(n_1536)
);

BUFx12f_ASAP7_75t_SL g1537 ( 
.A(n_1356),
.Y(n_1537)
);

BUFx2_ASAP7_75t_SL g1538 ( 
.A(n_1359),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1453),
.A2(n_1312),
.B1(n_1394),
.B2(n_1336),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1312),
.A2(n_1366),
.B1(n_1379),
.B2(n_1351),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1413),
.Y(n_1541)
);

AOI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1359),
.A2(n_1437),
.B1(n_1409),
.B2(n_1393),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1359),
.A2(n_1392),
.B1(n_1349),
.B2(n_1353),
.Y(n_1543)
);

INVx8_ASAP7_75t_L g1544 ( 
.A(n_1433),
.Y(n_1544)
);

INVx6_ASAP7_75t_L g1545 ( 
.A(n_1433),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1392),
.A2(n_1341),
.B1(n_1365),
.B2(n_1417),
.Y(n_1546)
);

OAI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1388),
.A2(n_1406),
.B1(n_1328),
.B2(n_1316),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1433),
.Y(n_1548)
);

INVx6_ASAP7_75t_L g1549 ( 
.A(n_1447),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1407),
.Y(n_1550)
);

CKINVDCx11_ASAP7_75t_R g1551 ( 
.A(n_1318),
.Y(n_1551)
);

INVx1_ASAP7_75t_SL g1552 ( 
.A(n_1387),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1365),
.A2(n_1370),
.B1(n_1358),
.B2(n_1443),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1400),
.B(n_1404),
.Y(n_1554)
);

INVx3_ASAP7_75t_L g1555 ( 
.A(n_1400),
.Y(n_1555)
);

INVxp67_ASAP7_75t_L g1556 ( 
.A(n_1342),
.Y(n_1556)
);

BUFx12f_ASAP7_75t_L g1557 ( 
.A(n_1327),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1358),
.A2(n_1434),
.B1(n_1443),
.B2(n_1364),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1434),
.A2(n_1443),
.B1(n_1450),
.B2(n_1448),
.Y(n_1559)
);

BUFx10_ASAP7_75t_L g1560 ( 
.A(n_1428),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_SL g1561 ( 
.A1(n_1438),
.A2(n_1446),
.B1(n_1374),
.B2(n_1396),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1313),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1313),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1324),
.A2(n_1323),
.B1(n_1317),
.B2(n_1331),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1310),
.A2(n_1451),
.B1(n_1456),
.B2(n_1321),
.Y(n_1565)
);

BUFx12f_ASAP7_75t_L g1566 ( 
.A(n_1321),
.Y(n_1566)
);

AOI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1314),
.A2(n_1352),
.B1(n_1329),
.B2(n_1322),
.Y(n_1567)
);

BUFx10_ASAP7_75t_L g1568 ( 
.A(n_1321),
.Y(n_1568)
);

BUFx8_ASAP7_75t_L g1569 ( 
.A(n_1424),
.Y(n_1569)
);

INVx3_ASAP7_75t_SL g1570 ( 
.A(n_1427),
.Y(n_1570)
);

BUFx6f_ASAP7_75t_L g1571 ( 
.A(n_1463),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1325),
.Y(n_1572)
);

CKINVDCx11_ASAP7_75t_R g1573 ( 
.A(n_1449),
.Y(n_1573)
);

INVx2_ASAP7_75t_SL g1574 ( 
.A(n_1311),
.Y(n_1574)
);

INVx4_ASAP7_75t_L g1575 ( 
.A(n_1461),
.Y(n_1575)
);

INVx6_ASAP7_75t_L g1576 ( 
.A(n_1408),
.Y(n_1576)
);

AOI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1355),
.A2(n_834),
.B1(n_975),
.B2(n_855),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_1461),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1423),
.A2(n_806),
.B1(n_1039),
.B2(n_659),
.Y(n_1579)
);

BUFx6f_ASAP7_75t_L g1580 ( 
.A(n_1357),
.Y(n_1580)
);

BUFx3_ASAP7_75t_L g1581 ( 
.A(n_1311),
.Y(n_1581)
);

BUFx2_ASAP7_75t_SL g1582 ( 
.A(n_1410),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1423),
.A2(n_806),
.B1(n_1039),
.B2(n_659),
.Y(n_1583)
);

INVx4_ASAP7_75t_L g1584 ( 
.A(n_1461),
.Y(n_1584)
);

CKINVDCx20_ASAP7_75t_R g1585 ( 
.A(n_1311),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1423),
.A2(n_806),
.B1(n_1039),
.B2(n_659),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1355),
.A2(n_1422),
.B1(n_1431),
.B2(n_1423),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_SL g1588 ( 
.A(n_1408),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_SL g1589 ( 
.A1(n_1423),
.A2(n_607),
.B1(n_659),
.B2(n_834),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1423),
.A2(n_806),
.B1(n_1039),
.B2(n_659),
.Y(n_1590)
);

CKINVDCx20_ASAP7_75t_R g1591 ( 
.A(n_1311),
.Y(n_1591)
);

CKINVDCx11_ASAP7_75t_R g1592 ( 
.A(n_1449),
.Y(n_1592)
);

CKINVDCx11_ASAP7_75t_R g1593 ( 
.A(n_1449),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1325),
.Y(n_1594)
);

CKINVDCx6p67_ASAP7_75t_R g1595 ( 
.A(n_1449),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1354),
.B(n_1367),
.Y(n_1596)
);

INVx6_ASAP7_75t_L g1597 ( 
.A(n_1408),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1423),
.A2(n_806),
.B1(n_1039),
.B2(n_659),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_SL g1599 ( 
.A1(n_1423),
.A2(n_607),
.B1(n_659),
.B2(n_834),
.Y(n_1599)
);

OAI22x1_ASAP7_75t_L g1600 ( 
.A1(n_1422),
.A2(n_1431),
.B1(n_1355),
.B2(n_1423),
.Y(n_1600)
);

BUFx6f_ASAP7_75t_SL g1601 ( 
.A(n_1311),
.Y(n_1601)
);

BUFx4f_ASAP7_75t_SL g1602 ( 
.A(n_1449),
.Y(n_1602)
);

OAI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1423),
.A2(n_1444),
.B1(n_1422),
.B2(n_1431),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1325),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1423),
.A2(n_806),
.B1(n_1039),
.B2(n_659),
.Y(n_1605)
);

BUFx8_ASAP7_75t_L g1606 ( 
.A(n_1449),
.Y(n_1606)
);

OAI21xp5_ASAP7_75t_SL g1607 ( 
.A1(n_1355),
.A2(n_1444),
.B(n_1423),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_SL g1608 ( 
.A1(n_1423),
.A2(n_607),
.B1(n_659),
.B2(n_834),
.Y(n_1608)
);

CKINVDCx20_ASAP7_75t_R g1609 ( 
.A(n_1311),
.Y(n_1609)
);

BUFx6f_ASAP7_75t_L g1610 ( 
.A(n_1357),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1325),
.Y(n_1611)
);

BUFx3_ASAP7_75t_L g1612 ( 
.A(n_1311),
.Y(n_1612)
);

OAI22xp33_ASAP7_75t_R g1613 ( 
.A1(n_1355),
.A2(n_494),
.B1(n_229),
.B2(n_246),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1346),
.B(n_1418),
.Y(n_1614)
);

BUFx3_ASAP7_75t_L g1615 ( 
.A(n_1311),
.Y(n_1615)
);

CKINVDCx11_ASAP7_75t_R g1616 ( 
.A(n_1449),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1423),
.A2(n_806),
.B1(n_1039),
.B2(n_659),
.Y(n_1617)
);

BUFx10_ASAP7_75t_L g1618 ( 
.A(n_1315),
.Y(n_1618)
);

INVx8_ASAP7_75t_L g1619 ( 
.A(n_1357),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1325),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1355),
.A2(n_1422),
.B1(n_1431),
.B2(n_1423),
.Y(n_1621)
);

AOI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1613),
.A2(n_1621),
.B1(n_1587),
.B2(n_1471),
.Y(n_1622)
);

BUFx4f_ASAP7_75t_L g1623 ( 
.A(n_1469),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1497),
.Y(n_1624)
);

INVx3_ASAP7_75t_L g1625 ( 
.A(n_1569),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_1478),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1507),
.Y(n_1627)
);

INVx3_ASAP7_75t_L g1628 ( 
.A(n_1569),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1566),
.Y(n_1629)
);

A2O1A1Ixp33_ASAP7_75t_L g1630 ( 
.A1(n_1577),
.A2(n_1607),
.B(n_1589),
.C(n_1599),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1562),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1563),
.Y(n_1632)
);

BUFx8_ASAP7_75t_L g1633 ( 
.A(n_1601),
.Y(n_1633)
);

AOI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1600),
.A2(n_1470),
.B1(n_1603),
.B2(n_1472),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1533),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1554),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1620),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1467),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1468),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1474),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1525),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1475),
.Y(n_1642)
);

OAI21x1_ASAP7_75t_L g1643 ( 
.A1(n_1564),
.A2(n_1540),
.B(n_1546),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1481),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1572),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1594),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1470),
.A2(n_1603),
.B1(n_1485),
.B2(n_1500),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1500),
.B(n_1568),
.Y(n_1648)
);

BUFx4f_ASAP7_75t_SL g1649 ( 
.A(n_1585),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1604),
.Y(n_1650)
);

INVx3_ASAP7_75t_L g1651 ( 
.A(n_1571),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1611),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1490),
.Y(n_1653)
);

CKINVDCx6p67_ASAP7_75t_R g1654 ( 
.A(n_1573),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1520),
.Y(n_1655)
);

A2O1A1Ixp33_ASAP7_75t_L g1656 ( 
.A1(n_1589),
.A2(n_1599),
.B(n_1608),
.C(n_1479),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1516),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_SL g1658 ( 
.A(n_1532),
.B(n_1535),
.Y(n_1658)
);

INVxp67_ASAP7_75t_L g1659 ( 
.A(n_1494),
.Y(n_1659)
);

AO21x2_ASAP7_75t_L g1660 ( 
.A1(n_1521),
.A2(n_1565),
.B(n_1567),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1568),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1555),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1555),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1571),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1489),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1496),
.B(n_1529),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1513),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1536),
.B(n_1556),
.Y(n_1668)
);

AO21x2_ASAP7_75t_L g1669 ( 
.A1(n_1521),
.A2(n_1509),
.B(n_1547),
.Y(n_1669)
);

INVxp67_ASAP7_75t_SL g1670 ( 
.A(n_1556),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1515),
.Y(n_1671)
);

NOR2x1_ASAP7_75t_SL g1672 ( 
.A(n_1486),
.B(n_1557),
.Y(n_1672)
);

OAI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1496),
.A2(n_1608),
.B(n_1526),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1552),
.Y(n_1674)
);

BUFx12f_ASAP7_75t_L g1675 ( 
.A(n_1592),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1523),
.Y(n_1676)
);

HB1xp67_ASAP7_75t_L g1677 ( 
.A(n_1512),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1529),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1484),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1558),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1558),
.Y(n_1681)
);

OAI21x1_ASAP7_75t_L g1682 ( 
.A1(n_1540),
.A2(n_1546),
.B(n_1543),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1551),
.Y(n_1683)
);

OAI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1479),
.A2(n_1477),
.B1(n_1487),
.B2(n_1526),
.Y(n_1684)
);

BUFx2_ASAP7_75t_L g1685 ( 
.A(n_1570),
.Y(n_1685)
);

BUFx3_ASAP7_75t_L g1686 ( 
.A(n_1469),
.Y(n_1686)
);

HB1xp67_ASAP7_75t_L g1687 ( 
.A(n_1550),
.Y(n_1687)
);

OAI21x1_ASAP7_75t_L g1688 ( 
.A1(n_1543),
.A2(n_1553),
.B(n_1559),
.Y(n_1688)
);

BUFx6f_ASAP7_75t_L g1689 ( 
.A(n_1549),
.Y(n_1689)
);

OR2x6_ASAP7_75t_L g1690 ( 
.A(n_1506),
.B(n_1476),
.Y(n_1690)
);

AO21x2_ASAP7_75t_L g1691 ( 
.A1(n_1547),
.A2(n_1614),
.B(n_1499),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1559),
.B(n_1553),
.Y(n_1692)
);

CKINVDCx20_ASAP7_75t_R g1693 ( 
.A(n_1593),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1482),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1482),
.Y(n_1695)
);

INVxp67_ASAP7_75t_SL g1696 ( 
.A(n_1493),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1522),
.Y(n_1697)
);

OAI21x1_ASAP7_75t_L g1698 ( 
.A1(n_1539),
.A2(n_1493),
.B(n_1541),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1503),
.Y(n_1699)
);

BUFx3_ASAP7_75t_L g1700 ( 
.A(n_1476),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1570),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1487),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1561),
.Y(n_1703)
);

OAI21x1_ASAP7_75t_L g1704 ( 
.A1(n_1539),
.A2(n_1528),
.B(n_1491),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1596),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1561),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1488),
.Y(n_1707)
);

CKINVDCx6p67_ASAP7_75t_R g1708 ( 
.A(n_1616),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1488),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1560),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1560),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1532),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1480),
.B(n_1473),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1542),
.Y(n_1714)
);

OR2x6_ASAP7_75t_L g1715 ( 
.A(n_1476),
.B(n_1597),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1480),
.Y(n_1716)
);

AOI21x1_ASAP7_75t_L g1717 ( 
.A1(n_1508),
.A2(n_1483),
.B(n_1534),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1524),
.Y(n_1718)
);

OAI21x1_ASAP7_75t_L g1719 ( 
.A1(n_1527),
.A2(n_1579),
.B(n_1617),
.Y(n_1719)
);

AO21x2_ASAP7_75t_L g1720 ( 
.A1(n_1579),
.A2(n_1586),
.B(n_1583),
.Y(n_1720)
);

INVx4_ASAP7_75t_L g1721 ( 
.A(n_1495),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1537),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1538),
.Y(n_1723)
);

INVx4_ASAP7_75t_L g1724 ( 
.A(n_1495),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1495),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1576),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1582),
.B(n_1590),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1498),
.B(n_1575),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1498),
.B(n_1575),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1584),
.B(n_1597),
.Y(n_1730)
);

OAI21x1_ASAP7_75t_L g1731 ( 
.A1(n_1583),
.A2(n_1586),
.B(n_1617),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1580),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1502),
.Y(n_1733)
);

OA21x2_ASAP7_75t_L g1734 ( 
.A1(n_1590),
.A2(n_1605),
.B(n_1598),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1580),
.Y(n_1735)
);

HB1xp67_ASAP7_75t_L g1736 ( 
.A(n_1530),
.Y(n_1736)
);

OAI21x1_ASAP7_75t_L g1737 ( 
.A1(n_1598),
.A2(n_1605),
.B(n_1588),
.Y(n_1737)
);

INVx2_ASAP7_75t_SL g1738 ( 
.A(n_1618),
.Y(n_1738)
);

OA21x2_ASAP7_75t_L g1739 ( 
.A1(n_1531),
.A2(n_1548),
.B(n_1511),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1610),
.Y(n_1740)
);

OAI21x1_ASAP7_75t_L g1741 ( 
.A1(n_1588),
.A2(n_1545),
.B(n_1504),
.Y(n_1741)
);

AND2x6_ASAP7_75t_SL g1742 ( 
.A(n_1602),
.B(n_1606),
.Y(n_1742)
);

BUFx12f_ASAP7_75t_L g1743 ( 
.A(n_1606),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1657),
.B(n_1584),
.Y(n_1744)
);

A2O1A1Ixp33_ASAP7_75t_L g1745 ( 
.A1(n_1630),
.A2(n_1518),
.B(n_1505),
.C(n_1574),
.Y(n_1745)
);

AND2x4_ASAP7_75t_L g1746 ( 
.A(n_1690),
.B(n_1492),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1659),
.B(n_1581),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1676),
.B(n_1615),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1637),
.Y(n_1749)
);

OAI22xp5_ASAP7_75t_SL g1750 ( 
.A1(n_1622),
.A2(n_1578),
.B1(n_1517),
.B2(n_1591),
.Y(n_1750)
);

AOI221xp5_ASAP7_75t_L g1751 ( 
.A1(n_1684),
.A2(n_1601),
.B1(n_1501),
.B2(n_1612),
.C(n_1518),
.Y(n_1751)
);

AO21x2_ASAP7_75t_L g1752 ( 
.A1(n_1673),
.A2(n_1618),
.B(n_1514),
.Y(n_1752)
);

INVx5_ASAP7_75t_SL g1753 ( 
.A(n_1654),
.Y(n_1753)
);

AOI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1647),
.A2(n_1619),
.B(n_1544),
.Y(n_1754)
);

OAI31xp33_ASAP7_75t_SL g1755 ( 
.A1(n_1666),
.A2(n_1519),
.A3(n_1619),
.B(n_1544),
.Y(n_1755)
);

OAI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1622),
.A2(n_1609),
.B(n_1510),
.Y(n_1756)
);

INVxp67_ASAP7_75t_L g1757 ( 
.A(n_1677),
.Y(n_1757)
);

AOI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1666),
.A2(n_1595),
.B1(n_1610),
.B2(n_1619),
.Y(n_1758)
);

INVx3_ASAP7_75t_L g1759 ( 
.A(n_1625),
.Y(n_1759)
);

OAI211xp5_ASAP7_75t_L g1760 ( 
.A1(n_1634),
.A2(n_1655),
.B(n_1703),
.C(n_1706),
.Y(n_1760)
);

AO32x2_ASAP7_75t_L g1761 ( 
.A1(n_1738),
.A2(n_1724),
.A3(n_1721),
.B1(n_1696),
.B2(n_1687),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1649),
.B(n_1739),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1641),
.B(n_1652),
.Y(n_1763)
);

AOI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1669),
.A2(n_1672),
.B(n_1656),
.Y(n_1764)
);

BUFx12f_ASAP7_75t_L g1765 ( 
.A(n_1742),
.Y(n_1765)
);

AO32x1_ASAP7_75t_L g1766 ( 
.A1(n_1678),
.A2(n_1702),
.A3(n_1710),
.B1(n_1711),
.B2(n_1712),
.Y(n_1766)
);

OAI21xp5_ASAP7_75t_L g1767 ( 
.A1(n_1682),
.A2(n_1702),
.B(n_1648),
.Y(n_1767)
);

OR2x6_ASAP7_75t_L g1768 ( 
.A(n_1658),
.B(n_1625),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1629),
.B(n_1736),
.Y(n_1769)
);

INVx4_ASAP7_75t_L g1770 ( 
.A(n_1715),
.Y(n_1770)
);

OAI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1643),
.A2(n_1713),
.B(n_1678),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1637),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1728),
.B(n_1729),
.Y(n_1773)
);

A2O1A1Ixp33_ASAP7_75t_L g1774 ( 
.A1(n_1683),
.A2(n_1737),
.B(n_1731),
.C(n_1694),
.Y(n_1774)
);

AOI211xp5_ASAP7_75t_L g1775 ( 
.A1(n_1683),
.A2(n_1703),
.B(n_1706),
.C(n_1692),
.Y(n_1775)
);

A2O1A1Ixp33_ASAP7_75t_L g1776 ( 
.A1(n_1737),
.A2(n_1731),
.B(n_1695),
.C(n_1727),
.Y(n_1776)
);

AOI221xp5_ASAP7_75t_L g1777 ( 
.A1(n_1716),
.A2(n_1681),
.B1(n_1680),
.B2(n_1669),
.C(n_1692),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1739),
.B(n_1626),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1638),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1639),
.B(n_1640),
.Y(n_1780)
);

NAND2x1_ASAP7_75t_L g1781 ( 
.A(n_1711),
.B(n_1625),
.Y(n_1781)
);

AO32x2_ASAP7_75t_L g1782 ( 
.A1(n_1738),
.A2(n_1721),
.A3(n_1724),
.B1(n_1716),
.B2(n_1691),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1639),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1640),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1730),
.B(n_1690),
.Y(n_1785)
);

O2A1O1Ixp33_ASAP7_75t_SL g1786 ( 
.A1(n_1693),
.A2(n_1742),
.B(n_1708),
.C(n_1654),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1730),
.B(n_1733),
.Y(n_1787)
);

OR2x6_ASAP7_75t_L g1788 ( 
.A(n_1628),
.B(n_1712),
.Y(n_1788)
);

BUFx8_ASAP7_75t_SL g1789 ( 
.A(n_1743),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1628),
.B(n_1715),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1628),
.B(n_1741),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1642),
.Y(n_1792)
);

BUFx2_ASAP7_75t_L g1793 ( 
.A(n_1739),
.Y(n_1793)
);

OA21x2_ASAP7_75t_L g1794 ( 
.A1(n_1688),
.A2(n_1698),
.B(n_1704),
.Y(n_1794)
);

BUFx2_ASAP7_75t_L g1795 ( 
.A(n_1739),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1722),
.B(n_1726),
.Y(n_1796)
);

OAI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1674),
.A2(n_1698),
.B(n_1719),
.Y(n_1797)
);

A2O1A1Ixp33_ASAP7_75t_L g1798 ( 
.A1(n_1719),
.A2(n_1707),
.B(n_1709),
.C(n_1704),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_L g1799 ( 
.A(n_1686),
.B(n_1700),
.Y(n_1799)
);

INVx4_ASAP7_75t_L g1800 ( 
.A(n_1623),
.Y(n_1800)
);

OR2x6_ASAP7_75t_L g1801 ( 
.A(n_1674),
.B(n_1661),
.Y(n_1801)
);

OAI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1734),
.A2(n_1707),
.B1(n_1709),
.B2(n_1714),
.Y(n_1802)
);

O2A1O1Ixp33_ASAP7_75t_L g1803 ( 
.A1(n_1660),
.A2(n_1714),
.B(n_1723),
.C(n_1661),
.Y(n_1803)
);

AO21x1_ASAP7_75t_L g1804 ( 
.A1(n_1653),
.A2(n_1650),
.B(n_1644),
.Y(n_1804)
);

INVx2_ASAP7_75t_SL g1805 ( 
.A(n_1633),
.Y(n_1805)
);

AO22x2_ASAP7_75t_L g1806 ( 
.A1(n_1680),
.A2(n_1681),
.B1(n_1679),
.B2(n_1653),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1627),
.B(n_1667),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1644),
.B(n_1645),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1645),
.B(n_1646),
.Y(n_1809)
);

OA21x2_ASAP7_75t_L g1810 ( 
.A1(n_1624),
.A2(n_1662),
.B(n_1663),
.Y(n_1810)
);

OAI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1734),
.A2(n_1670),
.B(n_1718),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1627),
.B(n_1667),
.Y(n_1812)
);

INVx11_ASAP7_75t_L g1813 ( 
.A(n_1675),
.Y(n_1813)
);

OA21x2_ASAP7_75t_L g1814 ( 
.A1(n_1624),
.A2(n_1663),
.B(n_1662),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1650),
.B(n_1685),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_L g1816 ( 
.A(n_1708),
.B(n_1675),
.Y(n_1816)
);

AO32x2_ASAP7_75t_L g1817 ( 
.A1(n_1721),
.A2(n_1724),
.A3(n_1660),
.B1(n_1699),
.B2(n_1665),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1685),
.B(n_1725),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1817),
.B(n_1701),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_L g1820 ( 
.A1(n_1777),
.A2(n_1720),
.B1(n_1734),
.B2(n_1679),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1804),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1810),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1793),
.B(n_1636),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1749),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1810),
.Y(n_1825)
);

HB1xp67_ASAP7_75t_L g1826 ( 
.A(n_1814),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1817),
.B(n_1761),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1772),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1779),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1761),
.B(n_1668),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1761),
.B(n_1808),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1795),
.B(n_1671),
.Y(n_1832)
);

AOI22xp33_ASAP7_75t_L g1833 ( 
.A1(n_1764),
.A2(n_1720),
.B1(n_1734),
.B2(n_1665),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1783),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1784),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1792),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1767),
.B(n_1815),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1807),
.Y(n_1838)
);

BUFx2_ASAP7_75t_L g1839 ( 
.A(n_1801),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1807),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_SL g1841 ( 
.A(n_1755),
.B(n_1778),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1812),
.Y(n_1842)
);

INVx1_ASAP7_75t_SL g1843 ( 
.A(n_1744),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1763),
.B(n_1635),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1780),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_L g1846 ( 
.A1(n_1802),
.A2(n_1720),
.B1(n_1697),
.B2(n_1699),
.Y(n_1846)
);

INVx4_ASAP7_75t_L g1847 ( 
.A(n_1765),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1809),
.Y(n_1848)
);

BUFx2_ASAP7_75t_L g1849 ( 
.A(n_1801),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1812),
.Y(n_1850)
);

INVx1_ASAP7_75t_SL g1851 ( 
.A(n_1769),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1806),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1782),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1782),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1806),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1782),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1786),
.B(n_1743),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_L g1858 ( 
.A(n_1762),
.B(n_1723),
.Y(n_1858)
);

AOI22xp33_ASAP7_75t_L g1859 ( 
.A1(n_1802),
.A2(n_1697),
.B1(n_1633),
.B2(n_1705),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1773),
.B(n_1651),
.Y(n_1860)
);

INVxp67_ASAP7_75t_L g1861 ( 
.A(n_1818),
.Y(n_1861)
);

AND2x4_ASAP7_75t_L g1862 ( 
.A(n_1791),
.B(n_1664),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1794),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1803),
.B(n_1632),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_SL g1865 ( 
.A(n_1755),
.B(n_1689),
.Y(n_1865)
);

NOR3xp33_ASAP7_75t_L g1866 ( 
.A(n_1821),
.B(n_1756),
.C(n_1750),
.Y(n_1866)
);

INVxp67_ASAP7_75t_L g1867 ( 
.A(n_1821),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1825),
.Y(n_1868)
);

INVx3_ASAP7_75t_SL g1869 ( 
.A(n_1847),
.Y(n_1869)
);

INVx2_ASAP7_75t_SL g1870 ( 
.A(n_1830),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1838),
.B(n_1840),
.Y(n_1871)
);

OAI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1833),
.A2(n_1775),
.B1(n_1756),
.B2(n_1760),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1837),
.B(n_1757),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1837),
.B(n_1787),
.Y(n_1874)
);

HB1xp67_ASAP7_75t_L g1875 ( 
.A(n_1832),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1824),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1824),
.Y(n_1877)
);

OAI21xp33_ASAP7_75t_L g1878 ( 
.A1(n_1827),
.A2(n_1775),
.B(n_1771),
.Y(n_1878)
);

INVx4_ASAP7_75t_L g1879 ( 
.A(n_1847),
.Y(n_1879)
);

AND2x4_ASAP7_75t_L g1880 ( 
.A(n_1830),
.B(n_1788),
.Y(n_1880)
);

INVx3_ASAP7_75t_L g1881 ( 
.A(n_1862),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1845),
.B(n_1771),
.Y(n_1882)
);

OAI221xp5_ASAP7_75t_L g1883 ( 
.A1(n_1833),
.A2(n_1751),
.B1(n_1750),
.B2(n_1745),
.C(n_1774),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1863),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1831),
.B(n_1785),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1845),
.B(n_1811),
.Y(n_1886)
);

BUFx2_ASAP7_75t_L g1887 ( 
.A(n_1862),
.Y(n_1887)
);

NAND2x1p5_ASAP7_75t_L g1888 ( 
.A(n_1865),
.B(n_1770),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1828),
.Y(n_1889)
);

INVx3_ASAP7_75t_L g1890 ( 
.A(n_1862),
.Y(n_1890)
);

OAI221xp5_ASAP7_75t_L g1891 ( 
.A1(n_1820),
.A2(n_1811),
.B1(n_1776),
.B2(n_1797),
.C(n_1798),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1845),
.B(n_1748),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1828),
.Y(n_1893)
);

OR2x2_ASAP7_75t_L g1894 ( 
.A(n_1848),
.B(n_1797),
.Y(n_1894)
);

NAND4xp25_ASAP7_75t_SL g1895 ( 
.A(n_1827),
.B(n_1758),
.C(n_1754),
.D(n_1753),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1831),
.B(n_1747),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1829),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1829),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1863),
.Y(n_1899)
);

BUFx2_ASAP7_75t_L g1900 ( 
.A(n_1862),
.Y(n_1900)
);

HB1xp67_ASAP7_75t_L g1901 ( 
.A(n_1832),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1851),
.B(n_1788),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1834),
.Y(n_1903)
);

INVx4_ASAP7_75t_L g1904 ( 
.A(n_1847),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1838),
.B(n_1631),
.Y(n_1905)
);

HB1xp67_ASAP7_75t_L g1906 ( 
.A(n_1823),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1863),
.Y(n_1907)
);

INVx3_ASAP7_75t_L g1908 ( 
.A(n_1862),
.Y(n_1908)
);

NAND4xp25_ASAP7_75t_L g1909 ( 
.A(n_1857),
.B(n_1816),
.C(n_1758),
.D(n_1759),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1834),
.Y(n_1910)
);

AOI221xp5_ASAP7_75t_SL g1911 ( 
.A1(n_1827),
.A2(n_1796),
.B1(n_1725),
.B2(n_1735),
.C(n_1732),
.Y(n_1911)
);

OAI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1864),
.A2(n_1768),
.B(n_1781),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1835),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1822),
.Y(n_1914)
);

OAI31xp33_ASAP7_75t_L g1915 ( 
.A1(n_1820),
.A2(n_1746),
.A3(n_1766),
.B(n_1790),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1835),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1836),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1822),
.Y(n_1918)
);

OAI22xp5_ASAP7_75t_L g1919 ( 
.A1(n_1846),
.A2(n_1768),
.B1(n_1753),
.B2(n_1800),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1906),
.B(n_1840),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1906),
.B(n_1875),
.Y(n_1921)
);

NOR2x1_ASAP7_75t_L g1922 ( 
.A(n_1879),
.B(n_1847),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1901),
.B(n_1842),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1911),
.B(n_1842),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1876),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1868),
.Y(n_1926)
);

BUFx3_ASAP7_75t_L g1927 ( 
.A(n_1869),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1876),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1885),
.B(n_1843),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1885),
.B(n_1843),
.Y(n_1930)
);

AND2x4_ASAP7_75t_SL g1931 ( 
.A(n_1902),
.B(n_1847),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1870),
.B(n_1861),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1877),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1877),
.Y(n_1934)
);

AND2x4_ASAP7_75t_L g1935 ( 
.A(n_1880),
.B(n_1839),
.Y(n_1935)
);

BUFx4f_ASAP7_75t_SL g1936 ( 
.A(n_1869),
.Y(n_1936)
);

NOR2x1_ASAP7_75t_L g1937 ( 
.A(n_1879),
.B(n_1904),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1889),
.Y(n_1938)
);

NAND2x1_ASAP7_75t_SL g1939 ( 
.A(n_1869),
.B(n_1819),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1870),
.B(n_1861),
.Y(n_1940)
);

OR2x2_ASAP7_75t_L g1941 ( 
.A(n_1871),
.B(n_1844),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1911),
.B(n_1850),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1889),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1893),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1870),
.B(n_1860),
.Y(n_1945)
);

INVx1_ASAP7_75t_SL g1946 ( 
.A(n_1892),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1893),
.Y(n_1947)
);

NOR2xp33_ASAP7_75t_L g1948 ( 
.A(n_1879),
.B(n_1789),
.Y(n_1948)
);

NOR4xp25_ASAP7_75t_SL g1949 ( 
.A(n_1878),
.B(n_1841),
.C(n_1849),
.D(n_1839),
.Y(n_1949)
);

HB1xp67_ASAP7_75t_L g1950 ( 
.A(n_1871),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1887),
.B(n_1860),
.Y(n_1951)
);

NOR2xp67_ASAP7_75t_L g1952 ( 
.A(n_1895),
.B(n_1826),
.Y(n_1952)
);

INVxp67_ASAP7_75t_SL g1953 ( 
.A(n_1867),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1897),
.Y(n_1954)
);

BUFx3_ASAP7_75t_L g1955 ( 
.A(n_1879),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1887),
.B(n_1860),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1868),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1897),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1900),
.B(n_1874),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1873),
.B(n_1850),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1884),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1873),
.B(n_1823),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1898),
.Y(n_1963)
);

AOI21xp5_ASAP7_75t_L g1964 ( 
.A1(n_1872),
.A2(n_1878),
.B(n_1895),
.Y(n_1964)
);

OR2x2_ASAP7_75t_L g1965 ( 
.A(n_1892),
.B(n_1844),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1898),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1903),
.Y(n_1967)
);

OR2x2_ASAP7_75t_L g1968 ( 
.A(n_1882),
.B(n_1844),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1925),
.Y(n_1969)
);

OAI22xp5_ASAP7_75t_L g1970 ( 
.A1(n_1964),
.A2(n_1872),
.B1(n_1883),
.B2(n_1866),
.Y(n_1970)
);

INVx3_ASAP7_75t_L g1971 ( 
.A(n_1927),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1925),
.Y(n_1972)
);

OR2x2_ASAP7_75t_L g1973 ( 
.A(n_1924),
.B(n_1867),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1928),
.Y(n_1974)
);

NOR2xp33_ASAP7_75t_L g1975 ( 
.A(n_1948),
.B(n_1813),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1928),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1933),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1959),
.B(n_1900),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1933),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1959),
.B(n_1881),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1926),
.Y(n_1981)
);

OR2x2_ASAP7_75t_L g1982 ( 
.A(n_1942),
.B(n_1905),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1953),
.B(n_1866),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1934),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1950),
.B(n_1903),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1921),
.B(n_1910),
.Y(n_1986)
);

HB1xp67_ASAP7_75t_L g1987 ( 
.A(n_1934),
.Y(n_1987)
);

OR2x2_ASAP7_75t_L g1988 ( 
.A(n_1941),
.B(n_1905),
.Y(n_1988)
);

OR2x2_ASAP7_75t_L g1989 ( 
.A(n_1941),
.B(n_1910),
.Y(n_1989)
);

AND2x4_ASAP7_75t_L g1990 ( 
.A(n_1927),
.B(n_1904),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1931),
.B(n_1881),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1931),
.B(n_1881),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1931),
.B(n_1932),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1938),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1938),
.Y(n_1995)
);

BUFx2_ASAP7_75t_L g1996 ( 
.A(n_1939),
.Y(n_1996)
);

OR2x2_ASAP7_75t_L g1997 ( 
.A(n_1968),
.B(n_1913),
.Y(n_1997)
);

OAI31xp33_ASAP7_75t_L g1998 ( 
.A1(n_1949),
.A2(n_1915),
.A3(n_1891),
.B(n_1883),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1932),
.B(n_1881),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1940),
.B(n_1929),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1943),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1943),
.Y(n_2002)
);

INVx4_ASAP7_75t_L g2003 ( 
.A(n_1936),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1940),
.B(n_1890),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1944),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1929),
.B(n_1890),
.Y(n_2006)
);

HB1xp67_ASAP7_75t_L g2007 ( 
.A(n_1944),
.Y(n_2007)
);

INVx4_ASAP7_75t_L g2008 ( 
.A(n_1927),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1962),
.B(n_1913),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1947),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1960),
.B(n_1916),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1947),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1954),
.Y(n_2013)
);

OAI33xp33_ASAP7_75t_L g2014 ( 
.A1(n_1920),
.A2(n_1894),
.A3(n_1886),
.B1(n_1914),
.B2(n_1918),
.B3(n_1917),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1930),
.B(n_1890),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1926),
.Y(n_2016)
);

OR2x6_ASAP7_75t_L g2017 ( 
.A(n_1922),
.B(n_1904),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1930),
.B(n_1951),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1954),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_2018),
.B(n_1955),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1970),
.B(n_1923),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_2000),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1987),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1983),
.B(n_1968),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_2018),
.B(n_1955),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_2007),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1969),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1969),
.Y(n_2028)
);

AND2x4_ASAP7_75t_L g2029 ( 
.A(n_1996),
.B(n_1952),
.Y(n_2029)
);

NAND2x1_ASAP7_75t_L g2030 ( 
.A(n_1996),
.B(n_1922),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1972),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1981),
.Y(n_2032)
);

OR2x2_ASAP7_75t_L g2033 ( 
.A(n_1982),
.B(n_1965),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1972),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_2000),
.B(n_1955),
.Y(n_2035)
);

AND2x4_ASAP7_75t_L g2036 ( 
.A(n_1993),
.B(n_1952),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1982),
.B(n_1965),
.Y(n_2037)
);

AND2x2_ASAP7_75t_SL g2038 ( 
.A(n_2003),
.B(n_1904),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_SL g2039 ( 
.A(n_1998),
.B(n_1935),
.Y(n_2039)
);

HB1xp67_ASAP7_75t_L g2040 ( 
.A(n_1973),
.Y(n_2040)
);

AOI22xp5_ASAP7_75t_L g2041 ( 
.A1(n_2014),
.A2(n_1891),
.B1(n_1752),
.B2(n_1919),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1976),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1993),
.B(n_1951),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1978),
.B(n_1956),
.Y(n_2044)
);

OR2x2_ASAP7_75t_L g2045 ( 
.A(n_1988),
.B(n_1958),
.Y(n_2045)
);

INVxp67_ASAP7_75t_SL g2046 ( 
.A(n_1971),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1981),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1976),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1973),
.B(n_1946),
.Y(n_2049)
);

NOR2xp33_ASAP7_75t_L g2050 ( 
.A(n_2003),
.B(n_1909),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1977),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1977),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_1978),
.B(n_1956),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_1991),
.B(n_1945),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_2016),
.Y(n_2055)
);

NAND4xp25_ASAP7_75t_L g2056 ( 
.A(n_2008),
.B(n_1937),
.C(n_1915),
.D(n_1909),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1979),
.Y(n_2057)
);

INVx1_ASAP7_75t_SL g2058 ( 
.A(n_2003),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_2016),
.Y(n_2059)
);

AOI21xp5_ASAP7_75t_L g2060 ( 
.A1(n_1985),
.A2(n_1912),
.B(n_1937),
.Y(n_2060)
);

O2A1O1Ixp33_ASAP7_75t_L g2061 ( 
.A1(n_2039),
.A2(n_1971),
.B(n_1984),
.C(n_1979),
.Y(n_2061)
);

AOI221xp5_ASAP7_75t_SL g2062 ( 
.A1(n_2056),
.A2(n_1971),
.B1(n_1980),
.B2(n_2004),
.C(n_1999),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_2022),
.Y(n_2063)
);

OAI221xp5_ASAP7_75t_SL g2064 ( 
.A1(n_2041),
.A2(n_1997),
.B1(n_1853),
.B2(n_1856),
.C(n_1854),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_2044),
.B(n_1990),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_SL g2066 ( 
.A(n_2029),
.B(n_2008),
.Y(n_2066)
);

AOI32xp33_ASAP7_75t_L g2067 ( 
.A1(n_2029),
.A2(n_1856),
.A3(n_1854),
.B1(n_1853),
.B2(n_1914),
.Y(n_2067)
);

OR2x2_ASAP7_75t_L g2068 ( 
.A(n_2033),
.B(n_2024),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2027),
.Y(n_2069)
);

INVxp67_ASAP7_75t_L g2070 ( 
.A(n_2050),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_2040),
.B(n_2008),
.Y(n_2071)
);

OR2x2_ASAP7_75t_L g2072 ( 
.A(n_2022),
.B(n_1986),
.Y(n_2072)
);

AOI22xp5_ASAP7_75t_L g2073 ( 
.A1(n_2041),
.A2(n_1854),
.B1(n_1853),
.B2(n_1856),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_2021),
.B(n_1988),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2027),
.Y(n_2075)
);

OAI22xp5_ASAP7_75t_L g2076 ( 
.A1(n_2036),
.A2(n_1935),
.B1(n_2017),
.B2(n_1888),
.Y(n_2076)
);

OAI32xp33_ASAP7_75t_L g2077 ( 
.A1(n_2033),
.A2(n_1997),
.A3(n_1989),
.B1(n_1888),
.B2(n_1999),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2028),
.Y(n_2078)
);

NAND4xp75_ASAP7_75t_L g2079 ( 
.A(n_2038),
.B(n_1912),
.C(n_1992),
.D(n_1991),
.Y(n_2079)
);

OAI22xp5_ASAP7_75t_L g2080 ( 
.A1(n_2036),
.A2(n_1935),
.B1(n_2017),
.B2(n_1888),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2023),
.B(n_2011),
.Y(n_2081)
);

OAI32xp33_ASAP7_75t_L g2082 ( 
.A1(n_2049),
.A2(n_1989),
.A3(n_2004),
.B1(n_1980),
.B2(n_1992),
.Y(n_2082)
);

INVx2_ASAP7_75t_L g2083 ( 
.A(n_2032),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_2023),
.B(n_2009),
.Y(n_2084)
);

OAI22xp33_ASAP7_75t_SL g2085 ( 
.A1(n_2029),
.A2(n_1855),
.B1(n_1852),
.B2(n_1882),
.Y(n_2085)
);

AOI211xp5_ASAP7_75t_L g2086 ( 
.A1(n_2029),
.A2(n_1919),
.B(n_1990),
.C(n_2019),
.Y(n_2086)
);

HB1xp67_ASAP7_75t_L g2087 ( 
.A(n_2028),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_2032),
.Y(n_2088)
);

AOI21xp33_ASAP7_75t_SL g2089 ( 
.A1(n_2061),
.A2(n_2038),
.B(n_2036),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_2065),
.B(n_2058),
.Y(n_2090)
);

AOI222xp33_ASAP7_75t_L g2091 ( 
.A1(n_2074),
.A2(n_2036),
.B1(n_2059),
.B2(n_2032),
.C1(n_2055),
.C2(n_2047),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2087),
.Y(n_2092)
);

OAI21xp5_ASAP7_75t_SL g2093 ( 
.A1(n_2065),
.A2(n_2035),
.B(n_2025),
.Y(n_2093)
);

NOR2xp33_ASAP7_75t_L g2094 ( 
.A(n_2070),
.B(n_2038),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2087),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_SL g2096 ( 
.A(n_2062),
.B(n_2046),
.Y(n_2096)
);

NAND4xp25_ASAP7_75t_L g2097 ( 
.A(n_2086),
.B(n_2026),
.C(n_2035),
.D(n_2060),
.Y(n_2097)
);

OAI22xp5_ASAP7_75t_SL g2098 ( 
.A1(n_2068),
.A2(n_2030),
.B1(n_2026),
.B2(n_1975),
.Y(n_2098)
);

AOI22xp5_ASAP7_75t_L g2099 ( 
.A1(n_2073),
.A2(n_2059),
.B1(n_2055),
.B2(n_2047),
.Y(n_2099)
);

OAI21xp5_ASAP7_75t_L g2100 ( 
.A1(n_2064),
.A2(n_2030),
.B(n_2025),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_2068),
.B(n_2020),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2063),
.B(n_2044),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2063),
.Y(n_2103)
);

AOI211xp5_ASAP7_75t_L g2104 ( 
.A1(n_2077),
.A2(n_2031),
.B(n_2057),
.C(n_2042),
.Y(n_2104)
);

NAND3xp33_ASAP7_75t_L g2105 ( 
.A(n_2071),
.B(n_2066),
.C(n_2067),
.Y(n_2105)
);

OAI21xp33_ASAP7_75t_L g2106 ( 
.A1(n_2082),
.A2(n_2020),
.B(n_2037),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2072),
.B(n_2053),
.Y(n_2107)
);

NOR2xp33_ASAP7_75t_L g2108 ( 
.A(n_2066),
.B(n_2043),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_2079),
.B(n_2053),
.Y(n_2109)
);

AOI322xp5_ASAP7_75t_L g2110 ( 
.A1(n_2083),
.A2(n_2059),
.A3(n_2055),
.B1(n_2057),
.B2(n_2031),
.C1(n_2052),
.C2(n_2051),
.Y(n_2110)
);

OAI31xp33_ASAP7_75t_L g2111 ( 
.A1(n_2085),
.A2(n_2034),
.A3(n_2052),
.B(n_2051),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2101),
.B(n_2043),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2107),
.Y(n_2113)
);

AOI22xp5_ASAP7_75t_L g2114 ( 
.A1(n_2099),
.A2(n_2088),
.B1(n_2083),
.B2(n_2080),
.Y(n_2114)
);

AOI21xp33_ASAP7_75t_L g2115 ( 
.A1(n_2091),
.A2(n_2088),
.B(n_2075),
.Y(n_2115)
);

INVxp67_ASAP7_75t_L g2116 ( 
.A(n_2094),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2107),
.Y(n_2117)
);

OAI21xp33_ASAP7_75t_L g2118 ( 
.A1(n_2097),
.A2(n_2084),
.B(n_2081),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2102),
.Y(n_2119)
);

NOR2x1_ASAP7_75t_L g2120 ( 
.A(n_2092),
.B(n_2069),
.Y(n_2120)
);

OAI22xp5_ASAP7_75t_L g2121 ( 
.A1(n_2098),
.A2(n_2076),
.B1(n_2045),
.B2(n_2054),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_SL g2122 ( 
.A(n_2111),
.B(n_1990),
.Y(n_2122)
);

NOR2xp67_ASAP7_75t_SL g2123 ( 
.A(n_2090),
.B(n_1633),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2095),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_2103),
.Y(n_2125)
);

INVx1_ASAP7_75t_SL g2126 ( 
.A(n_2109),
.Y(n_2126)
);

NAND4xp75_ASAP7_75t_L g2127 ( 
.A(n_2120),
.B(n_2096),
.C(n_2094),
.D(n_2100),
.Y(n_2127)
);

AOI221xp5_ASAP7_75t_L g2128 ( 
.A1(n_2115),
.A2(n_2096),
.B1(n_2105),
.B2(n_2089),
.C(n_2104),
.Y(n_2128)
);

INVxp33_ASAP7_75t_L g2129 ( 
.A(n_2112),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_2126),
.B(n_2108),
.Y(n_2130)
);

NOR2xp33_ASAP7_75t_L g2131 ( 
.A(n_2123),
.B(n_2093),
.Y(n_2131)
);

NAND3xp33_ASAP7_75t_L g2132 ( 
.A(n_2116),
.B(n_2110),
.C(n_2108),
.Y(n_2132)
);

HB1xp67_ASAP7_75t_L g2133 ( 
.A(n_2113),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_2117),
.B(n_2106),
.Y(n_2134)
);

OAI221xp5_ASAP7_75t_L g2135 ( 
.A1(n_2114),
.A2(n_2078),
.B1(n_1939),
.B2(n_2048),
.C(n_2034),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2125),
.Y(n_2136)
);

AOI221xp5_ASAP7_75t_SL g2137 ( 
.A1(n_2122),
.A2(n_2048),
.B1(n_2042),
.B2(n_2054),
.C(n_2045),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_SL g2138 ( 
.A(n_2121),
.B(n_1935),
.Y(n_2138)
);

OAI221xp5_ASAP7_75t_L g2139 ( 
.A1(n_2128),
.A2(n_2118),
.B1(n_2122),
.B2(n_2116),
.C(n_2125),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2133),
.Y(n_2140)
);

OAI22xp33_ASAP7_75t_L g2141 ( 
.A1(n_2132),
.A2(n_2130),
.B1(n_2135),
.B2(n_2134),
.Y(n_2141)
);

AOI221xp5_ASAP7_75t_L g2142 ( 
.A1(n_2136),
.A2(n_2124),
.B1(n_2119),
.B2(n_1914),
.C(n_1918),
.Y(n_2142)
);

AOI21xp33_ASAP7_75t_SL g2143 ( 
.A1(n_2129),
.A2(n_2017),
.B(n_1805),
.Y(n_2143)
);

AOI221xp5_ASAP7_75t_L g2144 ( 
.A1(n_2137),
.A2(n_1918),
.B1(n_1984),
.B2(n_2013),
.C(n_2012),
.Y(n_2144)
);

AOI22xp5_ASAP7_75t_L g2145 ( 
.A1(n_2127),
.A2(n_1884),
.B1(n_1907),
.B2(n_1899),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2138),
.Y(n_2146)
);

AOI22xp5_ASAP7_75t_L g2147 ( 
.A1(n_2131),
.A2(n_1907),
.B1(n_1899),
.B2(n_1858),
.Y(n_2147)
);

OAI221xp5_ASAP7_75t_L g2148 ( 
.A1(n_2139),
.A2(n_2017),
.B1(n_2019),
.B2(n_2010),
.C(n_2013),
.Y(n_2148)
);

OAI221xp5_ASAP7_75t_L g2149 ( 
.A1(n_2142),
.A2(n_2147),
.B1(n_2140),
.B2(n_2145),
.C(n_2146),
.Y(n_2149)
);

OAI21xp5_ASAP7_75t_L g2150 ( 
.A1(n_2141),
.A2(n_1995),
.B(n_1994),
.Y(n_2150)
);

AOI221xp5_ASAP7_75t_L g2151 ( 
.A1(n_2144),
.A2(n_2143),
.B1(n_2012),
.B2(n_2010),
.C(n_2005),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2140),
.Y(n_2152)
);

OAI211xp5_ASAP7_75t_L g2153 ( 
.A1(n_2139),
.A2(n_1995),
.B(n_1994),
.C(n_2005),
.Y(n_2153)
);

AOI221xp5_ASAP7_75t_L g2154 ( 
.A1(n_2141),
.A2(n_2002),
.B1(n_2001),
.B2(n_1974),
.C(n_1899),
.Y(n_2154)
);

AOI222xp33_ASAP7_75t_L g2155 ( 
.A1(n_2139),
.A2(n_1926),
.B1(n_1957),
.B2(n_1855),
.C1(n_1852),
.C2(n_2002),
.Y(n_2155)
);

NOR2x1p5_ASAP7_75t_L g2156 ( 
.A(n_2152),
.B(n_1633),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_2155),
.B(n_2006),
.Y(n_2157)
);

XNOR2xp5_ASAP7_75t_L g2158 ( 
.A(n_2149),
.B(n_1717),
.Y(n_2158)
);

AOI22xp5_ASAP7_75t_L g2159 ( 
.A1(n_2154),
.A2(n_1957),
.B1(n_2006),
.B2(n_2015),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_2148),
.Y(n_2160)
);

NAND4xp75_ASAP7_75t_L g2161 ( 
.A(n_2150),
.B(n_2015),
.C(n_1858),
.D(n_1902),
.Y(n_2161)
);

AOI22xp5_ASAP7_75t_L g2162 ( 
.A1(n_2153),
.A2(n_2151),
.B1(n_1957),
.B2(n_1907),
.Y(n_2162)
);

NOR2xp33_ASAP7_75t_L g2163 ( 
.A(n_2157),
.B(n_1958),
.Y(n_2163)
);

NAND3xp33_ASAP7_75t_L g2164 ( 
.A(n_2160),
.B(n_1966),
.C(n_1963),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2161),
.B(n_1967),
.Y(n_2165)
);

INVxp67_ASAP7_75t_L g2166 ( 
.A(n_2156),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_2159),
.B(n_1945),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2167),
.B(n_2158),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2165),
.Y(n_2169)
);

OAI22x1_ASAP7_75t_L g2170 ( 
.A1(n_2169),
.A2(n_2166),
.B1(n_2163),
.B2(n_2164),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2170),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2170),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_2171),
.Y(n_2173)
);

OAI21xp33_ASAP7_75t_L g2174 ( 
.A1(n_2172),
.A2(n_2168),
.B(n_2162),
.Y(n_2174)
);

AOI21xp5_ASAP7_75t_L g2175 ( 
.A1(n_2174),
.A2(n_1896),
.B(n_1963),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_2175),
.B(n_2173),
.Y(n_2176)
);

NAND2xp67_ASAP7_75t_L g2177 ( 
.A(n_2176),
.B(n_1896),
.Y(n_2177)
);

INVxp67_ASAP7_75t_L g2178 ( 
.A(n_2177),
.Y(n_2178)
);

OAI221xp5_ASAP7_75t_R g2179 ( 
.A1(n_2178),
.A2(n_1967),
.B1(n_1966),
.B2(n_1859),
.C(n_1908),
.Y(n_2179)
);

AOI211xp5_ASAP7_75t_L g2180 ( 
.A1(n_2179),
.A2(n_1799),
.B(n_1740),
.C(n_1961),
.Y(n_2180)
);


endmodule