module fake_jpeg_21546_n_256 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_256);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx8_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_28),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

CKINVDCx9p33_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_32),
.Y(n_35)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_28),
.A2(n_13),
.B1(n_21),
.B2(n_24),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_34),
.A2(n_21),
.B1(n_13),
.B2(n_24),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_11),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_13),
.Y(n_53)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_23),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_53),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_53),
.Y(n_78)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_54),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_33),
.B1(n_26),
.B2(n_29),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_35),
.B1(n_38),
.B2(n_24),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_56),
.A2(n_60),
.B1(n_35),
.B2(n_21),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_14),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_57),
.B(n_59),
.Y(n_72)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_17),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_31),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_34),
.B1(n_35),
.B2(n_42),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_35),
.B1(n_38),
.B2(n_12),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_61),
.A2(n_42),
.B1(n_21),
.B2(n_13),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_60),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_61),
.A2(n_21),
.B1(n_24),
.B2(n_41),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_50),
.B1(n_61),
.B2(n_45),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_79),
.B(n_11),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_74),
.B1(n_49),
.B2(n_58),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_25),
.B1(n_38),
.B2(n_35),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_48),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_80),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_19),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_60),
.A2(n_11),
.B1(n_14),
.B2(n_23),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_30),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_78),
.Y(n_109)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_55),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_88),
.C(n_71),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_44),
.B1(n_14),
.B2(n_23),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_87),
.B(n_92),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_17),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_75),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_72),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_12),
.B(n_17),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_77),
.B1(n_74),
.B2(n_73),
.Y(n_106)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_93),
.B(n_49),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_63),
.B(n_16),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_95),
.B(n_96),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_69),
.B(n_16),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_97),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_94),
.A2(n_68),
.B1(n_62),
.B2(n_77),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_99),
.A2(n_106),
.B1(n_113),
.B2(n_18),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_94),
.A2(n_69),
.B(n_77),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_102),
.B(n_116),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_69),
.B(n_77),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_104),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_72),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_108),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_84),
.B(n_78),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_111),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_70),
.Y(n_112)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_92),
.A2(n_70),
.B1(n_79),
.B2(n_67),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_93),
.A2(n_67),
.B1(n_54),
.B2(n_65),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_66),
.Y(n_117)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_88),
.C(n_82),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_120),
.B(n_136),
.C(n_19),
.Y(n_162)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_126),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_83),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_129),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_90),
.B(n_97),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_110),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_110),
.Y(n_127)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_82),
.B(n_86),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_130),
.B(n_119),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_91),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_65),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_134),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_65),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_43),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_135),
.B(n_16),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_43),
.C(n_19),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_100),
.A2(n_17),
.B(n_18),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_140),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_17),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_43),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_114),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_118),
.B1(n_115),
.B2(n_117),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_118),
.A2(n_101),
.B(n_98),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_18),
.Y(n_156)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_143),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_147),
.B(n_1),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_129),
.A2(n_118),
.B1(n_98),
.B2(n_106),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_150),
.A2(n_153),
.B1(n_158),
.B2(n_159),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_125),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_151),
.B(n_157),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_119),
.A2(n_107),
.B(n_85),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_136),
.B(n_1),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_156),
.A2(n_18),
.B(n_16),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_22),
.B1(n_20),
.B2(n_15),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_162),
.C(n_163),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_16),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_161),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_120),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_132),
.A2(n_22),
.B1(n_20),
.B2(n_15),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_15),
.Y(n_185)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_140),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_138),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_135),
.Y(n_169)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

NOR4xp25_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_133),
.C(n_123),
.D(n_128),
.Y(n_175)
);

INVxp67_ASAP7_75t_SL g195 ( 
.A(n_175),
.Y(n_195)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_180),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_178),
.A2(n_179),
.B(n_156),
.Y(n_189)
);

BUFx12f_ASAP7_75t_SL g179 ( 
.A(n_144),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_155),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_0),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_181),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_0),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_182),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_186),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_0),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_184),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_185),
.A2(n_159),
.B1(n_162),
.B2(n_144),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_189),
.A2(n_183),
.B(n_188),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_190),
.A2(n_172),
.B1(n_180),
.B2(n_168),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_163),
.C(n_148),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_193),
.C(n_201),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_154),
.C(n_160),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_179),
.B(n_147),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_186),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_180),
.A2(n_154),
.B(n_157),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_199),
.B(n_1),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_169),
.C(n_174),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_195),
.C(n_193),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_209),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_204),
.A2(n_210),
.B1(n_211),
.B2(n_197),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_171),
.Y(n_205)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_171),
.Y(n_206)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_207),
.B(n_200),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_178),
.C(n_174),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_212),
.C(n_199),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_176),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_196),
.A2(n_185),
.B1(n_168),
.B2(n_22),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_19),
.C(n_20),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_213),
.A2(n_188),
.B(n_194),
.Y(n_219)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_216),
.Y(n_227)
);

OA21x2_ASAP7_75t_L g216 ( 
.A1(n_206),
.A2(n_198),
.B(n_189),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_4),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_200),
.C(n_22),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_223),
.C(n_212),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_222),
.B(n_207),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_20),
.C(n_16),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_208),
.A2(n_2),
.B(n_3),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_224),
.A2(n_2),
.B(n_4),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_222),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_229),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_16),
.C(n_3),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_230),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_4),
.C(n_5),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_216),
.Y(n_236)
);

NOR2xp67_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_5),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_232),
.A2(n_220),
.B(n_216),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_227),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_236),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_235),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_214),
.C(n_223),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_238),
.B(n_240),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_5),
.Y(n_245)
);

OAI21x1_ASAP7_75t_L g242 ( 
.A1(n_236),
.A2(n_225),
.B(n_6),
.Y(n_242)
);

AOI21xp33_ASAP7_75t_L g248 ( 
.A1(n_242),
.A2(n_245),
.B(n_6),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_239),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_247),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_248),
.A2(n_246),
.B(n_7),
.Y(n_249)
);

OAI21x1_ASAP7_75t_SL g251 ( 
.A1(n_249),
.A2(n_244),
.B(n_237),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_250),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_6),
.C(n_7),
.Y(n_253)
);

MAJx2_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_7),
.C(n_8),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_254),
.A2(n_8),
.B(n_9),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_8),
.C(n_10),
.Y(n_256)
);


endmodule