module fake_jpeg_3588_n_293 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_293);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_293;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_241;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_13),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_41),
.B(n_44),
.Y(n_81)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_51),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_28),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_0),
.Y(n_58)
);

AOI21xp33_ASAP7_75t_L g94 ( 
.A1(n_58),
.A2(n_25),
.B(n_18),
.Y(n_94)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g104 ( 
.A(n_60),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_24),
.B1(n_34),
.B2(n_35),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_62),
.A2(n_70),
.B1(n_71),
.B2(n_101),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_54),
.A2(n_19),
.B1(n_31),
.B2(n_40),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_64),
.A2(n_80),
.B1(n_83),
.B2(n_88),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_58),
.A2(n_24),
.B1(n_34),
.B2(n_35),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_24),
.B1(n_34),
.B2(n_32),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_27),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_73),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_44),
.B(n_27),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_31),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_78),
.B(n_94),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_32),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_84),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_53),
.A2(n_26),
.B1(n_37),
.B2(n_21),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_53),
.A2(n_40),
.B1(n_37),
.B2(n_22),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_22),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_30),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_87),
.Y(n_122)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_53),
.A2(n_50),
.B1(n_26),
.B2(n_29),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_30),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_90),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_29),
.Y(n_90)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_60),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_96),
.Y(n_127)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_25),
.Y(n_96)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_55),
.A2(n_18),
.B1(n_36),
.B2(n_20),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_20),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_48),
.B(n_17),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_106),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_52),
.A2(n_18),
.B1(n_36),
.B2(n_20),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_52),
.A2(n_18),
.B1(n_36),
.B2(n_20),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_121)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx3_ASAP7_75t_SL g167 ( 
.A(n_107),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_124),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_110),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_20),
.C(n_2),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_112),
.B(n_132),
.C(n_74),
.Y(n_158)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_17),
.B(n_16),
.C(n_15),
.Y(n_116)
);

AOI21xp33_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_99),
.B(n_10),
.Y(n_143)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_82),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_76),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_98),
.A2(n_4),
.B(n_5),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_125),
.Y(n_168)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_90),
.A2(n_6),
.B(n_8),
.C(n_9),
.Y(n_128)
);

O2A1O1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_128),
.A2(n_82),
.B(n_11),
.C(n_12),
.Y(n_165)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_72),
.B(n_14),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_131),
.B(n_9),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_78),
.B(n_6),
.Y(n_132)
);

BUFx10_ASAP7_75t_L g133 ( 
.A(n_69),
.Y(n_133)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_78),
.B(n_8),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_137),
.B(n_105),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_138),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_139),
.B(n_150),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_117),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_142),
.B(n_148),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_143),
.B(n_157),
.Y(n_191)
);

AO22x1_ASAP7_75t_SL g147 ( 
.A1(n_118),
.A2(n_77),
.B1(n_68),
.B2(n_104),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_158),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_68),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_77),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_152),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_115),
.A2(n_91),
.B1(n_104),
.B2(n_74),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_153),
.A2(n_161),
.B1(n_170),
.B2(n_107),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_97),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_66),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_163),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_115),
.A2(n_63),
.B1(n_95),
.B2(n_92),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_162),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_102),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_127),
.A2(n_105),
.B1(n_63),
.B2(n_65),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_164),
.A2(n_111),
.B(n_123),
.Y(n_176)
);

OAI21x1_ASAP7_75t_SL g186 ( 
.A1(n_165),
.A2(n_133),
.B(n_137),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_112),
.B(n_65),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_130),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_109),
.A2(n_67),
.B1(n_102),
.B2(n_12),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_171),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_168),
.A2(n_125),
.B(n_109),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_175),
.A2(n_176),
.B(n_183),
.Y(n_205)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_177),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_160),
.A2(n_132),
.B1(n_119),
.B2(n_113),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_178),
.A2(n_192),
.B1(n_193),
.B2(n_167),
.Y(n_217)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_179),
.B(n_182),
.Y(n_203)
);

BUFx12_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_180),
.Y(n_201)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_154),
.A2(n_128),
.B(n_116),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_184),
.B(n_189),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_163),
.A2(n_132),
.B1(n_129),
.B2(n_67),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_185),
.A2(n_166),
.B1(n_151),
.B2(n_170),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_164),
.Y(n_204)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_190),
.B(n_153),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_161),
.A2(n_120),
.B1(n_108),
.B2(n_110),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_154),
.A2(n_134),
.B(n_108),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_194),
.A2(n_155),
.B(n_134),
.Y(n_218)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_144),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_195),
.B(n_171),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_149),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_199),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_149),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_176),
.A2(n_154),
.B(n_165),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_200),
.A2(n_204),
.B(n_218),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_207),
.A2(n_212),
.B1(n_217),
.B2(n_199),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_158),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_208),
.B(n_210),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_181),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_175),
.C(n_185),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_182),
.A2(n_156),
.B1(n_167),
.B2(n_110),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_172),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_214),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_173),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_184),
.A2(n_181),
.B1(n_187),
.B2(n_188),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_220),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_155),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_219),
.B(n_179),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_174),
.Y(n_220)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_221),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_227),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_202),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_225),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_196),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_187),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_228),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_205),
.A2(n_200),
.B(n_204),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_194),
.C(n_178),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_205),
.A2(n_183),
.B(n_191),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_238),
.Y(n_248)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_234),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_235),
.A2(n_211),
.B1(n_215),
.B2(n_210),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_216),
.B(n_177),
.Y(n_236)
);

XNOR2x1_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_211),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_203),
.Y(n_237)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_237),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_214),
.B(n_196),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_239),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_207),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_251),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_239),
.A2(n_220),
.B1(n_206),
.B2(n_212),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_247),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_231),
.A2(n_156),
.B1(n_186),
.B2(n_215),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_252),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_232),
.A2(n_229),
.B1(n_231),
.B2(n_233),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_236),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_L g252 ( 
.A1(n_224),
.A2(n_201),
.B1(n_198),
.B2(n_197),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_254),
.A2(n_247),
.B1(n_246),
.B2(n_251),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_222),
.C(n_228),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_259),
.Y(n_271)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_257),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_230),
.C(n_227),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_230),
.C(n_201),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_261),
.C(n_244),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_224),
.C(n_195),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_189),
.Y(n_262)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_262),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_253),
.Y(n_264)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_264),
.Y(n_269)
);

NOR2xp67_ASAP7_75t_SL g277 ( 
.A(n_266),
.B(n_180),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_258),
.A2(n_255),
.B1(n_254),
.B2(n_264),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_169),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_252),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_270),
.B(n_272),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_120),
.C(n_169),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_180),
.C(n_152),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_145),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_274),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_275),
.A2(n_277),
.B(n_279),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_135),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_271),
.A2(n_145),
.B(n_180),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_280),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_266),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_273),
.C(n_270),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_278),
.B(n_265),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_284),
.B(n_268),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_287),
.Y(n_289)
);

AOI322xp5_ASAP7_75t_L g288 ( 
.A1(n_286),
.A2(n_281),
.A3(n_283),
.B1(n_267),
.B2(n_282),
.C1(n_146),
.C2(n_133),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_288),
.B(n_289),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_133),
.B(n_11),
.Y(n_291)
);

OAI21xp33_ASAP7_75t_SL g292 ( 
.A1(n_291),
.A2(n_10),
.B(n_13),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_13),
.Y(n_293)
);


endmodule