module fake_jpeg_14093_n_618 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_618);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_618;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_6),
.B(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_18),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_11),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_16),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_62),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_63),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_31),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_64),
.B(n_80),
.Y(n_144)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_68),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_36),
.B(n_0),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_69),
.B(n_74),
.Y(n_211)
);

INVx11_ASAP7_75t_SL g70 ( 
.A(n_60),
.Y(n_70)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_70),
.Y(n_150)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_71),
.Y(n_139)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_72),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_73),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_36),
.B(n_0),
.Y(n_74)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_75),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_76),
.Y(n_154)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_78),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_79),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_31),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_81),
.Y(n_152)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_82),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_83),
.Y(n_175)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_84),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_85),
.Y(n_156)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_86),
.Y(n_188)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_87),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_88),
.Y(n_187)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_90),
.Y(n_191)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_91),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_31),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_92),
.B(n_108),
.Y(n_160)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_93),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_25),
.Y(n_94)
);

NAND2x1_ASAP7_75t_SL g132 ( 
.A(n_94),
.B(n_34),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_95),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_19),
.Y(n_97)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_27),
.B(n_0),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_98),
.B(n_105),
.Y(n_129)
);

BUFx12_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

BUFx4f_ASAP7_75t_SL g190 ( 
.A(n_99),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_100),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_29),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_101),
.B(n_57),
.Y(n_143)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_19),
.Y(n_103)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_103),
.Y(n_158)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_104),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_27),
.B(n_3),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_29),
.Y(n_106)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_29),
.Y(n_107)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_107),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_31),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_109),
.Y(n_179)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_26),
.Y(n_110)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_110),
.Y(n_198)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_30),
.Y(n_111)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_111),
.Y(n_199)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_19),
.Y(n_112)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_112),
.Y(n_208)
);

BUFx12_ASAP7_75t_L g113 ( 
.A(n_34),
.Y(n_113)
);

CKINVDCx10_ASAP7_75t_R g159 ( 
.A(n_113),
.Y(n_159)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

INVx3_ASAP7_75t_SL g137 ( 
.A(n_114),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_115),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_116),
.Y(n_178)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_30),
.Y(n_117)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_117),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

INVx3_ASAP7_75t_SL g195 ( 
.A(n_118),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_32),
.B(n_18),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_119),
.B(n_3),
.Y(n_134)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_37),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_120),
.B(n_124),
.Y(n_177)
);

INVx4_ASAP7_75t_SL g121 ( 
.A(n_34),
.Y(n_121)
);

INVx13_ASAP7_75t_L g209 ( 
.A(n_121),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_53),
.Y(n_122)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_123),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_31),
.Y(n_124)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_22),
.Y(n_125)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_125),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_126),
.Y(n_210)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_51),
.Y(n_127)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_127),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_78),
.A2(n_33),
.B1(n_22),
.B2(n_51),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_128),
.A2(n_57),
.B1(n_83),
.B2(n_79),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_132),
.B(n_169),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_134),
.B(n_194),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_70),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_135),
.B(n_145),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_143),
.B(n_153),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_99),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_102),
.B(n_51),
.Y(n_153)
);

INVx2_ASAP7_75t_R g162 ( 
.A(n_121),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_162),
.B(n_196),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_89),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_163),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_113),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_164),
.B(n_167),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_61),
.A2(n_22),
.B1(n_58),
.B2(n_59),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_165),
.A2(n_197),
.B1(n_207),
.B2(n_54),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_75),
.Y(n_167)
);

HAxp5_ASAP7_75t_SL g169 ( 
.A(n_94),
.B(n_60),
.CON(n_169),
.SN(n_169)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_123),
.B(n_37),
.C(n_41),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_180),
.B(n_56),
.C(n_8),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_67),
.B(n_32),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_181),
.B(n_183),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_67),
.B(n_42),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_95),
.B(n_55),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_186),
.B(n_50),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g192 ( 
.A(n_95),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_192),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_106),
.B(n_42),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_127),
.B(n_51),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_114),
.A2(n_43),
.B1(n_59),
.B2(n_44),
.Y(n_197)
);

BUFx10_ASAP7_75t_L g201 ( 
.A(n_116),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_201),
.Y(n_213)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_125),
.Y(n_204)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_204),
.Y(n_212)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_62),
.Y(n_205)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_63),
.A2(n_48),
.B1(n_45),
.B2(n_46),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_177),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_214),
.B(n_245),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_157),
.Y(n_215)
);

INVx6_ASAP7_75t_L g331 ( 
.A(n_215),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_216),
.A2(n_226),
.B1(n_247),
.B2(n_272),
.Y(n_293)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_219),
.Y(n_297)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_221),
.Y(n_300)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_137),
.Y(n_222)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_222),
.Y(n_306)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_223),
.Y(n_294)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_224),
.Y(n_299)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_178),
.Y(n_225)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_225),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_211),
.A2(n_76),
.B1(n_122),
.B2(n_118),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_169),
.A2(n_48),
.B(n_46),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_227),
.A2(n_268),
.B(n_273),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_157),
.Y(n_228)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_228),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_156),
.A2(n_52),
.B1(n_45),
.B2(n_41),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_229),
.Y(n_305)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_166),
.Y(n_231)
);

INVx5_ASAP7_75t_L g335 ( 
.A(n_231),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_156),
.A2(n_52),
.B1(n_93),
.B2(n_126),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_232),
.Y(n_314)
);

INVx11_ASAP7_75t_L g233 ( 
.A(n_147),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_233),
.Y(n_311)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_210),
.Y(n_234)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_234),
.Y(n_312)
);

BUFx16f_ASAP7_75t_L g235 ( 
.A(n_150),
.Y(n_235)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_235),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_132),
.A2(n_100),
.B1(n_51),
.B2(n_57),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_237),
.A2(n_262),
.B1(n_267),
.B2(n_280),
.Y(n_286)
);

AOI21xp33_ASAP7_75t_SL g239 ( 
.A1(n_143),
.A2(n_60),
.B(n_116),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_239),
.B(n_263),
.C(n_258),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_129),
.B(n_43),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_241),
.B(n_256),
.Y(n_336)
);

INVx8_ASAP7_75t_L g242 ( 
.A(n_166),
.Y(n_242)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_242),
.Y(n_329)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_133),
.Y(n_243)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_243),
.Y(n_287)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_210),
.Y(n_244)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_244),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_139),
.B(n_55),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_174),
.Y(n_246)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_246),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_207),
.A2(n_109),
.B1(n_96),
.B2(n_90),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_200),
.Y(n_248)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_248),
.Y(n_310)
);

INVx8_ASAP7_75t_L g249 ( 
.A(n_200),
.Y(n_249)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_249),
.Y(n_315)
);

BUFx12f_ASAP7_75t_L g251 ( 
.A(n_141),
.Y(n_251)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_251),
.Y(n_325)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_137),
.Y(n_252)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_252),
.Y(n_334)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_170),
.Y(n_254)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_254),
.Y(n_301)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_184),
.Y(n_255)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_255),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_188),
.B(n_44),
.Y(n_256)
);

AND2x4_ASAP7_75t_L g258 ( 
.A(n_162),
.B(n_50),
.Y(n_258)
);

AND2x2_ASAP7_75t_SL g288 ( 
.A(n_258),
.B(n_279),
.Y(n_288)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_149),
.Y(n_259)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_259),
.Y(n_318)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_182),
.Y(n_260)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_260),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_198),
.B(n_54),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_261),
.B(n_271),
.Y(n_307)
);

AND2x2_ASAP7_75t_SL g263 ( 
.A(n_199),
.B(n_57),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_185),
.Y(n_264)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_264),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_203),
.Y(n_265)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_265),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_206),
.B(n_57),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_266),
.B(n_269),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_136),
.A2(n_146),
.B1(n_148),
.B2(n_170),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_153),
.A2(n_88),
.B1(n_73),
.B2(n_68),
.Y(n_268)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_149),
.Y(n_270)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_270),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_203),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_154),
.A2(n_175),
.B1(n_187),
.B2(n_191),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_L g273 ( 
.A1(n_140),
.A2(n_50),
.B1(n_56),
.B2(n_6),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_273),
.A2(n_281),
.B1(n_168),
.B2(n_175),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_141),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_275),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_144),
.B(n_3),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_148),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_276),
.B(n_277),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_160),
.B(n_4),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_150),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_278),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_140),
.A2(n_56),
.B1(n_8),
.B2(n_9),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_154),
.A2(n_56),
.B1(n_10),
.B2(n_11),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_142),
.B(n_7),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_282),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_136),
.A2(n_56),
.B1(n_10),
.B2(n_12),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_283),
.A2(n_195),
.B1(n_168),
.B2(n_191),
.Y(n_320)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_173),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_284),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_218),
.B(n_196),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_285),
.B(n_289),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_218),
.B(n_172),
.C(n_176),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_290),
.B(n_317),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_247),
.A2(n_151),
.B1(n_179),
.B2(n_173),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_295),
.A2(n_316),
.B1(n_330),
.B2(n_222),
.Y(n_384)
);

OAI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_217),
.A2(n_158),
.B1(n_208),
.B2(n_195),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g380 ( 
.A1(n_296),
.A2(n_309),
.B1(n_313),
.B2(n_339),
.Y(n_380)
);

AOI32xp33_ASAP7_75t_L g308 ( 
.A1(n_230),
.A2(n_146),
.A3(n_201),
.B1(n_192),
.B2(n_163),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_SL g368 ( 
.A(n_308),
.B(n_238),
.C(n_209),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_217),
.A2(n_138),
.B1(n_171),
.B2(n_152),
.Y(n_309)
);

AO22x2_ASAP7_75t_SL g313 ( 
.A1(n_239),
.A2(n_147),
.B1(n_201),
.B2(n_192),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_220),
.A2(n_151),
.B1(n_179),
.B2(n_187),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_320),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_321),
.Y(n_376)
);

AND2x2_ASAP7_75t_SL g327 ( 
.A(n_263),
.B(n_130),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_327),
.B(n_264),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_263),
.A2(n_138),
.B1(n_131),
.B2(n_193),
.Y(n_330)
);

OAI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_262),
.A2(n_161),
.B1(n_155),
.B2(n_159),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_268),
.A2(n_209),
.B1(n_190),
.B2(n_12),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_341),
.A2(n_240),
.B1(n_249),
.B2(n_242),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_307),
.B(n_279),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_342),
.B(n_343),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_327),
.B(n_227),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_327),
.B(n_258),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_344),
.B(n_355),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_324),
.B(n_257),
.Y(n_345)
);

NAND3xp33_ASAP7_75t_L g395 ( 
.A(n_345),
.B(n_350),
.C(n_354),
.Y(n_395)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_322),
.Y(n_346)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_346),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_338),
.B(n_304),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_347),
.B(n_348),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_336),
.B(n_253),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_323),
.Y(n_349)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_349),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_298),
.B(n_250),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_292),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_351),
.B(n_352),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_340),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_306),
.Y(n_353)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_353),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_287),
.B(n_220),
.Y(n_354)
);

AND2x6_ASAP7_75t_L g355 ( 
.A(n_313),
.B(n_258),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_288),
.B(n_212),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_356),
.B(n_357),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_288),
.B(n_221),
.Y(n_357)
);

INVx4_ASAP7_75t_SL g358 ( 
.A(n_313),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_358),
.Y(n_387)
);

INVx13_ASAP7_75t_L g360 ( 
.A(n_319),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_360),
.Y(n_390)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_329),
.Y(n_361)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_361),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_362),
.B(n_364),
.Y(n_414)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_306),
.Y(n_363)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_363),
.Y(n_418)
);

INVx2_ASAP7_75t_SL g364 ( 
.A(n_326),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_334),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_365),
.B(n_367),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_288),
.B(n_236),
.Y(n_367)
);

OR2x4_ASAP7_75t_L g421 ( 
.A(n_368),
.B(n_325),
.Y(n_421)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_329),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_369),
.B(n_370),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_291),
.B(n_260),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_289),
.B(n_259),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_371),
.B(n_385),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_302),
.B(n_235),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_372),
.B(n_374),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_300),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_305),
.A2(n_233),
.B(n_270),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_375),
.A2(n_377),
.B(n_378),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_285),
.B(n_254),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_290),
.B(n_235),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_379),
.A2(n_381),
.B1(n_314),
.B2(n_311),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_314),
.A2(n_276),
.B1(n_224),
.B2(n_234),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_334),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_382),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_319),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_383),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_384),
.A2(n_286),
.B1(n_341),
.B2(n_333),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_309),
.B(n_284),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_376),
.A2(n_293),
.B1(n_317),
.B2(n_321),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_389),
.A2(n_394),
.B1(n_398),
.B2(n_404),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_391),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_373),
.A2(n_293),
.B1(n_305),
.B2(n_330),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_396),
.A2(n_358),
.B1(n_355),
.B2(n_375),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_376),
.A2(n_380),
.B1(n_342),
.B2(n_357),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_359),
.B(n_318),
.C(n_301),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_400),
.B(n_403),
.C(n_405),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_359),
.B(n_371),
.C(n_356),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_376),
.A2(n_231),
.B1(n_310),
.B2(n_248),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_359),
.B(n_332),
.C(n_337),
.Y(n_405)
);

MAJx2_ASAP7_75t_L g409 ( 
.A(n_367),
.B(n_311),
.C(n_325),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_409),
.B(n_417),
.C(n_382),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_343),
.A2(n_366),
.B1(n_385),
.B2(n_344),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_L g427 ( 
.A1(n_412),
.A2(n_358),
.B1(n_355),
.B2(n_377),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_366),
.A2(n_335),
.B1(n_315),
.B2(n_310),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_413),
.A2(n_420),
.B1(n_364),
.B2(n_361),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_366),
.B(n_337),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_384),
.A2(n_335),
.B1(n_315),
.B2(n_331),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_421),
.A2(n_372),
.B(n_346),
.Y(n_439)
);

OAI32xp33_ASAP7_75t_L g422 ( 
.A1(n_362),
.A2(n_299),
.A3(n_252),
.B1(n_297),
.B2(n_328),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_422),
.B(n_370),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_414),
.B(n_352),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_423),
.B(n_431),
.Y(n_460)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_386),
.Y(n_424)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_424),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_403),
.B(n_378),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_425),
.B(n_449),
.C(n_405),
.Y(n_461)
);

AOI22xp33_ASAP7_75t_SL g477 ( 
.A1(n_426),
.A2(n_404),
.B1(n_416),
.B2(n_422),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_427),
.Y(n_485)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_386),
.Y(n_428)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_428),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_395),
.B(n_348),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_429),
.B(n_433),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_392),
.B(n_347),
.Y(n_430)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_430),
.B(n_439),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_414),
.B(n_351),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_432),
.A2(n_434),
.B1(n_456),
.B2(n_410),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_407),
.B(n_350),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_396),
.A2(n_368),
.B1(n_345),
.B2(n_354),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_435),
.B(n_420),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_397),
.B(n_383),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_436),
.B(n_440),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_387),
.B(n_374),
.Y(n_437)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_437),
.Y(n_462)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_393),
.Y(n_438)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_438),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_408),
.B(n_349),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_415),
.B(n_361),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_441),
.A2(n_445),
.B(n_413),
.Y(n_464)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_393),
.Y(n_442)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_442),
.Y(n_475)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_418),
.Y(n_443)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_443),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_387),
.B(n_364),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_444),
.B(n_448),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_402),
.A2(n_369),
.B(n_297),
.Y(n_445)
);

INVx13_ASAP7_75t_L g446 ( 
.A(n_390),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_446),
.Y(n_478)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_418),
.Y(n_448)
);

INVx13_ASAP7_75t_L g451 ( 
.A(n_390),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_451),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_452),
.B(n_400),
.Y(n_458)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_401),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_453),
.B(n_454),
.Y(n_486)
);

NOR2x1_ASAP7_75t_R g454 ( 
.A(n_417),
.B(n_365),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_388),
.B(n_363),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_455),
.B(n_388),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_402),
.A2(n_331),
.B1(n_303),
.B2(n_271),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_458),
.B(n_461),
.C(n_463),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_425),
.B(n_399),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_464),
.B(n_471),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_445),
.A2(n_415),
.B(n_399),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_465),
.B(n_466),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_447),
.A2(n_398),
.B1(n_389),
.B2(n_412),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_470),
.A2(n_477),
.B1(n_450),
.B2(n_436),
.Y(n_490)
);

A2O1A1Ixp33_ASAP7_75t_L g471 ( 
.A1(n_439),
.A2(n_410),
.B(n_419),
.C(n_421),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_472),
.A2(n_431),
.B1(n_437),
.B2(n_444),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_435),
.A2(n_419),
.B(n_411),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_473),
.B(n_484),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_449),
.B(n_409),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_474),
.B(n_476),
.C(n_480),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_452),
.B(n_411),
.C(n_416),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_455),
.B(n_312),
.C(n_353),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_441),
.B(n_312),
.C(n_294),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_482),
.B(n_443),
.C(n_442),
.Y(n_505)
);

CKINVDCx14_ASAP7_75t_R g504 ( 
.A(n_483),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_453),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_490),
.A2(n_497),
.B1(n_506),
.B2(n_510),
.Y(n_525)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_469),
.Y(n_491)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_491),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_488),
.A2(n_429),
.B1(n_433),
.B2(n_450),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_493),
.Y(n_518)
);

NOR2x1_ASAP7_75t_L g494 ( 
.A(n_479),
.B(n_441),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_494),
.B(n_500),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_458),
.B(n_423),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_495),
.B(n_505),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_483),
.A2(n_432),
.B1(n_456),
.B2(n_434),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_498),
.A2(n_501),
.B1(n_515),
.B2(n_473),
.Y(n_524)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_467),
.Y(n_499)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_499),
.Y(n_522)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_467),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_485),
.A2(n_441),
.B1(n_426),
.B2(n_454),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_488),
.A2(n_430),
.B1(n_440),
.B2(n_448),
.Y(n_503)
);

CKINVDCx14_ASAP7_75t_R g519 ( 
.A(n_503),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_472),
.A2(n_454),
.B1(n_428),
.B2(n_438),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_469),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_508),
.B(n_511),
.Y(n_537)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_460),
.Y(n_509)
);

INVx1_ASAP7_75t_SL g539 ( 
.A(n_509),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_470),
.A2(n_424),
.B1(n_446),
.B2(n_451),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_457),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_461),
.B(n_406),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_512),
.B(n_514),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_476),
.B(n_406),
.C(n_294),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_513),
.B(n_487),
.C(n_478),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_474),
.B(n_451),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_483),
.A2(n_446),
.B1(n_303),
.B2(n_265),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_457),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_516),
.B(n_481),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_463),
.B(n_244),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_517),
.B(n_480),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_494),
.A2(n_465),
.B(n_464),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g543 ( 
.A1(n_523),
.A2(n_504),
.B(n_510),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_524),
.A2(n_541),
.B1(n_459),
.B2(n_328),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_526),
.B(n_535),
.C(n_496),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_497),
.B(n_460),
.Y(n_527)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_527),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_528),
.B(n_489),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_507),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_529),
.B(n_530),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_512),
.B(n_482),
.C(n_485),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_506),
.A2(n_462),
.B1(n_486),
.B2(n_484),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_531),
.A2(n_492),
.B1(n_505),
.B2(n_502),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_492),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_532),
.B(n_468),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_496),
.B(n_486),
.C(n_462),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_515),
.B(n_481),
.Y(n_536)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_536),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_495),
.B(n_471),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_SL g547 ( 
.A(n_538),
.B(n_517),
.Y(n_547)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_540),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_498),
.A2(n_501),
.B1(n_491),
.B2(n_509),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_542),
.A2(n_556),
.B1(n_541),
.B2(n_536),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_543),
.A2(n_536),
.B(n_526),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_521),
.B(n_514),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_545),
.B(n_547),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_546),
.B(n_553),
.Y(n_561)
);

XNOR2x1_ASAP7_75t_L g548 ( 
.A(n_524),
.B(n_513),
.Y(n_548)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_548),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_527),
.B(n_475),
.Y(n_549)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_549),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_551),
.B(n_553),
.C(n_546),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_521),
.B(n_489),
.C(n_475),
.Y(n_553)
);

CKINVDCx14_ASAP7_75t_R g555 ( 
.A(n_537),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_555),
.B(n_559),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_518),
.A2(n_468),
.B1(n_459),
.B2(n_215),
.Y(n_556)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_557),
.Y(n_572)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_533),
.Y(n_558)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_558),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_539),
.B(n_522),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_560),
.A2(n_525),
.B1(n_531),
.B2(n_539),
.Y(n_562)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_562),
.Y(n_578)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_563),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_542),
.A2(n_518),
.B1(n_519),
.B2(n_530),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_564),
.B(n_567),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_560),
.A2(n_525),
.B1(n_544),
.B2(n_534),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_568),
.B(n_360),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_552),
.B(n_535),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_569),
.B(n_570),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_551),
.B(n_520),
.C(n_528),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_SL g573 ( 
.A1(n_554),
.A2(n_523),
.B(n_559),
.Y(n_573)
);

MAJx2_ASAP7_75t_L g583 ( 
.A(n_573),
.B(n_543),
.C(n_549),
.Y(n_583)
);

OAI21xp33_ASAP7_75t_SL g590 ( 
.A1(n_574),
.A2(n_240),
.B(n_223),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_550),
.B(n_522),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_577),
.B(n_299),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_568),
.B(n_548),
.C(n_545),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_580),
.B(n_582),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_561),
.B(n_556),
.Y(n_581)
);

NAND3xp33_ASAP7_75t_L g594 ( 
.A(n_581),
.B(n_589),
.C(n_572),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_570),
.B(n_520),
.C(n_554),
.Y(n_582)
);

AOI31xp67_ASAP7_75t_L g597 ( 
.A1(n_583),
.A2(n_562),
.A3(n_567),
.B(n_576),
.Y(n_597)
);

NOR2x1_ASAP7_75t_L g585 ( 
.A(n_566),
.B(n_538),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g593 ( 
.A1(n_585),
.A2(n_574),
.B(n_565),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_564),
.B(n_547),
.C(n_360),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_586),
.B(n_576),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_588),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g600 ( 
.A(n_590),
.B(n_578),
.Y(n_600)
);

MAJx2_ASAP7_75t_L g591 ( 
.A(n_587),
.B(n_573),
.C(n_571),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g604 ( 
.A(n_591),
.B(n_597),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_SL g592 ( 
.A(n_582),
.B(n_575),
.Y(n_592)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_592),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_593),
.B(n_594),
.Y(n_605)
);

NAND4xp25_ASAP7_75t_L g595 ( 
.A(n_579),
.B(n_565),
.C(n_571),
.D(n_563),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_595),
.A2(n_600),
.B1(n_590),
.B2(n_584),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_598),
.B(n_599),
.Y(n_601)
);

NOR3xp33_ASAP7_75t_L g609 ( 
.A(n_601),
.B(n_190),
.C(n_219),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_602),
.A2(n_606),
.B(n_225),
.Y(n_608)
);

AOI322xp5_ASAP7_75t_L g603 ( 
.A1(n_596),
.A2(n_583),
.A3(n_585),
.B1(n_228),
.B2(n_251),
.C1(n_274),
.C2(n_213),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_603),
.B(n_7),
.C(n_12),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_598),
.B(n_251),
.Y(n_606)
);

AOI322xp5_ASAP7_75t_L g612 ( 
.A1(n_608),
.A2(n_609),
.A3(n_610),
.B1(n_611),
.B2(n_607),
.C1(n_603),
.C2(n_14),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_605),
.A2(n_213),
.B(n_10),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_612),
.Y(n_614)
);

AOI322xp5_ASAP7_75t_L g613 ( 
.A1(n_608),
.A2(n_604),
.A3(n_13),
.B1(n_15),
.B2(n_16),
.C1(n_17),
.C2(n_18),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_614),
.B(n_613),
.C(n_13),
.Y(n_615)
);

OAI21xp5_ASAP7_75t_SL g616 ( 
.A1(n_615),
.A2(n_7),
.B(n_15),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_L g617 ( 
.A(n_616),
.B(n_7),
.Y(n_617)
);

XOR2xp5_ASAP7_75t_L g618 ( 
.A(n_617),
.B(n_16),
.Y(n_618)
);


endmodule