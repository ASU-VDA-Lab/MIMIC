module fake_jpeg_984_n_512 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_512);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_512;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx4f_ASAP7_75t_SL g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_3),
.B(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_6),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_14),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_32),
.B(n_15),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_59),
.B(n_82),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_2),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_60),
.B(n_63),
.Y(n_134)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_61),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_3),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_64),
.Y(n_147)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_65),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_67),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_68),
.Y(n_172)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_69),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_70),
.Y(n_154)
);

INVx6_ASAP7_75t_SL g71 ( 
.A(n_50),
.Y(n_71)
);

INVx6_ASAP7_75t_SL g132 ( 
.A(n_71),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_72),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_4),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_73),
.B(n_85),
.Y(n_139)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_75),
.Y(n_171)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_77),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_79),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_80),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_81),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_18),
.B(n_6),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_83),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_16),
.B(n_14),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_84),
.B(n_95),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_16),
.B(n_7),
.Y(n_85)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_86),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_87),
.Y(n_165)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_89),
.Y(n_136)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_21),
.Y(n_90)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_90),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_19),
.Y(n_93)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_93),
.Y(n_140)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_94),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_19),
.B(n_8),
.Y(n_95)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_22),
.B(n_8),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_97),
.B(n_99),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_17),
.B(n_14),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_100),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_17),
.B(n_41),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_101),
.B(n_112),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_102),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_22),
.B(n_9),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_103),
.B(n_111),
.Y(n_183)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_104),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_105),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_109),
.Y(n_167)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_110),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_27),
.B(n_11),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_56),
.B(n_11),
.Y(n_112)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_40),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_117),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_20),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_118),
.Y(n_148)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_31),
.Y(n_115)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_115),
.Y(n_186)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_40),
.Y(n_116)
);

AOI21xp33_ASAP7_75t_L g161 ( 
.A1(n_116),
.A2(n_35),
.B(n_29),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_20),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_23),
.B(n_11),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_40),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_120),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_20),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_27),
.B(n_12),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_121),
.B(n_36),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_98),
.A2(n_24),
.B1(n_41),
.B2(n_51),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_124),
.A2(n_187),
.B1(n_171),
.B2(n_177),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_102),
.A2(n_33),
.B1(n_51),
.B2(n_44),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_126),
.A2(n_141),
.B1(n_169),
.B2(n_185),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_112),
.A2(n_53),
.B1(n_39),
.B2(n_30),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_135),
.A2(n_150),
.B1(n_92),
.B2(n_88),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_117),
.A2(n_24),
.B1(n_39),
.B2(n_30),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_60),
.B(n_53),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_143),
.B(n_153),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_63),
.A2(n_29),
.B1(n_28),
.B2(n_55),
.Y(n_150)
);

CKINVDCx12_ASAP7_75t_R g152 ( 
.A(n_67),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_152),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_73),
.B(n_33),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_55),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_155),
.B(n_168),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_161),
.B(n_135),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_69),
.B(n_87),
.C(n_106),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_163),
.B(n_128),
.C(n_172),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_100),
.B(n_44),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_72),
.A2(n_28),
.B1(n_36),
.B2(n_23),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_173),
.B(n_174),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_100),
.B(n_35),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_109),
.B(n_35),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_176),
.B(n_188),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_65),
.A2(n_42),
.B1(n_13),
.B2(n_14),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_62),
.A2(n_75),
.B1(n_81),
.B2(n_80),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_66),
.B(n_12),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_68),
.B(n_83),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_189),
.B(n_190),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_86),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_72),
.A2(n_13),
.B1(n_42),
.B2(n_78),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_192),
.A2(n_169),
.B1(n_141),
.B2(n_150),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_77),
.B(n_94),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_193),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_90),
.B(n_113),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_195),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_123),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_197),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_198),
.B(n_199),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_132),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_127),
.Y(n_200)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_200),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_105),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_201),
.Y(n_273)
);

INVx11_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_202),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_123),
.Y(n_203)
);

INVx8_ASAP7_75t_L g296 ( 
.A(n_203),
.Y(n_296)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_157),
.Y(n_205)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_205),
.Y(n_307)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_144),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_206),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_148),
.A2(n_116),
.B1(n_108),
.B2(n_91),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_207),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_132),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_208),
.B(n_209),
.Y(n_271)
);

A2O1A1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_134),
.A2(n_96),
.B(n_89),
.C(n_70),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_210),
.Y(n_275)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_127),
.Y(n_211)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_211),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_213),
.A2(n_237),
.B1(n_250),
.B2(n_255),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_215),
.A2(n_226),
.B1(n_233),
.B2(n_239),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_164),
.B(n_159),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_216),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_154),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_217),
.Y(n_283)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_165),
.Y(n_219)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_219),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_184),
.Y(n_220)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_220),
.Y(n_280)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_165),
.Y(n_221)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_221),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_149),
.Y(n_222)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_222),
.Y(n_284)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_138),
.Y(n_223)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_223),
.Y(n_301)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_140),
.Y(n_224)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_224),
.Y(n_302)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_151),
.Y(n_225)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_225),
.Y(n_311)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_151),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_228),
.Y(n_263)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_L g229 ( 
.A1(n_146),
.A2(n_162),
.B(n_180),
.C(n_139),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_229),
.B(n_251),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_183),
.A2(n_124),
.B1(n_187),
.B2(n_131),
.Y(n_231)
);

OA21x2_ASAP7_75t_L g304 ( 
.A1(n_231),
.A2(n_232),
.B(n_225),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_159),
.A2(n_142),
.B1(n_184),
.B2(n_125),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_145),
.B(n_186),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_243),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_154),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_236),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_147),
.A2(n_191),
.B1(n_158),
.B2(n_125),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_142),
.Y(n_239)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_157),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_241),
.B(n_242),
.Y(n_292)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_182),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_163),
.B(n_182),
.Y(n_243)
);

NAND3xp33_ASAP7_75t_SL g244 ( 
.A(n_129),
.B(n_170),
.C(n_175),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_244),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_196),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_245),
.B(n_248),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_171),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_246),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_L g247 ( 
.A1(n_192),
.A2(n_160),
.B1(n_133),
.B2(n_122),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_247),
.A2(n_249),
.B1(n_239),
.B2(n_209),
.Y(n_286)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_175),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_177),
.A2(n_178),
.B1(n_129),
.B2(n_170),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_178),
.A2(n_181),
.B1(n_128),
.B2(n_172),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_130),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_122),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_252),
.B(n_254),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_156),
.C(n_137),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_130),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_181),
.A2(n_149),
.B1(n_194),
.B2(n_166),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_133),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_260),
.Y(n_268)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_136),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_257),
.B(n_222),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_194),
.A2(n_166),
.B1(n_136),
.B2(n_196),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_SL g288 ( 
.A(n_258),
.B(n_216),
.C(n_201),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_137),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_160),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_156),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_266),
.B(n_281),
.C(n_289),
.Y(n_347)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_269),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_243),
.B(n_253),
.C(n_232),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_286),
.A2(n_278),
.B1(n_279),
.B2(n_274),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g349 ( 
.A(n_288),
.B(n_304),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_218),
.B(n_235),
.C(n_234),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_218),
.B(n_235),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_290),
.B(n_293),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_231),
.A2(n_213),
.B1(n_212),
.B2(n_240),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_291),
.A2(n_298),
.B1(n_310),
.B2(n_308),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_230),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_200),
.B(n_211),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_294),
.B(n_295),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_238),
.B(n_216),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_247),
.A2(n_261),
.B1(n_201),
.B2(n_256),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_303),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_214),
.B(n_229),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_206),
.B(n_221),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_309),
.B(n_263),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_227),
.A2(n_242),
.B1(n_252),
.B2(n_203),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_210),
.A2(n_241),
.B1(n_219),
.B2(n_205),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_312),
.A2(n_197),
.B1(n_236),
.B2(n_246),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_313),
.B(n_315),
.Y(n_372)
);

AND2x2_ASAP7_75t_SL g315 ( 
.A(n_281),
.B(n_220),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_204),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_317),
.B(n_339),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_264),
.A2(n_217),
.B1(n_245),
.B2(n_226),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_318),
.A2(n_321),
.B1(n_324),
.B2(n_326),
.Y(n_353)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_311),
.Y(n_319)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_319),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_264),
.B(n_202),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_320),
.B(n_330),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_286),
.A2(n_271),
.B1(n_304),
.B2(n_287),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_296),
.Y(n_322)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_322),
.Y(n_357)
);

OA21x2_ASAP7_75t_L g323 ( 
.A1(n_291),
.A2(n_298),
.B(n_267),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_323),
.B(n_329),
.Y(n_361)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_294),
.Y(n_325)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_325),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_304),
.A2(n_274),
.B1(n_278),
.B2(n_290),
.Y(n_326)
);

INVx11_ASAP7_75t_L g327 ( 
.A(n_272),
.Y(n_327)
);

CKINVDCx10_ASAP7_75t_R g367 ( 
.A(n_327),
.Y(n_367)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_309),
.Y(n_328)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_328),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_289),
.B(n_295),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_270),
.Y(n_331)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_331),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_266),
.A2(n_273),
.B1(n_279),
.B2(n_285),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_332),
.A2(n_338),
.B1(n_341),
.B2(n_346),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_333),
.B(n_343),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_288),
.A2(n_268),
.B(n_300),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_334),
.A2(n_280),
.B(n_307),
.Y(n_364)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_311),
.Y(n_335)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_335),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_301),
.B(n_302),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_337),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_265),
.A2(n_297),
.B1(n_268),
.B2(n_284),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_301),
.B(n_302),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_270),
.B(n_276),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_340),
.B(n_345),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_310),
.A2(n_269),
.B1(n_305),
.B2(n_292),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_265),
.A2(n_297),
.B1(n_284),
.B2(n_283),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_342),
.Y(n_378)
);

CKINVDCx14_ASAP7_75t_R g344 ( 
.A(n_312),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_344),
.B(n_348),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_280),
.B(n_262),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_276),
.A2(n_275),
.B1(n_282),
.B2(n_277),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_283),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_275),
.Y(n_350)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_350),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_339),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_355),
.B(n_374),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_349),
.A2(n_277),
.B(n_282),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_359),
.A2(n_364),
.B(n_342),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_333),
.B(n_307),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_369),
.B(n_370),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_316),
.B(n_296),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_331),
.Y(n_371)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_371),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_340),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_346),
.Y(n_375)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_375),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_316),
.B(n_272),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_376),
.B(n_377),
.Y(n_390)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_350),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_341),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_379),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_349),
.A2(n_306),
.B(n_326),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_380),
.A2(n_320),
.B(n_332),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_381),
.B(n_382),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_317),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_380),
.A2(n_349),
.B(n_334),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_385),
.A2(n_386),
.B(n_401),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_353),
.A2(n_324),
.B1(n_336),
.B2(n_325),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_387),
.A2(n_391),
.B1(n_402),
.B2(n_405),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_356),
.B(n_347),
.C(n_315),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_388),
.B(n_389),
.C(n_393),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_356),
.B(n_347),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_353),
.A2(n_321),
.B1(n_323),
.B2(n_336),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_359),
.B(n_315),
.C(n_330),
.Y(n_393)
);

OA21x2_ASAP7_75t_L g394 ( 
.A1(n_361),
.A2(n_323),
.B(n_318),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_394),
.B(n_404),
.Y(n_420)
);

XOR2x1_ASAP7_75t_L g395 ( 
.A(n_361),
.B(n_323),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_395),
.B(n_372),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_355),
.B(n_328),
.Y(n_397)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_397),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_374),
.B(n_381),
.Y(n_398)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_398),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_351),
.B(n_315),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_399),
.B(n_352),
.C(n_360),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_352),
.A2(n_343),
.B1(n_314),
.B2(n_313),
.Y(n_402)
);

OA22x2_ASAP7_75t_L g404 ( 
.A1(n_375),
.A2(n_319),
.B1(n_335),
.B2(n_322),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_372),
.A2(n_314),
.B1(n_348),
.B2(n_306),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_368),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_406),
.B(n_407),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_368),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_370),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_408),
.B(n_371),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_409),
.Y(n_441)
);

OAI21xp33_ASAP7_75t_L g410 ( 
.A1(n_398),
.A2(n_364),
.B(n_382),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_410),
.B(n_416),
.Y(n_445)
);

AND2x6_ASAP7_75t_L g413 ( 
.A(n_406),
.B(n_372),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_413),
.A2(n_431),
.B1(n_408),
.B2(n_402),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_407),
.B(n_354),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_392),
.B(n_354),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_417),
.B(n_429),
.Y(n_446)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_390),
.Y(n_418)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_418),
.Y(n_450)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_390),
.Y(n_419)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_419),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_421),
.B(n_389),
.Y(n_439)
);

A2O1A1O1Ixp25_ASAP7_75t_L g424 ( 
.A1(n_393),
.A2(n_351),
.B(n_360),
.C(n_358),
.D(n_369),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_424),
.A2(n_427),
.B(n_428),
.Y(n_440)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_396),
.Y(n_425)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_425),
.Y(n_433)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_396),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_426),
.B(n_430),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_385),
.A2(n_378),
.B(n_376),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_386),
.A2(n_401),
.B(n_400),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_392),
.B(n_373),
.Y(n_429)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_397),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_411),
.B(n_388),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_SL g467 ( 
.A(n_434),
.B(n_435),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_411),
.B(n_388),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_422),
.A2(n_387),
.B1(n_391),
.B2(n_394),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_436),
.A2(n_438),
.B1(n_444),
.B2(n_449),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_439),
.B(n_443),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_421),
.B(n_389),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_442),
.B(n_399),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_427),
.B(n_393),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_414),
.A2(n_400),
.B1(n_394),
.B2(n_384),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_415),
.B(n_399),
.C(n_401),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_447),
.B(n_409),
.C(n_405),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_422),
.A2(n_403),
.B1(n_384),
.B2(n_395),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_448),
.A2(n_420),
.B1(n_424),
.B2(n_413),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_414),
.A2(n_394),
.B1(n_403),
.B2(n_358),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_428),
.A2(n_383),
.B(n_395),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_451),
.B(n_423),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_440),
.B(n_415),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_452),
.B(n_453),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_446),
.B(n_383),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_454),
.B(n_459),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_439),
.B(n_423),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_456),
.B(n_458),
.C(n_441),
.Y(n_473)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_457),
.B(n_443),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_450),
.B(n_430),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_436),
.A2(n_420),
.B1(n_431),
.B2(n_412),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_460),
.A2(n_461),
.B1(n_432),
.B2(n_437),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_445),
.A2(n_412),
.B1(n_419),
.B2(n_418),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_433),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_462),
.B(n_466),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_434),
.B(n_426),
.C(n_404),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_463),
.B(n_447),
.C(n_451),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_464),
.A2(n_432),
.B1(n_437),
.B2(n_433),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_442),
.B(n_404),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_468),
.A2(n_474),
.B1(n_453),
.B2(n_425),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_470),
.B(n_471),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_455),
.B(n_435),
.C(n_440),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_455),
.B(n_441),
.C(n_448),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_472),
.B(n_473),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_464),
.Y(n_476)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_476),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_477),
.A2(n_363),
.B1(n_377),
.B2(n_366),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_460),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_478),
.B(n_404),
.Y(n_487)
);

OAI21x1_ASAP7_75t_L g481 ( 
.A1(n_475),
.A2(n_456),
.B(n_467),
.Y(n_481)
);

NAND3xp33_ASAP7_75t_L g492 ( 
.A(n_481),
.B(n_471),
.C(n_470),
.Y(n_492)
);

INVx11_ASAP7_75t_L g482 ( 
.A(n_479),
.Y(n_482)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_482),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_476),
.A2(n_465),
.B(n_463),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_483),
.A2(n_484),
.B(n_487),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_468),
.A2(n_466),
.B(n_458),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_486),
.B(n_488),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_489),
.B(n_469),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_491),
.B(n_493),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_492),
.A2(n_496),
.B(n_480),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_484),
.B(n_472),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_489),
.B(n_357),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_495),
.A2(n_488),
.B1(n_363),
.B2(n_366),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_485),
.B(n_357),
.Y(n_496)
);

NOR3xp33_ASAP7_75t_L g504 ( 
.A(n_498),
.B(n_501),
.C(n_497),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_499),
.B(n_500),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_491),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_494),
.A2(n_483),
.B(n_467),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_490),
.B(n_482),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_503),
.B(n_404),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_504),
.B(n_505),
.Y(n_509)
);

OA21x2_ASAP7_75t_SL g505 ( 
.A1(n_500),
.A2(n_365),
.B(n_362),
.Y(n_505)
);

OAI311xp33_ASAP7_75t_L g508 ( 
.A1(n_506),
.A2(n_502),
.A3(n_367),
.B1(n_365),
.C1(n_362),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_508),
.B(n_507),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_510),
.B(n_509),
.C(n_367),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_511),
.B(n_327),
.Y(n_512)
);


endmodule