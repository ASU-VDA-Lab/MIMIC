module real_jpeg_29811_n_7 (n_5, n_4, n_0, n_1, n_2, n_6, n_3, n_7);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_3;

output n_7;

wire n_17;
wire n_8;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_57;
wire n_73;
wire n_65;
wire n_33;
wire n_35;
wire n_50;
wire n_38;
wire n_29;
wire n_55;
wire n_69;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_58;
wire n_67;
wire n_63;
wire n_12;
wire n_68;
wire n_76;
wire n_24;
wire n_75;
wire n_66;
wire n_34;
wire n_72;
wire n_44;
wire n_28;
wire n_60;
wire n_46;
wire n_62;
wire n_59;
wire n_64;
wire n_23;
wire n_11;
wire n_14;
wire n_51;
wire n_71;
wire n_47;
wire n_25;
wire n_61;
wire n_45;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_36;
wire n_40;
wire n_39;
wire n_70;
wire n_41;
wire n_26;
wire n_32;
wire n_56;
wire n_19;
wire n_20;
wire n_27;
wire n_30;
wire n_48;
wire n_74;
wire n_16;
wire n_15;
wire n_13;

INVx11_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

AOI21xp33_ASAP7_75t_L g14 ( 
.A1(n_2),
.A2(n_3),
.B(n_15),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_2),
.A2(n_12),
.B1(n_17),
.B2(n_26),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_2),
.A2(n_12),
.B1(n_15),
.B2(n_22),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_2),
.A2(n_5),
.B(n_62),
.C(n_63),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_2),
.A2(n_12),
.B1(n_63),
.B2(n_64),
.Y(n_72)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_3),
.A2(n_13),
.B1(n_15),
.B2(n_22),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx11_ASAP7_75t_SL g16 ( 
.A(n_6),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_56),
.Y(n_7)
);

OAI21xp5_ASAP7_75t_SL g8 ( 
.A1(n_9),
.A2(n_44),
.B(n_55),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_28),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_10),
.B(n_28),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_18),
.Y(n_10)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_11),
.A2(n_18),
.B1(n_19),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_13),
.B(n_14),
.C(n_17),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_12),
.B(n_21),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_12),
.B(n_51),
.Y(n_50)
);

OAI21xp33_ASAP7_75t_L g62 ( 
.A1(n_12),
.A2(n_26),
.B(n_36),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_13),
.A2(n_17),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_15),
.B(n_40),
.Y(n_41)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_17),
.A2(n_26),
.B1(n_34),
.B2(n_36),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_18),
.A2(n_19),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_18),
.A2(n_19),
.B1(n_68),
.B2(n_73),
.Y(n_67)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_19),
.B(n_30),
.C(n_43),
.Y(n_58)
);

AND2x2_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_27),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_23),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_22),
.B(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_37),
.B1(n_42),
.B2(n_43),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_33),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_33),
.B(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_34),
.A2(n_36),
.B1(n_63),
.B2(n_64),
.Y(n_71)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_43),
.B1(n_61),
.B2(n_65),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_43),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_43),
.B(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_52),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_48),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_75),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_59),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_66),
.B1(n_67),
.B2(n_74),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_68),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);


endmodule