module fake_jpeg_2404_n_537 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_537);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_537;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_12),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_48),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_52),
.B(n_53),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_48),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_54),
.Y(n_135)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_55),
.Y(n_153)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_56),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_57),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_59),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_60),
.B(n_62),
.Y(n_109)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_61),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_73),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_30),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_66),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_35),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_35),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_67),
.B(n_70),
.Y(n_112)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_50),
.Y(n_68)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_71),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_39),
.B(n_9),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_80),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_77),
.Y(n_124)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_78),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_25),
.B(n_0),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_81),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_82),
.Y(n_148)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_50),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_86),
.B(n_92),
.Y(n_125)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_19),
.B(n_26),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_88),
.B(n_32),
.Y(n_139)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_35),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_49),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_94),
.B(n_95),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_39),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_96),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_42),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_97),
.B(n_99),
.Y(n_149)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g136 ( 
.A(n_98),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_42),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_100),
.Y(n_132)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

INVx3_ASAP7_75t_SL g142 ( 
.A(n_101),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_28),
.B(n_1),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_1),
.Y(n_130)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_106),
.Y(n_165)
);

NOR2x1_ASAP7_75t_R g108 ( 
.A(n_51),
.B(n_23),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_108),
.B(n_133),
.Y(n_205)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_111),
.Y(n_180)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_118),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_62),
.A2(n_49),
.B1(n_32),
.B2(n_19),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_122),
.A2(n_123),
.B1(n_150),
.B2(n_155),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_55),
.A2(n_32),
.B1(n_69),
.B2(n_83),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_130),
.B(n_14),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_64),
.A2(n_23),
.B1(n_38),
.B2(n_37),
.Y(n_133)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_56),
.Y(n_138)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_88),
.Y(n_168)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_141),
.Y(n_198)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_147),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_73),
.A2(n_45),
.B1(n_47),
.B2(n_37),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_151),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_70),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_163),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_61),
.A2(n_19),
.B1(n_47),
.B2(n_45),
.Y(n_155)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_79),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_158),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_80),
.A2(n_31),
.B1(n_20),
.B2(n_29),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_159),
.A2(n_29),
.B1(n_31),
.B2(n_20),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_98),
.A2(n_19),
.B1(n_38),
.B2(n_44),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_160),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_102),
.B(n_33),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_164),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_149),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_167),
.B(n_176),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_168),
.B(n_144),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_112),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_170),
.B(n_181),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_103),
.B(n_88),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_171),
.B(n_177),
.C(n_196),
.Y(n_252)
);

O2A1O1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_159),
.A2(n_71),
.B(n_91),
.C(n_87),
.Y(n_172)
);

OA22x2_ASAP7_75t_L g246 ( 
.A1(n_172),
.A2(n_107),
.B1(n_126),
.B2(n_144),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_173),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_105),
.B(n_120),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_174),
.B(n_184),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_129),
.A2(n_46),
.B1(n_101),
.B2(n_33),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_175),
.A2(n_183),
.B1(n_187),
.B2(n_216),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_109),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_85),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_178),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_179),
.A2(n_217),
.B1(n_223),
.B2(n_146),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_125),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_136),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_182),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_148),
.A2(n_46),
.B1(n_93),
.B2(n_57),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_57),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_110),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_186),
.B(n_200),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_148),
.A2(n_93),
.B1(n_54),
.B2(n_84),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_132),
.B(n_68),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_188),
.B(n_202),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_113),
.B(n_96),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_190),
.Y(n_242)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_114),
.Y(n_192)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_192),
.Y(n_236)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_115),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_193),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_122),
.A2(n_90),
.B1(n_81),
.B2(n_75),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_194),
.A2(n_214),
.B1(n_219),
.B2(n_156),
.Y(n_224)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_127),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_195),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_131),
.B(n_72),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_142),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_197),
.B(n_206),
.Y(n_270)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_143),
.Y(n_199)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_199),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_152),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_143),
.Y(n_201)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_201),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_134),
.B(n_2),
.Y(n_202)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_117),
.Y(n_203)
);

INVx3_ASAP7_75t_SL g265 ( 
.A(n_203),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_155),
.B(n_3),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_204),
.B(n_208),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_104),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_153),
.B(n_4),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_104),
.Y(n_209)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_209),
.Y(n_249)
);

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_119),
.Y(n_210)
);

INVx11_ASAP7_75t_L g275 ( 
.A(n_210),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_SL g211 ( 
.A(n_160),
.B(n_82),
.C(n_15),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_211),
.B(n_221),
.C(n_222),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_123),
.A2(n_59),
.B(n_89),
.Y(n_212)
);

NAND2xp33_ASAP7_75t_SL g253 ( 
.A(n_212),
.B(n_18),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_213),
.B(n_166),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_106),
.A2(n_89),
.B1(n_14),
.B2(n_8),
.Y(n_214)
);

NAND2x1_ASAP7_75t_SL g215 ( 
.A(n_142),
.B(n_5),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_215),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_117),
.A2(n_5),
.B1(n_9),
.B2(n_10),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_111),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_135),
.Y(n_220)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_220),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_118),
.B(n_10),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_158),
.B(n_15),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_157),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_224),
.A2(n_226),
.B1(n_191),
.B2(n_185),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_225),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_169),
.A2(n_156),
.B1(n_146),
.B2(n_128),
.Y(n_226)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_210),
.Y(n_227)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_227),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_232),
.A2(n_233),
.B1(n_245),
.B2(n_250),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_204),
.A2(n_124),
.B1(n_128),
.B2(n_121),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_203),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_237),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_168),
.B(n_145),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_239),
.Y(n_281)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_180),
.Y(n_240)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_240),
.Y(n_292)
);

AO22x1_ASAP7_75t_L g244 ( 
.A1(n_194),
.A2(n_119),
.B1(n_162),
.B2(n_126),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_244),
.A2(n_191),
.B(n_190),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_168),
.A2(n_124),
.B1(n_121),
.B2(n_162),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_246),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_170),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_247),
.B(n_256),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_205),
.A2(n_107),
.B1(n_144),
.B2(n_137),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_253),
.A2(n_211),
.B(n_190),
.Y(n_279)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_180),
.Y(n_255)
);

INVx3_ASAP7_75t_SL g285 ( 
.A(n_255),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_197),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_181),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_257),
.B(n_266),
.Y(n_316)
);

INVx13_ASAP7_75t_L g258 ( 
.A(n_209),
.Y(n_258)
);

INVx13_ASAP7_75t_L g301 ( 
.A(n_258),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_205),
.A2(n_16),
.B1(n_17),
.B2(n_212),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_259),
.A2(n_262),
.B1(n_267),
.B2(n_269),
.Y(n_320)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_164),
.Y(n_260)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_260),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_172),
.A2(n_16),
.B1(n_208),
.B2(n_202),
.Y(n_262)
);

AND2x2_ASAP7_75t_SL g264 ( 
.A(n_188),
.B(n_177),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_264),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_215),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_221),
.A2(n_222),
.B1(n_171),
.B2(n_178),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_165),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_268),
.B(n_274),
.Y(n_319)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_230),
.Y(n_277)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_277),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_196),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_278),
.B(n_299),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_279),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_253),
.A2(n_207),
.B(n_189),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_280),
.A2(n_287),
.B(n_321),
.Y(n_332)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_230),
.Y(n_282)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_282),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_192),
.C(n_207),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_284),
.B(n_290),
.C(n_307),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_286),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_229),
.A2(n_198),
.B(n_189),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_234),
.Y(n_288)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_288),
.Y(n_344)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_234),
.Y(n_289)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_289),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_252),
.B(n_264),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_291),
.A2(n_320),
.B1(n_268),
.B2(n_265),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_198),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_294),
.B(n_296),
.Y(n_330)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_260),
.Y(n_295)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_295),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_251),
.B(n_218),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_270),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_297),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_228),
.B(n_218),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_298),
.B(n_304),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_231),
.B(n_185),
.Y(n_299)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_236),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_302),
.Y(n_324)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_236),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_303),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_241),
.B(n_165),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_254),
.B(n_210),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_305),
.B(n_306),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_231),
.B(n_214),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_264),
.B(n_191),
.C(n_239),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_272),
.A2(n_224),
.B1(n_226),
.B2(n_242),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_309),
.A2(n_312),
.B1(n_245),
.B2(n_246),
.Y(n_342)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_243),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_313),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_272),
.A2(n_271),
.B1(n_262),
.B2(n_239),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_243),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_254),
.B(n_248),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_249),
.Y(n_329)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_248),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_317),
.Y(n_345)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_238),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_259),
.A2(n_269),
.B(n_225),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_238),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_323),
.B(n_238),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_329),
.B(n_331),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_297),
.B(n_261),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_322),
.A2(n_244),
.B1(n_233),
.B2(n_225),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_334),
.B(n_360),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_316),
.A2(n_250),
.B(n_244),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_336),
.A2(n_341),
.B(n_349),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_338),
.A2(n_342),
.B1(n_358),
.B2(n_361),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_308),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_340),
.B(n_350),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_279),
.A2(n_246),
.B(n_249),
.Y(n_341)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_346),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_290),
.B(n_273),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_347),
.B(n_354),
.C(n_355),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_283),
.A2(n_246),
.B1(n_227),
.B2(n_265),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_319),
.B(n_235),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_284),
.B(n_235),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_351),
.B(n_357),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_301),
.Y(n_352)
);

BUFx24_ASAP7_75t_L g382 ( 
.A(n_352),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_301),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_353),
.B(n_300),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_307),
.B(n_278),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_318),
.B(n_240),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_299),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_309),
.A2(n_237),
.B1(n_255),
.B2(n_258),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_322),
.A2(n_275),
.B1(n_312),
.B2(n_286),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_306),
.A2(n_275),
.B1(n_321),
.B2(n_281),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_276),
.B(n_277),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_362),
.B(n_364),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_276),
.B(n_295),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_310),
.B(n_313),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_365),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_326),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_366),
.B(n_372),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_356),
.A2(n_287),
.B(n_311),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_368),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_370),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_342),
.A2(n_281),
.B1(n_288),
.B2(n_282),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_371),
.A2(n_386),
.B1(n_387),
.B2(n_380),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_326),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_354),
.B(n_289),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_374),
.B(n_400),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_345),
.B(n_302),
.Y(n_377)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_377),
.Y(n_409)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_362),
.Y(n_378)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_378),
.Y(n_411)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_364),
.Y(n_380)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_380),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_328),
.B(n_315),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_381),
.B(n_347),
.C(n_361),
.Y(n_402)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_324),
.Y(n_384)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_384),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_325),
.A2(n_303),
.B1(n_323),
.B2(n_317),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_345),
.Y(n_387)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_387),
.Y(n_427)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_324),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_388),
.Y(n_424)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_324),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_389),
.B(n_392),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_356),
.A2(n_341),
.B(n_332),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_391),
.A2(n_332),
.B(n_339),
.Y(n_405)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_333),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_363),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_393),
.Y(n_410)
);

OAI32xp33_ASAP7_75t_L g394 ( 
.A1(n_325),
.A2(n_280),
.A3(n_292),
.B1(n_285),
.B2(n_300),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_394),
.B(n_396),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_360),
.A2(n_285),
.B1(n_293),
.B2(n_292),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_395),
.A2(n_349),
.B1(n_358),
.B2(n_336),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_363),
.B(n_285),
.Y(n_396)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_333),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_398),
.B(n_399),
.Y(n_415)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_337),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_328),
.B(n_293),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_346),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_401),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_402),
.B(n_421),
.C(n_426),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_403),
.A2(n_407),
.B1(n_418),
.B2(n_395),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_SL g443 ( 
.A(n_405),
.B(n_371),
.C(n_390),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_381),
.B(n_355),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_412),
.B(n_419),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_370),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_414),
.B(n_417),
.Y(n_447)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_370),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_367),
.A2(n_327),
.B1(n_343),
.B2(n_335),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_374),
.B(n_330),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_383),
.B(n_339),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_420),
.B(n_397),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_383),
.B(n_343),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_337),
.C(n_344),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_379),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_429),
.B(n_430),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_377),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_385),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_431),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_396),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_432),
.B(n_376),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_434),
.B(n_421),
.Y(n_468)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_415),
.Y(n_435)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_435),
.Y(n_459)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_415),
.Y(n_436)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_436),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_437),
.A2(n_451),
.B1(n_403),
.B2(n_424),
.Y(n_476)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_404),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_438),
.B(n_441),
.Y(n_465)
);

XOR2x2_ASAP7_75t_SL g440 ( 
.A(n_408),
.B(n_391),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_440),
.B(n_443),
.Y(n_460)
);

BUFx24_ASAP7_75t_SL g441 ( 
.A(n_423),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_442),
.Y(n_478)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_404),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_444),
.B(n_445),
.Y(n_470)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_422),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_410),
.B(n_376),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_446),
.B(n_452),
.Y(n_469)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_422),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_448),
.B(n_449),
.Y(n_462)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_428),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_408),
.A2(n_369),
.B1(n_373),
.B2(n_378),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_411),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_416),
.B(n_368),
.C(n_375),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_453),
.B(n_456),
.C(n_457),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_432),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_454),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_416),
.B(n_375),
.C(n_386),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_426),
.B(n_369),
.C(n_390),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_409),
.A2(n_427),
.B(n_413),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_458),
.A2(n_427),
.B(n_413),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g464 ( 
.A(n_455),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_464),
.B(n_472),
.Y(n_491)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_466),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_468),
.B(n_479),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_446),
.B(n_409),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_471),
.Y(n_485)
);

CKINVDCx14_ASAP7_75t_R g472 ( 
.A(n_447),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_442),
.A2(n_411),
.B(n_406),
.Y(n_473)
);

NAND2x1_ASAP7_75t_L g492 ( 
.A(n_473),
.B(n_480),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_439),
.B(n_402),
.C(n_420),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_474),
.B(n_475),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_451),
.B(n_424),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_476),
.A2(n_425),
.B1(n_457),
.B2(n_405),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_439),
.B(n_412),
.C(n_406),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_477),
.B(n_433),
.Y(n_487)
);

AO22x1_ASAP7_75t_SL g479 ( 
.A1(n_440),
.A2(n_443),
.B1(n_334),
.B2(n_458),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_450),
.B(n_425),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_461),
.B(n_456),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_481),
.B(n_489),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_483),
.A2(n_486),
.B1(n_469),
.B2(n_478),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_480),
.A2(n_475),
.B1(n_459),
.B2(n_467),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_487),
.B(n_490),
.Y(n_499)
);

FAx1_ASAP7_75t_L g488 ( 
.A(n_479),
.B(n_394),
.CI(n_453),
.CON(n_488),
.SN(n_488)
);

A2O1A1Ixp33_ASAP7_75t_SL g500 ( 
.A1(n_488),
.A2(n_478),
.B(n_471),
.C(n_459),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_477),
.B(n_434),
.C(n_433),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_462),
.B(n_463),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_468),
.B(n_463),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_493),
.B(n_460),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_473),
.A2(n_388),
.B(n_399),
.Y(n_494)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_494),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_474),
.B(n_460),
.C(n_479),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_495),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_465),
.B(n_419),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_497),
.B(n_467),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_498),
.B(n_502),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_500),
.B(n_503),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_493),
.B(n_470),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_489),
.B(n_466),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_504),
.A2(n_508),
.B(n_510),
.Y(n_512)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_505),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_496),
.B(n_469),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_507),
.B(n_511),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_484),
.B(n_398),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_482),
.B(n_344),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_492),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_503),
.A2(n_491),
.B1(n_485),
.B2(n_495),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_514),
.B(n_517),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_508),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_499),
.A2(n_509),
.B(n_506),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_519),
.A2(n_520),
.B(n_521),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_501),
.A2(n_492),
.B(n_488),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_500),
.A2(n_488),
.B(n_483),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_515),
.B(n_486),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_523),
.B(n_524),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_518),
.B(n_482),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_513),
.B(n_500),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_526),
.B(n_527),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_512),
.A2(n_494),
.B1(n_352),
.B2(n_353),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_525),
.B(n_516),
.C(n_359),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_528),
.B(n_530),
.C(n_348),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_522),
.A2(n_516),
.B(n_359),
.Y(n_530)
);

NAND3xp33_ASAP7_75t_L g532 ( 
.A(n_531),
.B(n_348),
.C(n_382),
.Y(n_532)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_532),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_534),
.A2(n_529),
.B(n_533),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_535),
.B(n_382),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_536),
.B(n_382),
.Y(n_537)
);


endmodule