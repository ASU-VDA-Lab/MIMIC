module real_aes_239_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_815;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_0), .B(n_129), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_1), .A2(n_138), .B(n_143), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_2), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g819 ( .A(n_3), .Y(n_819) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_4), .B(n_145), .Y(n_184) );
INVx1_ASAP7_75t_L g136 ( .A(n_5), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_6), .B(n_145), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_7), .B(n_156), .Y(n_490) );
INVx1_ASAP7_75t_L g510 ( .A(n_8), .Y(n_510) );
CKINVDCx16_ASAP7_75t_R g452 ( .A(n_9), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g524 ( .A(n_10), .Y(n_524) );
NAND2xp33_ASAP7_75t_L g207 ( .A(n_11), .B(n_147), .Y(n_207) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_12), .A2(n_38), .B1(n_440), .B2(n_441), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_12), .Y(n_441) );
INVx2_ASAP7_75t_L g126 ( .A(n_13), .Y(n_126) );
AOI221x1_ASAP7_75t_L g231 ( .A1(n_14), .A2(n_28), .B1(n_129), .B2(n_138), .C(n_232), .Y(n_231) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_15), .Y(n_107) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_16), .B(n_129), .Y(n_203) );
AO21x2_ASAP7_75t_L g200 ( .A1(n_17), .A2(n_201), .B(n_202), .Y(n_200) );
INVx1_ASAP7_75t_L g499 ( .A(n_18), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_19), .B(n_149), .Y(n_235) );
XOR2xp5_ASAP7_75t_L g809 ( .A(n_20), .B(n_810), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_21), .B(n_145), .Y(n_160) );
AO21x1_ASAP7_75t_L g179 ( .A1(n_22), .A2(n_129), .B(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g111 ( .A(n_23), .Y(n_111) );
OAI22xp5_ASAP7_75t_L g810 ( .A1(n_24), .A2(n_59), .B1(n_811), .B2(n_812), .Y(n_810) );
CKINVDCx16_ASAP7_75t_R g812 ( .A(n_24), .Y(n_812) );
INVx1_ASAP7_75t_L g497 ( .A(n_25), .Y(n_497) );
INVx1_ASAP7_75t_SL g565 ( .A(n_26), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_27), .B(n_130), .Y(n_484) );
NAND2x1_ASAP7_75t_L g224 ( .A(n_29), .B(n_145), .Y(n_224) );
AOI33xp33_ASAP7_75t_L g543 ( .A1(n_30), .A2(n_55), .A3(n_472), .B1(n_481), .B2(n_544), .B3(n_545), .Y(n_543) );
NAND2x1_ASAP7_75t_L g170 ( .A(n_31), .B(n_147), .Y(n_170) );
INVx1_ASAP7_75t_L g518 ( .A(n_32), .Y(n_518) );
OA21x2_ASAP7_75t_L g125 ( .A1(n_33), .A2(n_89), .B(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g151 ( .A(n_33), .B(n_89), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_34), .B(n_508), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_35), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_36), .B(n_145), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_37), .B(n_147), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_38), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_39), .A2(n_138), .B(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g135 ( .A(n_40), .B(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g139 ( .A(n_40), .B(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g480 ( .A(n_40), .Y(n_480) );
OR2x6_ASAP7_75t_L g109 ( .A(n_41), .B(n_110), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_42), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_43), .B(n_129), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_44), .B(n_508), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g468 ( .A1(n_45), .A2(n_124), .B1(n_156), .B2(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_46), .B(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_47), .B(n_130), .Y(n_566) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_48), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_49), .B(n_147), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_50), .B(n_201), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_51), .B(n_130), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_52), .A2(n_138), .B(n_169), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g476 ( .A(n_53), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_54), .B(n_147), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_56), .B(n_130), .Y(n_536) );
INVx1_ASAP7_75t_L g132 ( .A(n_57), .Y(n_132) );
INVx1_ASAP7_75t_L g142 ( .A(n_57), .Y(n_142) );
AND2x2_ASAP7_75t_L g537 ( .A(n_58), .B(n_149), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g811 ( .A(n_59), .Y(n_811) );
AOI221xp5_ASAP7_75t_L g507 ( .A1(n_60), .A2(n_76), .B1(n_478), .B2(n_508), .C(n_509), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_61), .B(n_508), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_62), .B(n_145), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_63), .B(n_124), .Y(n_526) );
AOI21xp5_ASAP7_75t_SL g554 ( .A1(n_64), .A2(n_478), .B(n_555), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_65), .A2(n_138), .B(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g493 ( .A(n_66), .Y(n_493) );
AO21x1_ASAP7_75t_L g181 ( .A1(n_67), .A2(n_138), .B(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g128 ( .A(n_68), .B(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g535 ( .A(n_69), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_70), .B(n_129), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_71), .A2(n_478), .B(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g196 ( .A(n_72), .B(n_150), .Y(n_196) );
INVx1_ASAP7_75t_L g134 ( .A(n_73), .Y(n_134) );
INVx1_ASAP7_75t_L g140 ( .A(n_73), .Y(n_140) );
AND2x2_ASAP7_75t_L g174 ( .A(n_74), .B(n_123), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_75), .B(n_508), .Y(n_546) );
AND2x2_ASAP7_75t_L g567 ( .A(n_77), .B(n_123), .Y(n_567) );
INVx1_ASAP7_75t_L g494 ( .A(n_78), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_79), .A2(n_478), .B(n_564), .Y(n_563) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_80), .A2(n_478), .B(n_483), .C(n_488), .Y(n_477) );
INVx1_ASAP7_75t_L g112 ( .A(n_81), .Y(n_112) );
AND2x2_ASAP7_75t_L g122 ( .A(n_82), .B(n_123), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_83), .B(n_129), .Y(n_162) );
AND2x2_ASAP7_75t_SL g552 ( .A(n_84), .B(n_123), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_85), .B(n_445), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_86), .A2(n_478), .B1(n_541), .B2(n_542), .Y(n_540) );
AND2x2_ASAP7_75t_L g180 ( .A(n_87), .B(n_156), .Y(n_180) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_88), .A2(n_103), .B1(n_447), .B2(n_454), .C1(n_823), .C2(n_828), .Y(n_102) );
AOI22xp5_ASAP7_75t_L g113 ( .A1(n_88), .A2(n_114), .B1(n_442), .B2(n_443), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g443 ( .A(n_88), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_90), .B(n_147), .Y(n_161) );
AND2x2_ASAP7_75t_L g227 ( .A(n_91), .B(n_123), .Y(n_227) );
INVx1_ASAP7_75t_L g556 ( .A(n_92), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_93), .B(n_145), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_94), .A2(n_138), .B(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_95), .B(n_147), .Y(n_233) );
AND2x2_ASAP7_75t_L g547 ( .A(n_96), .B(n_123), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_97), .B(n_145), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_98), .A2(n_516), .B(n_517), .C(n_519), .Y(n_515) );
BUFx2_ASAP7_75t_L g453 ( .A(n_99), .Y(n_453) );
BUFx2_ASAP7_75t_SL g832 ( .A(n_99), .Y(n_832) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_100), .A2(n_138), .B(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_101), .B(n_130), .Y(n_557) );
OAI21x1_ASAP7_75t_SL g103 ( .A1(n_104), .A2(n_113), .B(n_444), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
BUFx2_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
BUFx2_ASAP7_75t_L g446 ( .A(n_106), .Y(n_446) );
BUFx2_ASAP7_75t_L g834 ( .A(n_106), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
OR2x6_ASAP7_75t_SL g459 ( .A(n_107), .B(n_108), .Y(n_459) );
AND2x6_ASAP7_75t_SL g808 ( .A(n_107), .B(n_109), .Y(n_808) );
OR2x2_ASAP7_75t_L g822 ( .A(n_107), .B(n_109), .Y(n_822) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
INVx2_ASAP7_75t_L g442 ( .A(n_114), .Y(n_442) );
XNOR2x1_ASAP7_75t_L g114 ( .A(n_115), .B(n_439), .Y(n_114) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_115), .A2(n_457), .B1(n_460), .B2(n_807), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_115), .A2(n_458), .B1(n_460), .B2(n_815), .Y(n_814) );
AND2x4_ASAP7_75t_L g115 ( .A(n_116), .B(n_324), .Y(n_115) );
NOR3xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_279), .C(n_308), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g117 ( .A(n_118), .B(n_252), .Y(n_117) );
AOI221xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_175), .B1(n_197), .B2(n_209), .C(n_213), .Y(n_118) );
INVx3_ASAP7_75t_SL g369 ( .A(n_119), .Y(n_369) );
AND2x2_ASAP7_75t_SL g119 ( .A(n_120), .B(n_152), .Y(n_119) );
NAND2x1p5_ASAP7_75t_L g215 ( .A(n_120), .B(n_165), .Y(n_215) );
INVx4_ASAP7_75t_L g250 ( .A(n_120), .Y(n_250) );
AND2x2_ASAP7_75t_L g272 ( .A(n_120), .B(n_166), .Y(n_272) );
AND2x2_ASAP7_75t_L g278 ( .A(n_120), .B(n_217), .Y(n_278) );
INVx5_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g247 ( .A(n_121), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_121), .B(n_165), .Y(n_323) );
AND2x2_ASAP7_75t_L g328 ( .A(n_121), .B(n_166), .Y(n_328) );
AND2x2_ASAP7_75t_L g340 ( .A(n_121), .B(n_200), .Y(n_340) );
NOR2x1_ASAP7_75t_SL g379 ( .A(n_121), .B(n_217), .Y(n_379) );
OR2x6_ASAP7_75t_L g121 ( .A(n_122), .B(n_127), .Y(n_121) );
INVx3_ASAP7_75t_L g195 ( .A(n_123), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_123), .A2(n_195), .B1(n_515), .B2(n_520), .Y(n_514) );
INVx4_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_124), .B(n_523), .Y(n_522) );
INVx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx4f_ASAP7_75t_L g201 ( .A(n_125), .Y(n_201) );
AND2x2_ASAP7_75t_SL g150 ( .A(n_126), .B(n_151), .Y(n_150) );
AND2x4_ASAP7_75t_L g156 ( .A(n_126), .B(n_151), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_137), .B(n_149), .Y(n_127) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_135), .Y(n_129) );
INVx1_ASAP7_75t_L g495 ( .A(n_130), .Y(n_495) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_133), .Y(n_130) );
AND2x6_ASAP7_75t_L g147 ( .A(n_131), .B(n_140), .Y(n_147) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x4_ASAP7_75t_L g145 ( .A(n_133), .B(n_142), .Y(n_145) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx5_ASAP7_75t_L g148 ( .A(n_135), .Y(n_148) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_135), .Y(n_519) );
AND2x2_ASAP7_75t_L g141 ( .A(n_136), .B(n_142), .Y(n_141) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_136), .Y(n_473) );
AND2x6_ASAP7_75t_L g138 ( .A(n_139), .B(n_141), .Y(n_138) );
BUFx3_ASAP7_75t_L g475 ( .A(n_139), .Y(n_475) );
INVx2_ASAP7_75t_L g482 ( .A(n_140), .Y(n_482) );
AND2x4_ASAP7_75t_L g478 ( .A(n_141), .B(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g472 ( .A(n_142), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_146), .B(n_148), .Y(n_143) );
INVxp67_ASAP7_75t_L g500 ( .A(n_145), .Y(n_500) );
INVxp67_ASAP7_75t_L g498 ( .A(n_147), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_148), .A2(n_160), .B(n_161), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_148), .A2(n_170), .B(n_171), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_148), .A2(n_183), .B(n_184), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_148), .A2(n_192), .B(n_193), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_148), .A2(n_206), .B(n_207), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_148), .A2(n_224), .B(n_225), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_148), .A2(n_233), .B(n_234), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_148), .A2(n_484), .B(n_485), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_148), .B(n_156), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_SL g509 ( .A1(n_148), .A2(n_487), .B(n_510), .C(n_511), .Y(n_509) );
O2A1O1Ixp33_ASAP7_75t_L g534 ( .A1(n_148), .A2(n_487), .B(n_535), .C(n_536), .Y(n_534) );
INVx1_ASAP7_75t_L g541 ( .A(n_148), .Y(n_541) );
O2A1O1Ixp33_ASAP7_75t_L g555 ( .A1(n_148), .A2(n_487), .B(n_556), .C(n_557), .Y(n_555) );
O2A1O1Ixp33_ASAP7_75t_SL g564 ( .A1(n_148), .A2(n_487), .B(n_565), .C(n_566), .Y(n_564) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_149), .Y(n_173) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_149), .A2(n_231), .B(n_235), .Y(n_230) );
OA21x2_ASAP7_75t_L g275 ( .A1(n_149), .A2(n_231), .B(n_235), .Y(n_275) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g208 ( .A(n_152), .Y(n_208) );
AND2x2_ASAP7_75t_L g312 ( .A(n_152), .B(n_261), .Y(n_312) );
AND2x2_ASAP7_75t_L g409 ( .A(n_152), .B(n_340), .Y(n_409) );
AND2x4_ASAP7_75t_L g152 ( .A(n_153), .B(n_165), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g241 ( .A(n_154), .Y(n_241) );
INVx2_ASAP7_75t_L g263 ( .A(n_154), .Y(n_263) );
AO21x2_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_157), .B(n_163), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_155), .B(n_164), .Y(n_163) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_155), .A2(n_157), .B(n_163), .Y(n_217) );
INVx1_ASAP7_75t_SL g155 ( .A(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_156), .B(n_186), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_156), .A2(n_203), .B(n_204), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_156), .A2(n_554), .B(n_558), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_158), .B(n_162), .Y(n_157) );
AND2x2_ASAP7_75t_L g238 ( .A(n_165), .B(n_199), .Y(n_238) );
INVx2_ASAP7_75t_L g242 ( .A(n_165), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_165), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g341 ( .A(n_165), .B(n_306), .Y(n_341) );
OR2x2_ASAP7_75t_L g388 ( .A(n_165), .B(n_200), .Y(n_388) );
INVx4_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_166), .Y(n_338) );
AO21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_173), .B(n_174), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_168), .B(n_172), .Y(n_167) );
AO21x2_ASAP7_75t_L g560 ( .A1(n_173), .A2(n_561), .B(n_567), .Y(n_560) );
AND2x2_ASAP7_75t_L g385 ( .A(n_175), .B(n_266), .Y(n_385) );
AND2x2_ASAP7_75t_L g435 ( .A(n_175), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
OR2x2_ASAP7_75t_L g311 ( .A(n_176), .B(n_255), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_177), .B(n_187), .Y(n_176) );
AND2x2_ASAP7_75t_L g244 ( .A(n_177), .B(n_245), .Y(n_244) );
OR2x2_ASAP7_75t_L g274 ( .A(n_177), .B(n_275), .Y(n_274) );
AND2x4_ASAP7_75t_L g295 ( .A(n_177), .B(n_275), .Y(n_295) );
AND2x4_ASAP7_75t_L g330 ( .A(n_177), .B(n_318), .Y(n_330) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g211 ( .A(n_178), .Y(n_211) );
OAI21x1_ASAP7_75t_SL g178 ( .A1(n_179), .A2(n_181), .B(n_185), .Y(n_178) );
INVx1_ASAP7_75t_L g186 ( .A(n_180), .Y(n_186) );
AND2x2_ASAP7_75t_L g257 ( .A(n_187), .B(n_210), .Y(n_257) );
AND2x2_ASAP7_75t_L g343 ( .A(n_187), .B(n_275), .Y(n_343) );
AND2x2_ASAP7_75t_L g354 ( .A(n_187), .B(n_219), .Y(n_354) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g218 ( .A(n_188), .B(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g285 ( .A(n_188), .B(n_220), .Y(n_285) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_195), .B(n_196), .Y(n_188) );
AO21x2_ASAP7_75t_L g212 ( .A1(n_189), .A2(n_195), .B(n_196), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_190), .B(n_194), .Y(n_189) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_195), .A2(n_221), .B(n_227), .Y(n_220) );
AO21x2_ASAP7_75t_L g245 ( .A1(n_195), .A2(n_221), .B(n_227), .Y(n_245) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_195), .A2(n_531), .B(n_537), .Y(n_530) );
AO21x2_ASAP7_75t_L g584 ( .A1(n_195), .A2(n_531), .B(n_537), .Y(n_584) );
INVx2_ASAP7_75t_SL g197 ( .A(n_198), .Y(n_197) );
OR2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_208), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_199), .B(n_250), .Y(n_307) );
AND2x2_ASAP7_75t_L g351 ( .A(n_199), .B(n_217), .Y(n_351) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_200), .B(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g261 ( .A(n_200), .Y(n_261) );
BUFx3_ASAP7_75t_L g270 ( .A(n_200), .Y(n_270) );
AND2x2_ASAP7_75t_L g293 ( .A(n_200), .B(n_263), .Y(n_293) );
INVx2_ASAP7_75t_SL g488 ( .A(n_201), .Y(n_488) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_201), .A2(n_507), .B(n_512), .Y(n_506) );
OAI322xp33_ASAP7_75t_L g213 ( .A1(n_208), .A2(n_214), .A3(n_218), .B1(n_228), .B2(n_236), .C1(n_243), .C2(n_248), .Y(n_213) );
INVx1_ASAP7_75t_L g374 ( .A(n_208), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_209), .B(n_249), .Y(n_248) );
AND2x4_ASAP7_75t_L g287 ( .A(n_209), .B(n_229), .Y(n_287) );
INVx2_ASAP7_75t_L g332 ( .A(n_209), .Y(n_332) );
AND2x2_ASAP7_75t_L g348 ( .A(n_209), .B(n_290), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_209), .B(n_366), .Y(n_396) );
AND2x4_ASAP7_75t_L g209 ( .A(n_210), .B(n_212), .Y(n_209) );
AND2x2_ASAP7_75t_SL g299 ( .A(n_210), .B(n_275), .Y(n_299) );
OR2x2_ASAP7_75t_L g320 ( .A(n_210), .B(n_237), .Y(n_320) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
BUFx2_ASAP7_75t_L g292 ( .A(n_211), .Y(n_292) );
INVx2_ASAP7_75t_L g237 ( .A(n_212), .Y(n_237) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_212), .Y(n_239) );
OR2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
INVx2_ASAP7_75t_L g282 ( .A(n_215), .Y(n_282) );
INVxp67_ASAP7_75t_SL g302 ( .A(n_216), .Y(n_302) );
INVx1_ASAP7_75t_L g400 ( .A(n_216), .Y(n_400) );
INVxp67_ASAP7_75t_SL g415 ( .A(n_216), .Y(n_415) );
NAND2x1_ASAP7_75t_L g425 ( .A(n_218), .B(n_229), .Y(n_425) );
INVx1_ASAP7_75t_L g432 ( .A(n_218), .Y(n_432) );
BUFx2_ASAP7_75t_L g266 ( .A(n_219), .Y(n_266) );
AND2x2_ASAP7_75t_L g342 ( .A(n_219), .B(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
BUFx3_ASAP7_75t_L g251 ( .A(n_220), .Y(n_251) );
INVxp67_ASAP7_75t_L g255 ( .A(n_220), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_222), .B(n_226), .Y(n_221) );
NAND3xp33_ASAP7_75t_L g243 ( .A(n_228), .B(n_244), .C(n_246), .Y(n_243) );
INVx1_ASAP7_75t_SL g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_SL g264 ( .A(n_229), .B(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_229), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g416 ( .A(n_229), .B(n_365), .Y(n_416) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx2_ASAP7_75t_L g318 ( .A(n_230), .Y(n_318) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_230), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B1(n_239), .B2(n_240), .Y(n_236) );
AND2x4_ASAP7_75t_SL g365 ( .A(n_237), .B(n_245), .Y(n_365) );
AND2x2_ASAP7_75t_L g378 ( .A(n_238), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_239), .Y(n_380) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
INVx2_ASAP7_75t_L g337 ( .A(n_241), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_241), .B(n_250), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_242), .B(n_260), .Y(n_259) );
AND3x2_ASAP7_75t_L g277 ( .A(n_242), .B(n_270), .C(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g301 ( .A(n_242), .Y(n_301) );
AND2x2_ASAP7_75t_L g414 ( .A(n_242), .B(n_415), .Y(n_414) );
BUFx2_ASAP7_75t_L g290 ( .A(n_245), .Y(n_290) );
INVx1_ASAP7_75t_L g368 ( .A(n_245), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_246), .B(n_269), .Y(n_407) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_247), .B(n_351), .Y(n_356) );
AND2x4_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
AND2x2_ASAP7_75t_L g347 ( .A(n_250), .B(n_293), .Y(n_347) );
INVx1_ASAP7_75t_SL g298 ( .A(n_251), .Y(n_298) );
AND2x2_ASAP7_75t_L g406 ( .A(n_251), .B(n_318), .Y(n_406) );
AND2x2_ASAP7_75t_L g427 ( .A(n_251), .B(n_299), .Y(n_427) );
AOI221xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_258), .B1(n_264), .B2(n_267), .C(n_273), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
INVx1_ASAP7_75t_L g419 ( .A(n_255), .Y(n_419) );
AOI21xp33_ASAP7_75t_SL g273 ( .A1(n_256), .A2(n_274), .B(n_276), .Y(n_273) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g265 ( .A(n_257), .B(n_266), .Y(n_265) );
AOI222xp33_ASAP7_75t_L g288 ( .A1(n_257), .A2(n_289), .B1(n_291), .B2(n_296), .C1(n_300), .C2(n_303), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_257), .B(n_406), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g309 ( .A1(n_258), .A2(n_287), .B1(n_310), .B2(n_312), .Y(n_309) );
INVx1_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx1_ASAP7_75t_L g294 ( .A(n_261), .Y(n_294) );
AND2x2_ASAP7_75t_L g413 ( .A(n_261), .B(n_379), .Y(n_413) );
OAI32xp33_ASAP7_75t_L g417 ( .A1(n_261), .A2(n_286), .A3(n_338), .B1(n_346), .B2(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g422 ( .A(n_261), .B(n_272), .Y(n_422) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g306 ( .A(n_263), .Y(n_306) );
OAI21xp5_ASAP7_75t_SL g313 ( .A1(n_264), .A2(n_314), .B(n_321), .Y(n_313) );
INVx1_ASAP7_75t_L g377 ( .A(n_266), .Y(n_377) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
AND2x2_ASAP7_75t_L g281 ( .A(n_269), .B(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx2_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g289 ( .A(n_272), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g362 ( .A(n_272), .B(n_293), .Y(n_362) );
INVx1_ASAP7_75t_SL g433 ( .A(n_274), .Y(n_433) );
AND2x2_ASAP7_75t_L g367 ( .A(n_275), .B(n_368), .Y(n_367) );
OAI222xp33_ASAP7_75t_L g420 ( .A1(n_276), .A2(n_329), .B1(n_408), .B2(n_421), .C1(n_423), .C2(n_425), .Y(n_420) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x4_ASAP7_75t_L g393 ( .A(n_278), .B(n_394), .Y(n_393) );
OAI21xp33_ASAP7_75t_SL g279 ( .A1(n_280), .A2(n_283), .B(n_288), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_282), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx1_ASAP7_75t_L g361 ( .A(n_284), .Y(n_361) );
INVx1_ASAP7_75t_L g329 ( .A(n_285), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_285), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g383 ( .A(n_290), .Y(n_383) );
AO22x1_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_293), .B1(n_294), .B2(n_295), .Y(n_291) );
OAI322xp33_ASAP7_75t_L g403 ( .A1(n_292), .A2(n_353), .A3(n_356), .B1(n_404), .B2(n_405), .C1(n_407), .C2(n_408), .Y(n_403) );
AND2x2_ASAP7_75t_SL g327 ( .A(n_293), .B(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g322 ( .A(n_294), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_SL g382 ( .A(n_295), .B(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g424 ( .A(n_295), .B(n_354), .Y(n_424) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
INVx1_ASAP7_75t_L g404 ( .A(n_298), .Y(n_404) );
INVx1_ASAP7_75t_SL g333 ( .A(n_299), .Y(n_333) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
OR2x2_ASAP7_75t_L g335 ( .A(n_307), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g373 ( .A(n_307), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_313), .Y(n_308) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_319), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g346 ( .A(n_317), .B(n_332), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_317), .B(n_354), .Y(n_353) );
BUFx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g376 ( .A(n_320), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NOR2x1_ASAP7_75t_L g324 ( .A(n_325), .B(n_389), .Y(n_324) );
NAND4xp25_ASAP7_75t_L g325 ( .A(n_326), .B(n_344), .C(n_357), .D(n_370), .Y(n_325) );
AOI322xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_329), .A3(n_330), .B1(n_331), .B2(n_334), .C1(n_339), .C2(n_342), .Y(n_326) );
AOI211xp5_ASAP7_75t_L g426 ( .A1(n_327), .A2(n_427), .B(n_428), .C(n_431), .Y(n_426) );
AND2x2_ASAP7_75t_L g438 ( .A(n_328), .B(n_415), .Y(n_438) );
INVx1_ASAP7_75t_L g360 ( .A(n_330), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_330), .B(n_365), .Y(n_402) );
NAND2xp33_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_338), .B(n_351), .Y(n_418) );
AND2x4_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
AOI222xp33_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_347), .B1(n_348), .B2(n_349), .C1(n_352), .C2(n_355), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AOI221xp5_ASAP7_75t_L g357 ( .A1(n_347), .A2(n_358), .B1(n_361), .B2(n_362), .C(n_363), .Y(n_357) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AOI21xp33_ASAP7_75t_SL g363 ( .A1(n_364), .A2(n_366), .B(n_369), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
AOI221xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_375), .B1(n_378), .B2(n_380), .C(n_381), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_SL g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g430 ( .A(n_379), .Y(n_430) );
AOI21xp33_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_384), .B(n_386), .Y(n_381) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
OR2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
INVx2_ASAP7_75t_L g394 ( .A(n_388), .Y(n_394) );
OR2x2_ASAP7_75t_L g429 ( .A(n_388), .B(n_430), .Y(n_429) );
NAND3xp33_ASAP7_75t_L g389 ( .A(n_390), .B(n_410), .C(n_426), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_403), .Y(n_390) );
OAI21xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_395), .B(n_397), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_401), .Y(n_397) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_416), .B1(n_417), .B2(n_419), .C(n_420), .Y(n_410) );
INVxp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NOR2x1_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_425), .B(n_429), .Y(n_428) );
O2A1O1Ixp33_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_433), .B(n_434), .C(n_437), .Y(n_431) );
INVxp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g824 ( .A(n_446), .B(n_825), .Y(n_824) );
INVx1_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_SL g450 ( .A(n_451), .B(n_453), .Y(n_450) );
INVx2_ASAP7_75t_L g827 ( .A(n_451), .Y(n_827) );
AOI21xp5_ASAP7_75t_L g829 ( .A1(n_451), .A2(n_830), .B(n_833), .Y(n_829) );
NAND2xp5_ASAP7_75t_SL g826 ( .A(n_453), .B(n_827), .Y(n_826) );
INVxp33_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
AOI221xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_809), .B1(n_813), .B2(n_817), .C(n_818), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_458), .Y(n_457) );
CKINVDCx11_ASAP7_75t_R g458 ( .A(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_741), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_462), .B(n_664), .Y(n_461) );
NAND3xp33_ASAP7_75t_L g462 ( .A(n_463), .B(n_611), .C(n_644), .Y(n_462) );
AOI211xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_568), .B(n_577), .C(n_601), .Y(n_463) );
OAI21xp33_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_502), .B(n_548), .Y(n_464) );
OR2x2_ASAP7_75t_L g621 ( .A(n_465), .B(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g776 ( .A(n_465), .B(n_777), .Y(n_776) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AOI22xp33_ASAP7_75t_SL g666 ( .A1(n_466), .A2(n_667), .B1(n_671), .B2(n_673), .Y(n_666) );
AND2x2_ASAP7_75t_L g703 ( .A(n_466), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_489), .Y(n_466) );
INVx1_ASAP7_75t_L g600 ( .A(n_467), .Y(n_600) );
AND2x4_ASAP7_75t_L g617 ( .A(n_467), .B(n_598), .Y(n_617) );
INVx2_ASAP7_75t_L g639 ( .A(n_467), .Y(n_639) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_467), .Y(n_722) );
AND2x2_ASAP7_75t_L g793 ( .A(n_467), .B(n_551), .Y(n_793) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_477), .Y(n_467) );
NOR3xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_474), .C(n_476), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AND2x4_ASAP7_75t_L g508 ( .A(n_471), .B(n_475), .Y(n_508) );
AND2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
OR2x6_ASAP7_75t_L g487 ( .A(n_472), .B(n_482), .Y(n_487) );
INVxp33_ASAP7_75t_L g544 ( .A(n_472), .Y(n_544) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVxp67_ASAP7_75t_L g525 ( .A(n_478), .Y(n_525) );
NOR2x1p5_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
INVx1_ASAP7_75t_L g545 ( .A(n_481), .Y(n_545) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_487), .A2(n_493), .B1(n_494), .B2(n_495), .Y(n_492) );
INVxp67_ASAP7_75t_L g516 ( .A(n_487), .Y(n_516) );
AO21x2_ASAP7_75t_L g538 ( .A1(n_488), .A2(n_539), .B(n_547), .Y(n_538) );
AO21x2_ASAP7_75t_L g582 ( .A1(n_488), .A2(n_539), .B(n_547), .Y(n_582) );
AND2x2_ASAP7_75t_L g559 ( .A(n_489), .B(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g587 ( .A(n_489), .Y(n_587) );
INVx3_ASAP7_75t_L g598 ( .A(n_489), .Y(n_598) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
OAI21xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_496), .B(n_501), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_495), .B(n_518), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B1(n_499), .B2(n_500), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_502), .A2(n_788), .B1(n_790), .B2(n_792), .Y(n_787) );
NAND2xp5_ASAP7_75t_SL g798 ( .A(n_502), .B(n_799), .Y(n_798) );
INVx2_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_528), .Y(n_503) );
INVx3_ASAP7_75t_L g571 ( .A(n_504), .Y(n_571) );
AND2x2_ASAP7_75t_L g579 ( .A(n_504), .B(n_580), .Y(n_579) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_504), .Y(n_609) );
NAND2x1_ASAP7_75t_SL g803 ( .A(n_504), .B(n_570), .Y(n_803) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_513), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g576 ( .A(n_506), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_506), .B(n_582), .Y(n_594) );
AND2x2_ASAP7_75t_L g607 ( .A(n_506), .B(n_513), .Y(n_607) );
AND2x4_ASAP7_75t_L g614 ( .A(n_506), .B(n_615), .Y(n_614) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_506), .Y(n_663) );
INVxp67_ASAP7_75t_L g670 ( .A(n_506), .Y(n_670) );
INVx1_ASAP7_75t_L g675 ( .A(n_506), .Y(n_675) );
INVx1_ASAP7_75t_L g527 ( .A(n_508), .Y(n_527) );
INVx1_ASAP7_75t_L g574 ( .A(n_513), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_513), .B(n_584), .Y(n_593) );
INVx2_ASAP7_75t_L g661 ( .A(n_513), .Y(n_661) );
INVx1_ASAP7_75t_L g700 ( .A(n_513), .Y(n_700) );
OR2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_521), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_525), .B1(n_526), .B2(n_527), .Y(n_521) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g630 ( .A(n_528), .B(n_607), .Y(n_630) );
AND2x2_ASAP7_75t_L g698 ( .A(n_528), .B(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g712 ( .A(n_528), .B(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_528), .B(n_727), .Y(n_726) );
AND2x4_ASAP7_75t_L g528 ( .A(n_529), .B(n_538), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NOR2x1_ASAP7_75t_L g575 ( .A(n_530), .B(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g668 ( .A(n_530), .B(n_661), .Y(n_668) );
AND2x2_ASAP7_75t_L g759 ( .A(n_530), .B(n_581), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
INVx1_ASAP7_75t_L g570 ( .A(n_538), .Y(n_570) );
INVx2_ASAP7_75t_L g615 ( .A(n_538), .Y(n_615) );
AND2x2_ASAP7_75t_L g660 ( .A(n_538), .B(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_540), .B(n_546), .Y(n_539) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_559), .Y(n_549) );
AND2x2_ASAP7_75t_L g702 ( .A(n_550), .B(n_703), .Y(n_702) );
OR2x6_ASAP7_75t_L g761 ( .A(n_550), .B(n_762), .Y(n_761) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx4_ASAP7_75t_L g591 ( .A(n_551), .Y(n_591) );
AND2x4_ASAP7_75t_L g599 ( .A(n_551), .B(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g634 ( .A(n_551), .B(n_560), .Y(n_634) );
INVx2_ASAP7_75t_L g683 ( .A(n_551), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g732 ( .A(n_551), .B(n_657), .Y(n_732) );
AND2x2_ASAP7_75t_L g769 ( .A(n_551), .B(n_587), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_551), .B(n_652), .Y(n_777) );
OR2x6_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
AND2x2_ASAP7_75t_L g610 ( .A(n_559), .B(n_599), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_559), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_SL g749 ( .A(n_559), .B(n_637), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_559), .B(n_650), .Y(n_771) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_560), .Y(n_589) );
AND2x2_ASAP7_75t_L g597 ( .A(n_560), .B(n_598), .Y(n_597) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_560), .Y(n_620) );
INVx2_ASAP7_75t_L g623 ( .A(n_560), .Y(n_623) );
INVx1_ASAP7_75t_L g656 ( .A(n_560), .Y(n_656) );
INVx1_ASAP7_75t_L g704 ( .A(n_560), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
NAND2xp33_ASAP7_75t_L g568 ( .A(n_569), .B(n_572), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_570), .B(n_573), .Y(n_646) );
OR2x2_ASAP7_75t_L g718 ( .A(n_570), .B(n_719), .Y(n_718) );
AND4x1_ASAP7_75t_SL g764 ( .A(n_570), .B(n_746), .C(n_765), .D(n_766), .Y(n_764) );
OR2x2_ASAP7_75t_L g788 ( .A(n_571), .B(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
AND2x2_ASAP7_75t_L g625 ( .A(n_574), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_574), .B(n_583), .Y(n_775) );
AND2x2_ASAP7_75t_L g800 ( .A(n_575), .B(n_660), .Y(n_800) );
OAI32xp33_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_585), .A3(n_590), .B1(n_592), .B2(n_595), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g673 ( .A(n_580), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g773 ( .A(n_580), .B(n_727), .Y(n_773) );
AND2x4_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
AND2x2_ASAP7_75t_L g669 ( .A(n_581), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g755 ( .A(n_581), .Y(n_755) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_582), .B(n_584), .Y(n_789) );
INVx3_ASAP7_75t_L g606 ( .A(n_583), .Y(n_606) );
NAND2x1p5_ASAP7_75t_L g784 ( .A(n_583), .B(n_711), .Y(n_784) );
INVx3_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_584), .Y(n_643) );
AND2x2_ASAP7_75t_L g662 ( .A(n_584), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g796 ( .A(n_586), .Y(n_796) );
NAND2x1_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g636 ( .A(n_587), .Y(n_636) );
NOR2x1_ASAP7_75t_L g737 ( .A(n_587), .B(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_590), .B(n_696), .Y(n_695) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g628 ( .A(n_591), .B(n_596), .Y(n_628) );
AND2x4_ASAP7_75t_L g650 ( .A(n_591), .B(n_600), .Y(n_650) );
AND2x4_ASAP7_75t_SL g721 ( .A(n_591), .B(n_722), .Y(n_721) );
NOR2x1_ASAP7_75t_L g747 ( .A(n_591), .B(n_672), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_592), .A2(n_715), .B1(n_718), .B2(n_720), .Y(n_714) );
OR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
INVx2_ASAP7_75t_SL g734 ( .A(n_593), .Y(n_734) );
INVx2_ASAP7_75t_L g626 ( .A(n_594), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_599), .Y(n_595) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_597), .B(n_603), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_597), .A2(n_733), .B1(n_736), .B2(n_739), .Y(n_735) );
INVx1_ASAP7_75t_L g657 ( .A(n_598), .Y(n_657) );
AND2x2_ASAP7_75t_L g680 ( .A(n_598), .B(n_639), .Y(n_680) );
INVx2_ASAP7_75t_L g603 ( .A(n_599), .Y(n_603) );
OAI21xp5_ASAP7_75t_SL g601 ( .A1(n_602), .A2(n_604), .B(n_608), .Y(n_601) );
INVx1_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_605), .A2(n_677), .B1(n_681), .B2(n_682), .Y(n_676) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_606), .B(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_606), .B(n_674), .Y(n_690) );
INVx1_ASAP7_75t_L g694 ( .A(n_606), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
NOR3xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_627), .C(n_631), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_616), .B1(n_621), .B2(n_624), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g641 ( .A(n_614), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g681 ( .A(n_614), .B(n_668), .Y(n_681) );
AND2x2_ASAP7_75t_L g733 ( .A(n_614), .B(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g750 ( .A(n_614), .B(n_700), .Y(n_750) );
AND2x2_ASAP7_75t_L g805 ( .A(n_614), .B(n_699), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
INVx4_ASAP7_75t_L g672 ( .A(n_617), .Y(n_672) );
AND2x2_ASAP7_75t_L g682 ( .A(n_617), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
BUFx2_ASAP7_75t_L g687 ( .A(n_620), .Y(n_687) );
AND2x2_ASAP7_75t_L g696 ( .A(n_620), .B(n_680), .Y(n_696) );
INVx1_ASAP7_75t_L g731 ( .A(n_622), .Y(n_731) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g652 ( .A(n_623), .Y(n_652) );
INVxp67_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_625), .B(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_626), .B(n_694), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_635), .B(n_640), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_633), .B(n_672), .Y(n_781) );
INVx2_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
AOI21xp33_ASAP7_75t_SL g644 ( .A1(n_636), .A2(n_645), .B(n_647), .Y(n_644) );
AND2x2_ASAP7_75t_L g791 ( .A(n_636), .B(n_650), .Y(n_791) );
AND2x4_ASAP7_75t_L g654 ( .A(n_637), .B(n_655), .Y(n_654) );
INVx2_ASAP7_75t_SL g688 ( .A(n_637), .Y(n_688) );
NAND2xp5_ASAP7_75t_SL g770 ( .A(n_637), .B(n_704), .Y(n_770) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AOI21xp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_653), .B(n_658), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_650), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_650), .B(n_655), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_651), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g713 ( .A(n_651), .Y(n_713) );
INVx1_ASAP7_75t_L g717 ( .A(n_651), .Y(n_717) );
AND2x2_ASAP7_75t_L g801 ( .A(n_651), .B(n_769), .Y(n_801) );
AND2x2_ASAP7_75t_L g804 ( .A(n_651), .B(n_721), .Y(n_804) );
INVx3_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AND2x4_ASAP7_75t_SL g655 ( .A(n_656), .B(n_657), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_656), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AND2x4_ASAP7_75t_L g659 ( .A(n_660), .B(n_662), .Y(n_659) );
INVx1_ASAP7_75t_L g783 ( .A(n_660), .Y(n_783) );
AND2x2_ASAP7_75t_L g674 ( .A(n_661), .B(n_675), .Y(n_674) );
NAND4xp75_ASAP7_75t_L g664 ( .A(n_665), .B(n_684), .C(n_705), .D(n_723), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_676), .Y(n_665) );
AND2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
NAND2x1p5_ASAP7_75t_L g754 ( .A(n_668), .B(n_755), .Y(n_754) );
NAND2x1p5_ASAP7_75t_L g740 ( .A(n_669), .B(n_734), .Y(n_740) );
NAND2xp5_ASAP7_75t_R g756 ( .A(n_672), .B(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g806 ( .A(n_672), .Y(n_806) );
INVx2_ASAP7_75t_L g719 ( .A(n_674), .Y(n_719) );
BUFx3_ASAP7_75t_L g711 ( .A(n_675), .Y(n_711) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
BUFx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g762 ( .A(n_680), .Y(n_762) );
AND2x2_ASAP7_75t_L g716 ( .A(n_682), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g738 ( .A(n_683), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_689), .B(n_691), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_688), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_687), .B(n_721), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_688), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_690), .Y(n_785) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_695), .B1(n_697), .B2(n_701), .Y(n_691) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
OA21x2_ASAP7_75t_L g706 ( .A1(n_699), .A2(n_707), .B(n_708), .Y(n_706) );
INVx1_ASAP7_75t_L g727 ( .A(n_699), .Y(n_727) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g758 ( .A(n_700), .B(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g766 ( .A(n_700), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_701), .B(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g736 ( .A(n_704), .B(n_737), .Y(n_736) );
AOI21xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_712), .B(n_714), .Y(n_705) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
OR2x2_ASAP7_75t_L g753 ( .A(n_710), .B(n_754), .Y(n_753) );
INVx3_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_717), .Y(n_765) );
INVx2_ASAP7_75t_SL g757 ( .A(n_721), .Y(n_757) );
AND2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_735), .Y(n_723) );
AOI22xp5_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_728), .B1(n_730), .B2(n_733), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g786 ( .A(n_730), .Y(n_786) );
NOR2x1_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
INVx3_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_742), .B(n_778), .Y(n_741) );
NAND3xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_751), .C(n_763), .Y(n_742) );
NOR2x1_ASAP7_75t_L g743 ( .A(n_744), .B(n_748), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
BUFx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
AND2x2_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
AOI22xp33_ASAP7_75t_SL g751 ( .A1(n_752), .A2(n_756), .B1(n_758), .B2(n_760), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
NOR3xp33_ASAP7_75t_L g763 ( .A(n_764), .B(n_767), .C(n_774), .Y(n_763) );
AOI21xp33_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_771), .B(n_772), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
NOR2xp33_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_779), .B(n_797), .Y(n_778) );
NOR3xp33_ASAP7_75t_L g779 ( .A(n_780), .B(n_787), .C(n_794), .Y(n_779) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_782), .B1(n_785), .B2(n_786), .Y(n_780) );
OR2x2_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .Y(n_782) );
NOR3xp33_ASAP7_75t_L g794 ( .A(n_788), .B(n_793), .C(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVxp67_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
AOI222xp33_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_801), .B1(n_802), .B2(n_804), .C1(n_805), .C2(n_806), .Y(n_797) );
INVx1_ASAP7_75t_SL g799 ( .A(n_800), .Y(n_799) );
INVx2_ASAP7_75t_SL g802 ( .A(n_803), .Y(n_802) );
CKINVDCx11_ASAP7_75t_R g807 ( .A(n_808), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g816 ( .A(n_808), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_809), .Y(n_817) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx3_ASAP7_75t_SL g815 ( .A(n_816), .Y(n_815) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .Y(n_818) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx3_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
BUFx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVxp67_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_SL g828 ( .A(n_829), .Y(n_828) );
CKINVDCx11_ASAP7_75t_R g830 ( .A(n_831), .Y(n_830) );
CKINVDCx8_ASAP7_75t_R g831 ( .A(n_832), .Y(n_831) );
INVx2_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
endmodule