module real_jpeg_9573_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_2),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_49),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_3),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_3),
.B(n_25),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_3),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_3),
.A2(n_26),
.B(n_41),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_3),
.A2(n_79),
.B1(n_81),
.B2(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_3),
.A2(n_29),
.B(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_3),
.B(n_29),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_3),
.A2(n_70),
.B1(n_72),
.B2(n_134),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_3),
.A2(n_25),
.B(n_66),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_4),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_4),
.A2(n_46),
.B1(n_47),
.B2(n_61),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_7),
.A2(n_35),
.B1(n_46),
.B2(n_47),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_148)
);

BUFx6f_ASAP7_75t_SL g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_SL g54 ( 
.A1(n_10),
.A2(n_29),
.B(n_55),
.C(n_56),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_10),
.B(n_29),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_11),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_12),
.A2(n_33),
.B1(n_81),
.B2(n_106),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_12),
.A2(n_33),
.B1(n_46),
.B2(n_47),
.Y(n_134)
);

BUFx10_ASAP7_75t_L g81 ( 
.A(n_13),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_15),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_15),
.A2(n_25),
.B1(n_26),
.B2(n_59),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_15),
.A2(n_46),
.B1(n_47),
.B2(n_59),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_110),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_108),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_74),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_19),
.B(n_74),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_53),
.C(n_62),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_20),
.A2(n_21),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_36),
.B1(n_37),
.B2(n_52),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_22),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_32),
.B2(n_34),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_23),
.A2(n_28),
.B1(n_34),
.B2(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_23),
.A2(n_28),
.B1(n_32),
.B2(n_155),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B(n_27),
.C(n_28),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_25),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_24),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_24),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_25),
.A2(n_26),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_28),
.B(n_79),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_29),
.B(n_31),
.Y(n_67)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_30),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_43),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_38),
.B(n_43),
.C(n_52),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_39),
.A2(n_102),
.B1(n_105),
.B2(n_107),
.Y(n_101)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_40),
.A2(n_42),
.B(n_81),
.C(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_42),
.A2(n_79),
.B(n_80),
.C(n_81),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_42),
.B(n_81),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_45),
.B1(n_48),
.B2(n_50),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_44),
.A2(n_45),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_46),
.B(n_57),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_46),
.B(n_139),
.Y(n_138)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_47),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_48),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_50),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_53),
.A2(n_62),
.B1(n_63),
.B2(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_53),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_56),
.B1(n_58),
.B2(n_60),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_54),
.A2(n_56),
.B1(n_123),
.B2(n_125),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_54),
.A2(n_56),
.B1(n_125),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_54),
.A2(n_56),
.B1(n_58),
.B2(n_148),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_55),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_56),
.B(n_79),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_60),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_69),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_64),
.B(n_69),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_70),
.A2(n_72),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_70),
.A2(n_72),
.B1(n_117),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_119),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_72),
.B(n_79),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_90),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_76),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_82),
.B2(n_83),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_81),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_87),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_101),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_98),
.B2(n_99),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_158),
.B(n_164),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_151),
.B(n_157),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_142),
.B(n_150),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_131),
.B(n_141),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_120),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_115),
.B(n_120),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_126),
.B2(n_130),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_121),
.B(n_130),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_124),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_126),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_136),
.B(n_140),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_135),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_143),
.B(n_144),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_145),
.B(n_152),
.Y(n_157)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_147),
.CI(n_149),
.CON(n_145),
.SN(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_152),
.Y(n_159)
);

FAx1_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_154),
.CI(n_156),
.CON(n_152),
.SN(n_152)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_159),
.B(n_160),
.Y(n_164)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);


endmodule