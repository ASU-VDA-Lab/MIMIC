module fake_netlist_6_1252_n_2116 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2116);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2116;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_343;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_1033;
wire n_462;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1202;
wire n_1030;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2111;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_206;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g197 ( 
.A(n_136),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_69),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_103),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_182),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_102),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_24),
.Y(n_202)
);

INVxp33_ASAP7_75t_SL g203 ( 
.A(n_122),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_191),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_118),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_159),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_100),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_66),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_36),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_163),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_21),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_71),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_174),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_2),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_167),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_83),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_140),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_194),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_190),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_137),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_84),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_187),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_195),
.Y(n_223)
);

BUFx10_ASAP7_75t_L g224 ( 
.A(n_79),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_71),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_152),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_183),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_4),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_148),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_16),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_106),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_72),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_105),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_45),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_172),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_80),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_139),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_65),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_84),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_76),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_3),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_121),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_7),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_2),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_58),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_50),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_132),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_53),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_115),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_80),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_185),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_20),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_46),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_108),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_33),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_21),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_170),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_39),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_69),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_60),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_120),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_119),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_155),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_15),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_128),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_52),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_109),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_186),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_96),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_53),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_45),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_178),
.Y(n_272)
);

INVxp33_ASAP7_75t_L g273 ( 
.A(n_57),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_97),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_24),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_6),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_26),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_193),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_63),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_68),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_51),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_59),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_177),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_19),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_196),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_82),
.Y(n_286)
);

BUFx5_ASAP7_75t_L g287 ( 
.A(n_87),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_125),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_112),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_52),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_35),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_87),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_83),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_93),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_70),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_124),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_104),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_154),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_129),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_56),
.Y(n_300)
);

BUFx2_ASAP7_75t_SL g301 ( 
.A(n_91),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_59),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_78),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_48),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_114),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_188),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_150),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_85),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_86),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_47),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_127),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_175),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_6),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_26),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_1),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_74),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_113),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_180),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_79),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_189),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_18),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_39),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_75),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_169),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_55),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_15),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_91),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_146),
.Y(n_328)
);

INVx2_ASAP7_75t_SL g329 ( 
.A(n_160),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_65),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_157),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_192),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_23),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_46),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_74),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_162),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_60),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_166),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_11),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_28),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_58),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_61),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_72),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_117),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_3),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_85),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_88),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_43),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_66),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_35),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_12),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_41),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_11),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_93),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_36),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_184),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_145),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_42),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_38),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_50),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_27),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_4),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_110),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_37),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_27),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_78),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_73),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_31),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_34),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_7),
.Y(n_370)
);

BUFx10_ASAP7_75t_L g371 ( 
.A(n_54),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_70),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_56),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_95),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_123),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_5),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_43),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_63),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_158),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_111),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_81),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_68),
.Y(n_382)
);

BUFx2_ASAP7_75t_SL g383 ( 
.A(n_25),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_133),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_81),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_23),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_42),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_51),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_92),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_88),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_99),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_12),
.Y(n_392)
);

INVxp33_ASAP7_75t_L g393 ( 
.A(n_290),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_287),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_287),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_199),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_200),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_287),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_287),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_201),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_218),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_287),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_290),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_367),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_204),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_287),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_210),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_205),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_287),
.B(n_0),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_287),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_367),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_287),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_287),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_215),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_213),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_214),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_220),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_214),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_213),
.B(n_0),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_226),
.B(n_1),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_205),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_291),
.Y(n_422)
);

INVxp33_ASAP7_75t_L g423 ( 
.A(n_198),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_222),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_219),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_241),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_226),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_214),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_223),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_231),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_214),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_214),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_233),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_214),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_219),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_235),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_291),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_214),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_248),
.Y(n_439)
);

INVxp33_ASAP7_75t_SL g440 ( 
.A(n_209),
.Y(n_440)
);

INVxp67_ASAP7_75t_SL g441 ( 
.A(n_248),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_257),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_247),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_248),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_313),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_313),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_291),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_249),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_313),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_241),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_269),
.B(n_5),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_251),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_208),
.Y(n_453)
);

INVxp33_ASAP7_75t_SL g454 ( 
.A(n_216),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_254),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_261),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_257),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_265),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_262),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_208),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_263),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_272),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_208),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_246),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_278),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_246),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_246),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_265),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_252),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_297),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_298),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_342),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_312),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_207),
.B(n_8),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_312),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_306),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_311),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_318),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_272),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_320),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_269),
.B(n_8),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_198),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_344),
.Y(n_483)
);

NOR2xp67_ASAP7_75t_L g484 ( 
.A(n_327),
.B(n_9),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_252),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_272),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_252),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_294),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_344),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_294),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_294),
.Y(n_491)
);

NOR2xp67_ASAP7_75t_L g492 ( 
.A(n_327),
.B(n_9),
.Y(n_492)
);

NAND2xp33_ASAP7_75t_SL g493 ( 
.A(n_393),
.B(n_273),
.Y(n_493)
);

NOR2x1_ASAP7_75t_L g494 ( 
.A(n_474),
.B(n_289),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_453),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_441),
.B(n_207),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_426),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_441),
.B(n_289),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_401),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_396),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_416),
.Y(n_501)
);

AND3x2_ASAP7_75t_L g502 ( 
.A(n_451),
.B(n_481),
.C(n_420),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_397),
.Y(n_503)
);

NAND3xp33_ASAP7_75t_L g504 ( 
.A(n_419),
.B(n_273),
.C(n_390),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_472),
.B(n_242),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_462),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_400),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_416),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_408),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_405),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_462),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_R g512 ( 
.A(n_407),
.B(n_380),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_414),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_418),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_418),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_428),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_428),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_472),
.B(n_242),
.Y(n_518)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_462),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_431),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_450),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_411),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_417),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_431),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_424),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_484),
.B(n_342),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_421),
.B(n_202),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_432),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_453),
.B(n_207),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_432),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_434),
.Y(n_531)
);

AND2x6_ASAP7_75t_L g532 ( 
.A(n_394),
.B(n_289),
.Y(n_532)
);

AND3x2_ASAP7_75t_L g533 ( 
.A(n_403),
.B(n_390),
.C(n_206),
.Y(n_533)
);

BUFx10_ASAP7_75t_L g534 ( 
.A(n_429),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_430),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_434),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_438),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_438),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_425),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_422),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_433),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_436),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_460),
.B(n_329),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_443),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_435),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_479),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_479),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_479),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_442),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_486),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_460),
.B(n_296),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_486),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_486),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_394),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_463),
.B(n_296),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_395),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_463),
.B(n_329),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_395),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_398),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_398),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_399),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_399),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_R g563 ( 
.A(n_448),
.B(n_380),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_402),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_452),
.Y(n_565)
);

CKINVDCx16_ASAP7_75t_R g566 ( 
.A(n_457),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_402),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_406),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_406),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_410),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_410),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_455),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_511),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_551),
.B(n_296),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_519),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_519),
.Y(n_576)
);

BUFx8_ASAP7_75t_SL g577 ( 
.A(n_499),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_494),
.B(n_456),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_498),
.B(n_464),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_511),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_532),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_522),
.B(n_440),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_511),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_511),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_494),
.B(n_459),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_511),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_511),
.Y(n_587)
);

AND2x2_ASAP7_75t_SL g588 ( 
.A(n_526),
.B(n_409),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_522),
.B(n_454),
.Y(n_589)
);

AND2x6_ASAP7_75t_L g590 ( 
.A(n_498),
.B(n_317),
.Y(n_590)
);

INVx1_ASAP7_75t_SL g591 ( 
.A(n_512),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_551),
.B(n_317),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_562),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_537),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_537),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_526),
.B(n_461),
.Y(n_596)
);

INVx1_ASAP7_75t_SL g597 ( 
.A(n_563),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_500),
.Y(n_598)
);

INVx4_ASAP7_75t_SL g599 ( 
.A(n_532),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_558),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_502),
.B(n_465),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_502),
.B(n_470),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_537),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_558),
.Y(n_604)
);

OR2x6_ASAP7_75t_L g605 ( 
.A(n_529),
.B(n_474),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_562),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_498),
.B(n_464),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_532),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_562),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_540),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g611 ( 
.A(n_521),
.B(n_411),
.Y(n_611)
);

BUFx4f_ASAP7_75t_L g612 ( 
.A(n_532),
.Y(n_612)
);

OR2x2_ASAP7_75t_L g613 ( 
.A(n_521),
.B(n_415),
.Y(n_613)
);

BUFx2_ASAP7_75t_L g614 ( 
.A(n_540),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_559),
.B(n_471),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_559),
.B(n_476),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_560),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_495),
.B(n_466),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_503),
.B(n_477),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_560),
.B(n_478),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_534),
.B(n_480),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_495),
.B(n_466),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_561),
.B(n_427),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_548),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_495),
.B(n_467),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_561),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_551),
.Y(n_627)
);

BUFx10_ASAP7_75t_L g628 ( 
.A(n_572),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_548),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_562),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_564),
.B(n_329),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_504),
.A2(n_202),
.B1(n_333),
.B2(n_302),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_507),
.B(n_403),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_555),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_564),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_562),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_548),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_567),
.B(n_412),
.Y(n_638)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_497),
.B(n_404),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_534),
.B(n_404),
.Y(n_640)
);

AND2x6_ASAP7_75t_L g641 ( 
.A(n_567),
.B(n_317),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_555),
.B(n_384),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_555),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_568),
.B(n_569),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_497),
.B(n_422),
.Y(n_645)
);

AND2x4_ASAP7_75t_L g646 ( 
.A(n_568),
.B(n_384),
.Y(n_646)
);

INVx4_ASAP7_75t_L g647 ( 
.A(n_562),
.Y(n_647)
);

NAND2xp33_ASAP7_75t_SL g648 ( 
.A(n_505),
.B(n_518),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_569),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_570),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_532),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_570),
.B(n_384),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_496),
.B(n_467),
.Y(n_653)
);

NOR2x1p5_ASAP7_75t_L g654 ( 
.A(n_504),
.B(n_348),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_532),
.B(n_412),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_571),
.Y(n_656)
);

INVx4_ASAP7_75t_L g657 ( 
.A(n_532),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_571),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_SL g659 ( 
.A(n_510),
.B(n_203),
.Y(n_659)
);

AO21x2_ASAP7_75t_L g660 ( 
.A1(n_496),
.A2(n_409),
.B(n_529),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_532),
.A2(n_359),
.B1(n_373),
.B2(n_348),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_571),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_532),
.B(n_413),
.Y(n_663)
);

AND2x6_ASAP7_75t_L g664 ( 
.A(n_554),
.B(n_197),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_554),
.B(n_413),
.Y(n_665)
);

BUFx2_ASAP7_75t_L g666 ( 
.A(n_493),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_513),
.B(n_423),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_554),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_534),
.B(n_324),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_554),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_506),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_543),
.B(n_197),
.Y(n_672)
);

INVx4_ASAP7_75t_L g673 ( 
.A(n_556),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_534),
.B(n_523),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_543),
.B(n_206),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_556),
.Y(n_676)
);

OAI22xp5_ASAP7_75t_L g677 ( 
.A1(n_525),
.A2(n_492),
.B1(n_484),
.B2(n_228),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_535),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_556),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_556),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_SL g681 ( 
.A1(n_527),
.A2(n_302),
.B1(n_349),
.B2(n_333),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_501),
.Y(n_682)
);

INVx6_ASAP7_75t_L g683 ( 
.A(n_506),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_533),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_506),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_506),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_501),
.Y(n_687)
);

AND2x6_ASAP7_75t_L g688 ( 
.A(n_508),
.B(n_217),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_508),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_514),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_557),
.A2(n_359),
.B1(n_373),
.B2(n_348),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_541),
.B(n_469),
.Y(n_692)
);

NAND2xp33_ASAP7_75t_L g693 ( 
.A(n_542),
.B(n_331),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_527),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_514),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_L g696 ( 
.A1(n_557),
.A2(n_373),
.B1(n_389),
.B2(n_359),
.Y(n_696)
);

INVx1_ASAP7_75t_SL g697 ( 
.A(n_509),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_515),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_515),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_516),
.B(n_237),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_516),
.B(n_237),
.Y(n_701)
);

BUFx10_ASAP7_75t_L g702 ( 
.A(n_544),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_517),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_552),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_566),
.B(n_437),
.Y(n_705)
);

BUFx8_ASAP7_75t_SL g706 ( 
.A(n_539),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_517),
.B(n_274),
.Y(n_707)
);

BUFx10_ASAP7_75t_L g708 ( 
.A(n_565),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_566),
.B(n_437),
.Y(n_709)
);

INVx1_ASAP7_75t_SL g710 ( 
.A(n_545),
.Y(n_710)
);

OR2x6_ASAP7_75t_L g711 ( 
.A(n_520),
.B(n_492),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_520),
.B(n_332),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_524),
.B(n_469),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_524),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_528),
.B(n_274),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_552),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_528),
.B(n_338),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_530),
.B(n_485),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_552),
.Y(n_719)
);

INVx6_ASAP7_75t_L g720 ( 
.A(n_552),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_549),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_530),
.B(n_485),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_531),
.B(n_491),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_531),
.A2(n_389),
.B1(n_212),
.B2(n_232),
.Y(n_724)
);

AND2x6_ASAP7_75t_L g725 ( 
.A(n_536),
.B(n_217),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_627),
.B(n_536),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_668),
.Y(n_727)
);

OR2x6_ASAP7_75t_L g728 ( 
.A(n_711),
.B(n_301),
.Y(n_728)
);

BUFx8_ASAP7_75t_L g729 ( 
.A(n_684),
.Y(n_729)
);

NAND2xp33_ASAP7_75t_L g730 ( 
.A(n_590),
.B(n_288),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_588),
.A2(n_229),
.B1(n_267),
.B2(n_227),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_627),
.B(n_538),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_667),
.B(n_458),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_634),
.B(n_538),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_634),
.B(n_227),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_643),
.B(n_229),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_643),
.B(n_267),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_653),
.B(n_268),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_645),
.B(n_225),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_633),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_588),
.A2(n_283),
.B1(n_285),
.B2(n_268),
.Y(n_741)
);

NOR2xp67_ASAP7_75t_L g742 ( 
.A(n_657),
.B(n_546),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_579),
.B(n_283),
.Y(n_743)
);

OR2x6_ASAP7_75t_L g744 ( 
.A(n_711),
.B(n_301),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_588),
.A2(n_648),
.B1(n_666),
.B2(n_601),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_653),
.B(n_285),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_575),
.B(n_299),
.Y(n_747)
);

NAND2xp33_ASAP7_75t_L g748 ( 
.A(n_590),
.B(n_288),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_600),
.Y(n_749)
);

NAND3xp33_ASAP7_75t_SL g750 ( 
.A(n_632),
.B(n_473),
.C(n_468),
.Y(n_750)
);

NOR3xp33_ASAP7_75t_L g751 ( 
.A(n_640),
.B(n_345),
.C(n_225),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_575),
.B(n_299),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_576),
.B(n_307),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_600),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_576),
.B(n_307),
.Y(n_755)
);

BUFx6f_ASAP7_75t_SL g756 ( 
.A(n_628),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_579),
.B(n_328),
.Y(n_757)
);

AND3x1_ASAP7_75t_L g758 ( 
.A(n_632),
.B(n_212),
.C(n_211),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_660),
.A2(n_328),
.B1(n_357),
.B2(n_336),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_604),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_666),
.A2(n_305),
.B1(n_489),
.B2(n_483),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_604),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_660),
.A2(n_336),
.B1(n_357),
.B2(n_379),
.Y(n_763)
);

AND2x2_ASAP7_75t_SL g764 ( 
.A(n_661),
.B(n_379),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_607),
.B(n_487),
.Y(n_765)
);

O2A1O1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_623),
.A2(n_482),
.B(n_447),
.C(n_487),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_607),
.B(n_305),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_605),
.B(n_546),
.Y(n_768)
);

BUFx2_ASAP7_75t_L g769 ( 
.A(n_614),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_605),
.B(n_553),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_605),
.A2(n_475),
.B1(n_374),
.B2(n_356),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_660),
.A2(n_590),
.B1(n_605),
.B2(n_654),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_617),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_605),
.B(n_547),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_617),
.B(n_547),
.Y(n_775)
);

O2A1O1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_700),
.A2(n_482),
.B(n_447),
.C(n_488),
.Y(n_776)
);

NAND2xp33_ASAP7_75t_L g777 ( 
.A(n_590),
.B(n_363),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_582),
.B(n_375),
.Y(n_778)
);

OR2x6_ASAP7_75t_L g779 ( 
.A(n_711),
.B(n_383),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_626),
.B(n_553),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_626),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_635),
.Y(n_782)
);

INVxp67_ASAP7_75t_L g783 ( 
.A(n_589),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_612),
.A2(n_550),
.B(n_490),
.Y(n_784)
);

BUFx3_ASAP7_75t_L g785 ( 
.A(n_577),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_635),
.B(n_550),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_692),
.B(n_391),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_649),
.Y(n_788)
);

NAND2xp33_ASAP7_75t_L g789 ( 
.A(n_590),
.B(n_345),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_649),
.B(n_533),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_706),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_650),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_650),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_687),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_590),
.A2(n_383),
.B1(n_389),
.B2(n_211),
.Y(n_795)
);

NOR2xp67_ASAP7_75t_L g796 ( 
.A(n_657),
.B(n_98),
.Y(n_796)
);

AOI221xp5_ASAP7_75t_L g797 ( 
.A1(n_614),
.A2(n_351),
.B1(n_349),
.B2(n_386),
.C(n_387),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_687),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_690),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_602),
.A2(n_491),
.B1(n_490),
.B2(n_488),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_698),
.B(n_714),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_610),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_690),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_698),
.B(n_439),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_610),
.B(n_221),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_612),
.B(n_230),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_574),
.B(n_439),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_695),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_612),
.B(n_236),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_698),
.B(n_444),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_695),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_699),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_590),
.A2(n_386),
.B1(n_351),
.B2(n_238),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_628),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_714),
.B(n_444),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_699),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_654),
.A2(n_250),
.B1(n_253),
.B2(n_388),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_703),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_615),
.B(n_616),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_672),
.A2(n_250),
.B1(n_253),
.B2(n_388),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_578),
.B(n_239),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_714),
.B(n_644),
.Y(n_822)
);

NOR2xp67_ASAP7_75t_SL g823 ( 
.A(n_581),
.B(n_608),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_672),
.A2(n_245),
.B1(n_243),
.B2(n_387),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_645),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_703),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_620),
.B(n_445),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_672),
.A2(n_245),
.B1(n_243),
.B2(n_385),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_585),
.B(n_240),
.Y(n_829)
);

A2O1A1Ixp33_ASAP7_75t_L g830 ( 
.A1(n_655),
.A2(n_340),
.B(n_234),
.C(n_259),
.Y(n_830)
);

OR2x2_ASAP7_75t_L g831 ( 
.A(n_639),
.B(n_232),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_618),
.B(n_445),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_619),
.B(n_244),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_574),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_591),
.B(n_255),
.Y(n_835)
);

AND2x2_ASAP7_75t_SL g836 ( 
.A(n_672),
.B(n_234),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_668),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_670),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_618),
.B(n_446),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_622),
.B(n_446),
.Y(n_840)
);

BUFx2_ASAP7_75t_L g841 ( 
.A(n_705),
.Y(n_841)
);

NAND2xp33_ASAP7_75t_L g842 ( 
.A(n_664),
.B(n_256),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_622),
.B(n_449),
.Y(n_843)
);

OAI22xp33_ASAP7_75t_L g844 ( 
.A1(n_711),
.A2(n_259),
.B1(n_266),
.B2(n_385),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_597),
.B(n_258),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_670),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_625),
.B(n_449),
.Y(n_847)
);

AND2x2_ASAP7_75t_SL g848 ( 
.A(n_675),
.B(n_266),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_625),
.B(n_260),
.Y(n_849)
);

INVx3_ASAP7_75t_L g850 ( 
.A(n_668),
.Y(n_850)
);

NOR3xp33_ASAP7_75t_L g851 ( 
.A(n_694),
.B(n_270),
.C(n_264),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_675),
.B(n_275),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_679),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_679),
.B(n_271),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_680),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_680),
.Y(n_856)
);

NOR2x1p5_ASAP7_75t_L g857 ( 
.A(n_705),
.B(n_275),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_673),
.B(n_276),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_673),
.B(n_277),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_658),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_657),
.B(n_280),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_596),
.B(n_281),
.Y(n_862)
);

AOI22xp5_ASAP7_75t_L g863 ( 
.A1(n_574),
.A2(n_392),
.B1(n_282),
.B2(n_284),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_574),
.A2(n_293),
.B1(n_300),
.B2(n_378),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_SL g865 ( 
.A(n_598),
.B(n_224),
.Y(n_865)
);

OAI22xp33_ASAP7_75t_L g866 ( 
.A1(n_711),
.A2(n_382),
.B1(n_381),
.B2(n_279),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_592),
.A2(n_303),
.B1(n_304),
.B2(n_377),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_657),
.B(n_308),
.Y(n_868)
);

INVx1_ASAP7_75t_SL g869 ( 
.A(n_709),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_673),
.B(n_309),
.Y(n_870)
);

INVx4_ASAP7_75t_L g871 ( 
.A(n_599),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_592),
.Y(n_872)
);

O2A1O1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_701),
.A2(n_382),
.B(n_381),
.C(n_376),
.Y(n_873)
);

OR2x2_ASAP7_75t_L g874 ( 
.A(n_639),
.B(n_279),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_595),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_709),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_673),
.B(n_310),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_592),
.B(n_314),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_592),
.B(n_315),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_658),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_659),
.B(n_316),
.Y(n_881)
);

INVxp67_ASAP7_75t_L g882 ( 
.A(n_611),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_595),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_595),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_684),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_642),
.B(n_319),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_675),
.B(n_718),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_594),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_594),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_676),
.Y(n_890)
);

NOR2x2_ASAP7_75t_L g891 ( 
.A(n_681),
.B(n_224),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_613),
.B(n_322),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_642),
.B(n_325),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_613),
.B(n_326),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_675),
.B(n_376),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_642),
.B(n_330),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_L g897 ( 
.A1(n_642),
.A2(n_323),
.B1(n_352),
.B2(n_286),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_838),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_769),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_769),
.Y(n_900)
);

AO22x1_ASAP7_75t_L g901 ( 
.A1(n_819),
.A2(n_641),
.B1(n_688),
.B2(n_725),
.Y(n_901)
);

NOR3xp33_ASAP7_75t_SL g902 ( 
.A(n_750),
.B(n_721),
.C(n_677),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_SL g903 ( 
.A1(n_758),
.A2(n_733),
.B1(n_783),
.B2(n_710),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_R g904 ( 
.A(n_785),
.B(n_678),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_745),
.A2(n_693),
.B1(n_674),
.B2(n_621),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_838),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_887),
.B(n_676),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_846),
.Y(n_908)
);

O2A1O1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_767),
.A2(n_707),
.B(n_715),
.C(n_631),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_R g910 ( 
.A(n_785),
.B(n_791),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_802),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_887),
.B(n_676),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_807),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_765),
.B(n_611),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_760),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_871),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_822),
.B(n_646),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_846),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_760),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_871),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_885),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_814),
.Y(n_922)
);

BUFx12f_ASAP7_75t_L g923 ( 
.A(n_729),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_814),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_876),
.Y(n_925)
);

BUFx2_ASAP7_75t_L g926 ( 
.A(n_841),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_853),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_R g928 ( 
.A(n_791),
.B(n_628),
.Y(n_928)
);

OR2x6_ASAP7_75t_L g929 ( 
.A(n_728),
.B(n_581),
.Y(n_929)
);

NAND2xp33_ASAP7_75t_SL g930 ( 
.A(n_823),
.B(n_669),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_SL g931 ( 
.A(n_756),
.B(n_628),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_871),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_853),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_R g934 ( 
.A(n_756),
.B(n_702),
.Y(n_934)
);

NOR2xp67_ASAP7_75t_L g935 ( 
.A(n_740),
.B(n_718),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_855),
.Y(n_936)
);

BUFx12f_ASAP7_75t_L g937 ( 
.A(n_729),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_765),
.B(n_722),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_762),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_833),
.B(n_697),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_882),
.B(n_702),
.Y(n_941)
);

AND2x2_ASAP7_75t_SL g942 ( 
.A(n_731),
.B(n_646),
.Y(n_942)
);

INVx4_ASAP7_75t_L g943 ( 
.A(n_727),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_834),
.A2(n_652),
.B1(n_646),
.B2(n_641),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_836),
.B(n_702),
.Y(n_945)
);

NOR3xp33_ASAP7_75t_SL g946 ( 
.A(n_797),
.B(n_337),
.C(n_334),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_855),
.Y(n_947)
);

NOR2xp67_ASAP7_75t_L g948 ( 
.A(n_845),
.B(n_722),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_762),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_773),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_773),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_856),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_836),
.B(n_723),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_848),
.B(n_702),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_749),
.B(n_646),
.Y(n_955)
);

AND3x1_ASAP7_75t_SL g956 ( 
.A(n_857),
.B(n_292),
.C(n_286),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_834),
.B(n_723),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_R g958 ( 
.A(n_756),
.B(n_708),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_727),
.Y(n_959)
);

BUFx8_ASAP7_75t_L g960 ( 
.A(n_841),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_856),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_872),
.B(n_652),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_794),
.Y(n_963)
);

INVxp67_ASAP7_75t_SL g964 ( 
.A(n_727),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_749),
.B(n_652),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_794),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_848),
.B(n_708),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_837),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_852),
.B(n_708),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_754),
.B(n_781),
.Y(n_970)
);

AO22x1_ASAP7_75t_L g971 ( 
.A1(n_751),
.A2(n_641),
.B1(n_688),
.B2(n_725),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_807),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_807),
.Y(n_973)
);

INVxp67_ASAP7_75t_SL g974 ( 
.A(n_837),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_754),
.B(n_652),
.Y(n_975)
);

INVx6_ASAP7_75t_L g976 ( 
.A(n_728),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_852),
.B(n_708),
.Y(n_977)
);

BUFx3_ASAP7_75t_L g978 ( 
.A(n_729),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_759),
.A2(n_663),
.B(n_665),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_799),
.Y(n_980)
);

INVx5_ASAP7_75t_L g981 ( 
.A(n_837),
.Y(n_981)
);

HB1xp67_ASAP7_75t_L g982 ( 
.A(n_869),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_781),
.B(n_638),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_799),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_808),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_872),
.Y(n_986)
);

NAND2x1p5_ASAP7_75t_L g987 ( 
.A(n_823),
.B(n_581),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_782),
.B(n_713),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_782),
.Y(n_989)
);

AND2x2_ASAP7_75t_SL g990 ( 
.A(n_741),
.B(n_691),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_808),
.Y(n_991)
);

NOR3xp33_ASAP7_75t_SL g992 ( 
.A(n_771),
.B(n_341),
.C(n_339),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_812),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_R g994 ( 
.A(n_842),
.B(n_641),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_788),
.B(n_792),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_788),
.B(n_656),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_812),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_761),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_792),
.B(n_656),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_739),
.B(n_681),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_881),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_816),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_825),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_816),
.Y(n_1004)
);

NAND3xp33_ASAP7_75t_SL g1005 ( 
.A(n_865),
.B(n_696),
.C(n_347),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_793),
.B(n_656),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_739),
.B(n_712),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_857),
.Y(n_1008)
);

BUFx3_ASAP7_75t_L g1009 ( 
.A(n_793),
.Y(n_1009)
);

A2O1A1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_862),
.A2(n_651),
.B(n_608),
.C(n_717),
.Y(n_1010)
);

NOR3xp33_ASAP7_75t_SL g1011 ( 
.A(n_805),
.B(n_350),
.C(n_346),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_826),
.Y(n_1012)
);

INVxp67_ASAP7_75t_L g1013 ( 
.A(n_892),
.Y(n_1013)
);

INVx1_ASAP7_75t_SL g1014 ( 
.A(n_831),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_826),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_888),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_895),
.B(n_608),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_798),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_798),
.B(n_656),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_888),
.Y(n_1020)
);

INVx1_ASAP7_75t_SL g1021 ( 
.A(n_831),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_895),
.B(n_651),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_764),
.A2(n_641),
.B1(n_725),
.B2(n_688),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_728),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_803),
.B(n_662),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_889),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_889),
.Y(n_1027)
);

NAND2xp33_ASAP7_75t_SL g1028 ( 
.A(n_772),
.B(n_682),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_803),
.Y(n_1029)
);

AOI22xp33_ASAP7_75t_L g1030 ( 
.A1(n_764),
.A2(n_641),
.B1(n_725),
.B2(n_688),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_743),
.B(n_651),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_811),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_811),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_874),
.B(n_849),
.Y(n_1034)
);

INVx2_ASAP7_75t_SL g1035 ( 
.A(n_743),
.Y(n_1035)
);

NAND3xp33_ASAP7_75t_SL g1036 ( 
.A(n_813),
.B(n_355),
.C(n_372),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_860),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_818),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_818),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_827),
.B(n_662),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_860),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_880),
.Y(n_1042)
);

INVx4_ASAP7_75t_L g1043 ( 
.A(n_850),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_850),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_874),
.B(n_724),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_738),
.B(n_662),
.Y(n_1046)
);

AND2x4_ASAP7_75t_L g1047 ( 
.A(n_743),
.B(n_599),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_768),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_875),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_875),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_883),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_883),
.Y(n_1052)
);

INVxp67_ASAP7_75t_L g1053 ( 
.A(n_894),
.Y(n_1053)
);

NOR3xp33_ASAP7_75t_SL g1054 ( 
.A(n_835),
.B(n_358),
.C(n_369),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_884),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_746),
.B(n_599),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_726),
.B(n_662),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_R g1058 ( 
.A(n_842),
.B(n_641),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_728),
.Y(n_1059)
);

OR2x2_ASAP7_75t_L g1060 ( 
.A(n_878),
.B(n_879),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_757),
.B(n_599),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_884),
.Y(n_1062)
);

BUFx2_ASAP7_75t_L g1063 ( 
.A(n_744),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_880),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_850),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_890),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_790),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_732),
.B(n_606),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_744),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_890),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_817),
.B(n_764),
.Y(n_1071)
);

NOR2xp67_ASAP7_75t_L g1072 ( 
.A(n_800),
.B(n_580),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_886),
.B(n_599),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_778),
.B(n_593),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_744),
.B(n_606),
.Y(n_1075)
);

INVx4_ASAP7_75t_L g1076 ( 
.A(n_890),
.Y(n_1076)
);

AND2x4_ASAP7_75t_L g1077 ( 
.A(n_744),
.B(n_779),
.Y(n_1077)
);

NOR3xp33_ASAP7_75t_SL g1078 ( 
.A(n_844),
.B(n_354),
.C(n_366),
.Y(n_1078)
);

INVx2_ASAP7_75t_SL g1079 ( 
.A(n_770),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_775),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_780),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_801),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_893),
.B(n_658),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_734),
.B(n_606),
.Y(n_1084)
);

NOR2xp67_ASAP7_75t_L g1085 ( 
.A(n_896),
.B(n_580),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_858),
.B(n_636),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_R g1087 ( 
.A(n_777),
.B(n_606),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_786),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_779),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_774),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_779),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_938),
.B(n_1013),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_938),
.B(n_735),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_1086),
.A2(n_763),
.B(n_804),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1053),
.B(n_736),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_914),
.B(n_737),
.Y(n_1096)
);

INVx2_ASAP7_75t_SL g1097 ( 
.A(n_900),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_916),
.A2(n_742),
.B(n_796),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_914),
.B(n_851),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_SL g1100 ( 
.A1(n_970),
.A2(n_752),
.B(n_747),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_990),
.A2(n_730),
.B(n_748),
.C(n_789),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1081),
.B(n_832),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_SL g1103 ( 
.A1(n_995),
.A2(n_755),
.B(n_753),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_916),
.A2(n_742),
.B(n_796),
.Y(n_1104)
);

HB1xp67_ASAP7_75t_L g1105 ( 
.A(n_899),
.Y(n_1105)
);

A2O1A1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_990),
.A2(n_730),
.B(n_748),
.C(n_789),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_916),
.A2(n_777),
.B(n_647),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_1071),
.A2(n_1028),
.B(n_1007),
.C(n_946),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1081),
.B(n_839),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_1073),
.A2(n_815),
.B(n_810),
.Y(n_1110)
);

NAND3xp33_ASAP7_75t_L g1111 ( 
.A(n_1001),
.B(n_864),
.C(n_863),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_916),
.A2(n_647),
.B(n_593),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_987),
.A2(n_999),
.B(n_996),
.Y(n_1113)
);

AOI21x1_ASAP7_75t_L g1114 ( 
.A1(n_917),
.A2(n_868),
.B(n_861),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_987),
.A2(n_784),
.B(n_630),
.Y(n_1115)
);

AOI211x1_ASAP7_75t_L g1116 ( 
.A1(n_1029),
.A2(n_866),
.B(n_854),
.C(n_829),
.Y(n_1116)
);

AOI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1085),
.A2(n_870),
.B(n_859),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_987),
.A2(n_630),
.B(n_609),
.Y(n_1118)
);

BUFx2_ASAP7_75t_L g1119 ( 
.A(n_900),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1088),
.B(n_840),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_916),
.A2(n_647),
.B(n_593),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1088),
.B(n_843),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_920),
.A2(n_647),
.B(n_593),
.Y(n_1123)
);

NOR4xp25_ASAP7_75t_L g1124 ( 
.A(n_1036),
.B(n_873),
.C(n_776),
.D(n_766),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_942),
.A2(n_795),
.B1(n_877),
.B2(n_779),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1034),
.B(n_847),
.Y(n_1126)
);

AND3x4_ASAP7_75t_L g1127 ( 
.A(n_902),
.B(n_891),
.C(n_867),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_920),
.A2(n_806),
.B(n_809),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_1006),
.A2(n_630),
.B(n_609),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_915),
.Y(n_1130)
);

BUFx2_ASAP7_75t_L g1131 ( 
.A(n_899),
.Y(n_1131)
);

AO31x2_ASAP7_75t_L g1132 ( 
.A1(n_1010),
.A2(n_830),
.A3(n_586),
.B(n_587),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1019),
.A2(n_630),
.B(n_609),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_1031),
.B(n_821),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1034),
.B(n_787),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_1090),
.B(n_636),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1080),
.B(n_897),
.Y(n_1137)
);

AOI21x1_ASAP7_75t_L g1138 ( 
.A1(n_984),
.A2(n_991),
.B(n_985),
.Y(n_1138)
);

CKINVDCx20_ASAP7_75t_R g1139 ( 
.A(n_960),
.Y(n_1139)
);

NOR2x1_ASAP7_75t_SL g1140 ( 
.A(n_920),
.B(n_636),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1025),
.A2(n_609),
.B(n_586),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_942),
.A2(n_905),
.B1(n_1009),
.B2(n_989),
.Y(n_1142)
);

AOI21x1_ASAP7_75t_L g1143 ( 
.A1(n_984),
.A2(n_586),
.B(n_587),
.Y(n_1143)
);

AOI21x1_ASAP7_75t_L g1144 ( 
.A1(n_985),
.A2(n_587),
.B(n_603),
.Y(n_1144)
);

NAND2xp33_ASAP7_75t_SL g1145 ( 
.A(n_920),
.B(n_820),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_898),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1001),
.A2(n_828),
.B1(n_824),
.B2(n_664),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_920),
.A2(n_636),
.B(n_583),
.Y(n_1148)
);

INVx3_ASAP7_75t_SL g1149 ( 
.A(n_1024),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_898),
.Y(n_1150)
);

O2A1O1Ixp5_ASAP7_75t_L g1151 ( 
.A1(n_930),
.A2(n_584),
.B(n_573),
.C(n_603),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1080),
.B(n_682),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_915),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_906),
.A2(n_573),
.B(n_584),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_SL g1155 ( 
.A1(n_932),
.A2(n_636),
.B(n_583),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_935),
.B(n_682),
.Y(n_1156)
);

OAI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1017),
.A2(n_664),
.B(n_584),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_906),
.A2(n_573),
.B(n_584),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_919),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_982),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_932),
.A2(n_636),
.B(n_583),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_1031),
.B(n_573),
.Y(n_1162)
);

OA21x2_ASAP7_75t_L g1163 ( 
.A1(n_979),
.A2(n_624),
.B(n_629),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_932),
.A2(n_981),
.B(n_943),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_948),
.B(n_953),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1017),
.A2(n_664),
.B(n_725),
.Y(n_1166)
);

BUFx12f_ASAP7_75t_L g1167 ( 
.A(n_923),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_953),
.B(n_940),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_988),
.B(n_682),
.Y(n_1169)
);

AO31x2_ASAP7_75t_L g1170 ( 
.A1(n_908),
.A2(n_292),
.A3(n_295),
.B(n_321),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_919),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1014),
.B(n_224),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_939),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_926),
.Y(n_1174)
);

AO32x2_ASAP7_75t_L g1175 ( 
.A1(n_1048),
.A2(n_891),
.A3(n_725),
.B1(n_688),
.B2(n_664),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1048),
.B(n_682),
.Y(n_1176)
);

AOI21x1_ASAP7_75t_L g1177 ( 
.A1(n_991),
.A2(n_624),
.B(n_629),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_939),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_927),
.A2(n_637),
.B(n_685),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_932),
.A2(n_583),
.B(n_689),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_904),
.Y(n_1181)
);

OA22x2_ASAP7_75t_L g1182 ( 
.A1(n_998),
.A2(n_353),
.B1(n_295),
.B2(n_321),
.Y(n_1182)
);

AO31x2_ASAP7_75t_L g1183 ( 
.A1(n_947),
.A2(n_323),
.A3(n_360),
.B(n_368),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_952),
.A2(n_637),
.B(n_716),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_949),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_907),
.A2(n_664),
.B(n_725),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_932),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_952),
.A2(n_637),
.B(n_716),
.Y(n_1188)
);

INVx2_ASAP7_75t_SL g1189 ( 
.A(n_926),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_949),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1090),
.B(n_682),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1079),
.B(n_1060),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_981),
.A2(n_1043),
.B(n_943),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_961),
.A2(n_335),
.A3(n_340),
.B(n_343),
.Y(n_1194)
);

INVx6_ASAP7_75t_L g1195 ( 
.A(n_960),
.Y(n_1195)
);

AOI211x1_ASAP7_75t_L g1196 ( 
.A1(n_1032),
.A2(n_353),
.B(n_335),
.C(n_343),
.Y(n_1196)
);

NOR4xp25_ASAP7_75t_L g1197 ( 
.A(n_909),
.B(n_368),
.C(n_352),
.D(n_360),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_981),
.A2(n_583),
.B(n_689),
.Y(n_1198)
);

BUFx2_ASAP7_75t_L g1199 ( 
.A(n_960),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1071),
.A2(n_370),
.B(n_361),
.C(n_362),
.Y(n_1200)
);

NAND2x1_ASAP7_75t_L g1201 ( 
.A(n_943),
.B(n_683),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_968),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1079),
.B(n_689),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_912),
.A2(n_664),
.B(n_688),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1060),
.B(n_689),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_989),
.B(n_1009),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_925),
.Y(n_1207)
);

OA21x2_ASAP7_75t_L g1208 ( 
.A1(n_961),
.A2(n_671),
.B(n_719),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1021),
.B(n_364),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_SL g1210 ( 
.A1(n_1035),
.A2(n_719),
.B(n_686),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1043),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1043),
.A2(n_1076),
.B(n_1028),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_959),
.A2(n_704),
.B(n_685),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_1090),
.B(n_685),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_968),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_1031),
.B(n_972),
.Y(n_1216)
);

OAI21xp33_ASAP7_75t_L g1217 ( 
.A1(n_998),
.A2(n_941),
.B(n_1045),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1002),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1018),
.A2(n_720),
.B1(n_683),
.B2(n_686),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_1076),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1018),
.B(n_688),
.Y(n_1221)
);

CKINVDCx8_ASAP7_75t_R g1222 ( 
.A(n_1077),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1033),
.B(n_671),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1002),
.A2(n_704),
.A3(n_13),
.B(n_14),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1083),
.A2(n_965),
.B(n_955),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1033),
.B(n_720),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_959),
.A2(n_704),
.B(n_720),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1022),
.A2(n_720),
.B1(n_683),
.B2(n_365),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_969),
.B(n_683),
.Y(n_1229)
);

NOR2x1_ASAP7_75t_L g1230 ( 
.A(n_922),
.B(n_224),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_950),
.Y(n_1231)
);

BUFx12f_ASAP7_75t_L g1232 ( 
.A(n_923),
.Y(n_1232)
);

A2O1A1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1045),
.A2(n_371),
.B(n_13),
.C(n_14),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_959),
.A2(n_181),
.B(n_179),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1076),
.A2(n_176),
.B(n_173),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_975),
.A2(n_171),
.B(n_168),
.Y(n_1236)
);

AO31x2_ASAP7_75t_L g1237 ( 
.A1(n_1004),
.A2(n_10),
.A3(n_16),
.B(n_17),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1083),
.A2(n_142),
.B(n_165),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_969),
.B(n_371),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_950),
.Y(n_1240)
);

OAI21xp33_ASAP7_75t_L g1241 ( 
.A1(n_1000),
.A2(n_1067),
.B(n_1003),
.Y(n_1241)
);

AO31x2_ASAP7_75t_L g1242 ( 
.A1(n_1004),
.A2(n_10),
.A3(n_17),
.B(n_18),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1012),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_951),
.A2(n_164),
.B(n_161),
.Y(n_1244)
);

AOI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1012),
.A2(n_156),
.B(n_153),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_951),
.A2(n_151),
.B(n_149),
.Y(n_1246)
);

CKINVDCx20_ASAP7_75t_R g1247 ( 
.A(n_928),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_963),
.A2(n_147),
.B(n_144),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1046),
.A2(n_143),
.B(n_141),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_977),
.B(n_371),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_963),
.A2(n_138),
.B(n_135),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_SL g1252 ( 
.A(n_1090),
.B(n_977),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1168),
.B(n_967),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1154),
.A2(n_980),
.B(n_966),
.Y(n_1254)
);

BUFx3_ASAP7_75t_L g1255 ( 
.A(n_1174),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1154),
.A2(n_980),
.B(n_966),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1130),
.Y(n_1257)
);

NOR2x1_ASAP7_75t_R g1258 ( 
.A(n_1167),
.B(n_937),
.Y(n_1258)
);

BUFx2_ASAP7_75t_L g1259 ( 
.A(n_1131),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1130),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1153),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1093),
.B(n_967),
.Y(n_1262)
);

OR2x2_ASAP7_75t_L g1263 ( 
.A(n_1165),
.B(n_1000),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_SL g1264 ( 
.A1(n_1238),
.A2(n_997),
.B(n_1038),
.Y(n_1264)
);

INVx2_ASAP7_75t_SL g1265 ( 
.A(n_1174),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1146),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1126),
.B(n_983),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1150),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1158),
.A2(n_1015),
.B(n_993),
.Y(n_1269)
);

OA21x2_ASAP7_75t_L g1270 ( 
.A1(n_1141),
.A2(n_1040),
.B(n_1068),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1158),
.A2(n_1015),
.B(n_993),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1187),
.Y(n_1272)
);

INVx4_ASAP7_75t_L g1273 ( 
.A(n_1187),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1111),
.A2(n_1005),
.B1(n_903),
.B2(n_1008),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1187),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1187),
.Y(n_1276)
);

A2O1A1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1108),
.A2(n_930),
.B(n_992),
.C(n_945),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1217),
.B(n_911),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1129),
.A2(n_1084),
.B(n_1052),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1092),
.B(n_954),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1129),
.A2(n_1055),
.B(n_1052),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_1181),
.Y(n_1282)
);

HB1xp67_ASAP7_75t_L g1283 ( 
.A(n_1105),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1133),
.A2(n_1062),
.B(n_1055),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1108),
.A2(n_1074),
.B(n_1056),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1096),
.B(n_1090),
.Y(n_1286)
);

INVx1_ASAP7_75t_SL g1287 ( 
.A(n_1119),
.Y(n_1287)
);

BUFx4f_ASAP7_75t_L g1288 ( 
.A(n_1216),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1101),
.A2(n_1056),
.B(n_1072),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1133),
.A2(n_1062),
.B(n_1016),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1141),
.A2(n_1027),
.B(n_1020),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1113),
.A2(n_1143),
.B(n_1118),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_1216),
.B(n_1035),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1127),
.A2(n_1063),
.B1(n_1022),
.B2(n_1077),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1207),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_SL g1296 ( 
.A1(n_1142),
.A2(n_997),
.B(n_1039),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1153),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1206),
.A2(n_976),
.B1(n_913),
.B2(n_1022),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1113),
.A2(n_1118),
.B(n_1144),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_1202),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1098),
.A2(n_1104),
.B(n_1155),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1192),
.B(n_957),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1222),
.A2(n_976),
.B1(n_913),
.B2(n_1077),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_1160),
.Y(n_1304)
);

NAND3xp33_ASAP7_75t_L g1305 ( 
.A(n_1200),
.B(n_1054),
.C(n_1011),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1252),
.B(n_918),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1212),
.A2(n_1027),
.B(n_1020),
.Y(n_1307)
);

AO21x1_ASAP7_75t_L g1308 ( 
.A1(n_1125),
.A2(n_1057),
.B(n_933),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1115),
.A2(n_1026),
.B(n_1065),
.Y(n_1309)
);

INVx4_ASAP7_75t_SL g1310 ( 
.A(n_1202),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1189),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1115),
.A2(n_1138),
.B(n_1177),
.Y(n_1312)
);

AO31x2_ASAP7_75t_L g1313 ( 
.A1(n_1101),
.A2(n_1026),
.A3(n_936),
.B(n_1051),
.Y(n_1313)
);

OR2x2_ASAP7_75t_L g1314 ( 
.A(n_1252),
.B(n_1082),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1095),
.B(n_921),
.Y(n_1315)
);

OR2x4_ASAP7_75t_L g1316 ( 
.A(n_1209),
.B(n_973),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1179),
.A2(n_1065),
.B(n_1066),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_1216),
.B(n_1134),
.Y(n_1318)
);

NAND2x1p5_ASAP7_75t_L g1319 ( 
.A(n_1211),
.B(n_1220),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1159),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1102),
.B(n_957),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_R g1322 ( 
.A(n_1181),
.B(n_931),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1179),
.A2(n_1070),
.B(n_1066),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1222),
.A2(n_976),
.B1(n_929),
.B2(n_1091),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1109),
.B(n_957),
.Y(n_1325)
);

CKINVDCx6p67_ASAP7_75t_R g1326 ( 
.A(n_1167),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1159),
.Y(n_1327)
);

INVx8_ASAP7_75t_L g1328 ( 
.A(n_1202),
.Y(n_1328)
);

AO21x2_ASAP7_75t_L g1329 ( 
.A1(n_1106),
.A2(n_1087),
.B(n_994),
.Y(n_1329)
);

AO31x2_ASAP7_75t_L g1330 ( 
.A1(n_1106),
.A2(n_1050),
.A3(n_1049),
.B(n_1070),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1184),
.A2(n_1042),
.B(n_1041),
.Y(n_1331)
);

OAI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1225),
.A2(n_944),
.B(n_1061),
.Y(n_1332)
);

OAI222xp33_ASAP7_75t_L g1333 ( 
.A1(n_1182),
.A2(n_1091),
.B1(n_1089),
.B2(n_1024),
.C1(n_1059),
.C2(n_1063),
.Y(n_1333)
);

BUFx12f_ASAP7_75t_L g1334 ( 
.A(n_1232),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1171),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1218),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1120),
.B(n_1078),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1184),
.A2(n_1188),
.B(n_1213),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1127),
.A2(n_976),
.B1(n_1069),
.B2(n_962),
.Y(n_1339)
);

BUFx12f_ASAP7_75t_L g1340 ( 
.A(n_1232),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1188),
.A2(n_1042),
.B(n_1041),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1122),
.B(n_1082),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1213),
.A2(n_1064),
.B(n_1037),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_1247),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1151),
.A2(n_1064),
.B(n_1037),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_SL g1346 ( 
.A1(n_1195),
.A2(n_958),
.B1(n_934),
.B2(n_1089),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1097),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_SL g1348 ( 
.A1(n_1140),
.A2(n_986),
.B(n_1030),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1243),
.Y(n_1349)
);

INVx4_ASAP7_75t_L g1350 ( 
.A(n_1202),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1110),
.A2(n_1061),
.B(n_974),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1135),
.A2(n_1023),
.B(n_962),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1205),
.B(n_1082),
.Y(n_1353)
);

BUFx2_ASAP7_75t_L g1354 ( 
.A(n_1162),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1099),
.B(n_986),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1134),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1239),
.B(n_1082),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1134),
.B(n_1069),
.Y(n_1358)
);

INVx3_ASAP7_75t_L g1359 ( 
.A(n_1211),
.Y(n_1359)
);

AO31x2_ASAP7_75t_L g1360 ( 
.A1(n_1200),
.A2(n_956),
.A3(n_1082),
.B(n_901),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1171),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1241),
.B(n_1059),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_SL g1363 ( 
.A1(n_1245),
.A2(n_1128),
.B(n_1103),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1173),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1250),
.B(n_922),
.Y(n_1365)
);

AOI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1247),
.A2(n_1075),
.B1(n_962),
.B2(n_924),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1147),
.A2(n_1075),
.B1(n_929),
.B2(n_1047),
.Y(n_1367)
);

AOI21xp33_ASAP7_75t_L g1368 ( 
.A1(n_1209),
.A2(n_1075),
.B(n_929),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_SL g1369 ( 
.A1(n_1100),
.A2(n_929),
.B(n_971),
.Y(n_1369)
);

OAI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1137),
.A2(n_964),
.B(n_1047),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1173),
.Y(n_1371)
);

INVxp67_ASAP7_75t_L g1372 ( 
.A(n_1172),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1110),
.A2(n_1058),
.B(n_901),
.Y(n_1373)
);

INVx6_ASAP7_75t_L g1374 ( 
.A(n_1215),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1107),
.A2(n_1044),
.B(n_968),
.Y(n_1375)
);

AND2x6_ASAP7_75t_SL g1376 ( 
.A(n_1139),
.B(n_937),
.Y(n_1376)
);

CKINVDCx8_ASAP7_75t_R g1377 ( 
.A(n_1199),
.Y(n_1377)
);

AO21x1_ASAP7_75t_L g1378 ( 
.A1(n_1145),
.A2(n_1047),
.B(n_971),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1244),
.A2(n_1044),
.B(n_968),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1162),
.B(n_1178),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1211),
.A2(n_1220),
.B1(n_1221),
.B2(n_1169),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1139),
.Y(n_1382)
);

NAND2x1p5_ASAP7_75t_L g1383 ( 
.A(n_1220),
.B(n_1044),
.Y(n_1383)
);

AO31x2_ASAP7_75t_L g1384 ( 
.A1(n_1233),
.A2(n_1044),
.A3(n_968),
.B(n_22),
.Y(n_1384)
);

NAND2xp33_ASAP7_75t_SL g1385 ( 
.A(n_1215),
.B(n_1044),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1164),
.A2(n_924),
.B(n_978),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1152),
.A2(n_978),
.B1(n_910),
.B2(n_371),
.Y(n_1387)
);

INVx3_ASAP7_75t_L g1388 ( 
.A(n_1215),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1178),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1244),
.A2(n_134),
.B(n_131),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1185),
.B(n_19),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1162),
.Y(n_1392)
);

NAND2xp33_ASAP7_75t_L g1393 ( 
.A(n_1215),
.B(n_130),
.Y(n_1393)
);

BUFx2_ASAP7_75t_L g1394 ( 
.A(n_1185),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_R g1395 ( 
.A1(n_1228),
.A2(n_20),
.B(n_22),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1190),
.Y(n_1396)
);

O2A1O1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1233),
.A2(n_25),
.B(n_28),
.C(n_29),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1190),
.Y(n_1398)
);

AND2x2_ASAP7_75t_SL g1399 ( 
.A(n_1197),
.B(n_29),
.Y(n_1399)
);

OAI221xp5_ASAP7_75t_L g1400 ( 
.A1(n_1230),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.C(n_33),
.Y(n_1400)
);

OAI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1094),
.A2(n_126),
.B(n_116),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1246),
.A2(n_107),
.B(n_101),
.Y(n_1402)
);

OA21x2_ASAP7_75t_L g1403 ( 
.A1(n_1094),
.A2(n_30),
.B(n_32),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1246),
.A2(n_34),
.B(n_37),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1231),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1248),
.A2(n_38),
.B(n_40),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1231),
.Y(n_1407)
);

CKINVDCx6p67_ASAP7_75t_R g1408 ( 
.A(n_1149),
.Y(n_1408)
);

O2A1O1Ixp33_ASAP7_75t_L g1409 ( 
.A1(n_1124),
.A2(n_1156),
.B(n_1229),
.C(n_1191),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1248),
.A2(n_1251),
.B(n_1227),
.Y(n_1410)
);

AO32x2_ASAP7_75t_L g1411 ( 
.A1(n_1196),
.A2(n_40),
.A3(n_41),
.B1(n_44),
.B2(n_47),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1240),
.B(n_44),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1166),
.A2(n_94),
.B(n_49),
.Y(n_1413)
);

AO21x2_ASAP7_75t_L g1414 ( 
.A1(n_1117),
.A2(n_48),
.B(n_49),
.Y(n_1414)
);

INVx3_ASAP7_75t_L g1415 ( 
.A(n_1201),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_SL g1416 ( 
.A1(n_1193),
.A2(n_1249),
.B(n_1235),
.Y(n_1416)
);

A2O1A1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1145),
.A2(n_54),
.B(n_55),
.C(n_57),
.Y(n_1417)
);

AO32x2_ASAP7_75t_L g1418 ( 
.A1(n_1116),
.A2(n_61),
.A3(n_62),
.B1(n_64),
.B2(n_67),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_1149),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1182),
.A2(n_62),
.B1(n_64),
.B2(n_67),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1240),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1253),
.B(n_1170),
.Y(n_1422)
);

CKINVDCx6p67_ASAP7_75t_R g1423 ( 
.A(n_1334),
.Y(n_1423)
);

OAI221xp5_ASAP7_75t_L g1424 ( 
.A1(n_1274),
.A2(n_1195),
.B1(n_1204),
.B2(n_1186),
.C(n_1114),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1267),
.A2(n_1195),
.B1(n_1226),
.B2(n_1203),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1295),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1253),
.B(n_1194),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1319),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1257),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1262),
.B(n_1223),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1262),
.B(n_1194),
.Y(n_1431)
);

NAND3xp33_ASAP7_75t_SL g1432 ( 
.A(n_1397),
.B(n_1176),
.C(n_1191),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1399),
.A2(n_1214),
.B1(n_1163),
.B2(n_1136),
.Y(n_1433)
);

AND2x2_ASAP7_75t_SL g1434 ( 
.A(n_1399),
.B(n_1175),
.Y(n_1434)
);

AOI221xp5_ASAP7_75t_L g1435 ( 
.A1(n_1400),
.A2(n_1210),
.B1(n_1157),
.B2(n_1214),
.C(n_1219),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1372),
.A2(n_1136),
.B1(n_1180),
.B2(n_1198),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1295),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1420),
.A2(n_1163),
.B1(n_1234),
.B2(n_1236),
.Y(n_1438)
);

BUFx3_ASAP7_75t_L g1439 ( 
.A(n_1255),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1263),
.B(n_1183),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1266),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1260),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1301),
.A2(n_1112),
.B(n_1121),
.Y(n_1443)
);

BUFx3_ASAP7_75t_L g1444 ( 
.A(n_1255),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1260),
.Y(n_1445)
);

BUFx4_ASAP7_75t_SL g1446 ( 
.A(n_1376),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1355),
.B(n_1170),
.Y(n_1447)
);

BUFx3_ASAP7_75t_L g1448 ( 
.A(n_1259),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1268),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1261),
.Y(n_1450)
);

INVx3_ASAP7_75t_L g1451 ( 
.A(n_1319),
.Y(n_1451)
);

AOI21xp33_ASAP7_75t_L g1452 ( 
.A1(n_1263),
.A2(n_1163),
.B(n_1236),
.Y(n_1452)
);

INVx6_ASAP7_75t_L g1453 ( 
.A(n_1328),
.Y(n_1453)
);

BUFx3_ASAP7_75t_L g1454 ( 
.A(n_1259),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1261),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1315),
.B(n_1170),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1413),
.A2(n_1234),
.B1(n_1251),
.B2(n_1208),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1297),
.Y(n_1458)
);

AOI221xp5_ASAP7_75t_L g1459 ( 
.A1(n_1417),
.A2(n_1148),
.B1(n_1161),
.B2(n_1123),
.C(n_1194),
.Y(n_1459)
);

INVx5_ASAP7_75t_SL g1460 ( 
.A(n_1408),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_SL g1461 ( 
.A1(n_1362),
.A2(n_1175),
.B1(n_1208),
.B2(n_1227),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1305),
.A2(n_1208),
.B1(n_1237),
.B2(n_1242),
.Y(n_1462)
);

NAND2xp33_ASAP7_75t_SL g1463 ( 
.A(n_1322),
.B(n_1175),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1355),
.B(n_1183),
.Y(n_1464)
);

BUFx2_ASAP7_75t_L g1465 ( 
.A(n_1265),
.Y(n_1465)
);

NAND2xp33_ASAP7_75t_R g1466 ( 
.A(n_1358),
.B(n_1337),
.Y(n_1466)
);

OAI221xp5_ASAP7_75t_L g1467 ( 
.A1(n_1278),
.A2(n_1175),
.B1(n_1170),
.B2(n_1183),
.C(n_1194),
.Y(n_1467)
);

BUFx6f_ASAP7_75t_L g1468 ( 
.A(n_1272),
.Y(n_1468)
);

AND2x4_ASAP7_75t_SL g1469 ( 
.A(n_1408),
.B(n_1183),
.Y(n_1469)
);

BUFx3_ASAP7_75t_L g1470 ( 
.A(n_1265),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1337),
.B(n_1242),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1320),
.Y(n_1472)
);

AND2x4_ASAP7_75t_L g1473 ( 
.A(n_1318),
.B(n_1132),
.Y(n_1473)
);

BUFx8_ASAP7_75t_L g1474 ( 
.A(n_1334),
.Y(n_1474)
);

OAI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1316),
.A2(n_1242),
.B1(n_1237),
.B2(n_1224),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1354),
.B(n_1242),
.Y(n_1476)
);

INVx6_ASAP7_75t_L g1477 ( 
.A(n_1328),
.Y(n_1477)
);

CKINVDCx16_ASAP7_75t_R g1478 ( 
.A(n_1419),
.Y(n_1478)
);

BUFx6f_ASAP7_75t_L g1479 ( 
.A(n_1272),
.Y(n_1479)
);

NAND3xp33_ASAP7_75t_SL g1480 ( 
.A(n_1277),
.B(n_1237),
.C(n_1224),
.Y(n_1480)
);

INVx3_ASAP7_75t_SL g1481 ( 
.A(n_1282),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1283),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1318),
.B(n_1132),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_SL g1484 ( 
.A1(n_1393),
.A2(n_1237),
.B1(n_1224),
.B2(n_1132),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1336),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1308),
.A2(n_1224),
.B1(n_75),
.B2(n_76),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1280),
.B(n_1333),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1316),
.A2(n_1132),
.B1(n_77),
.B2(n_82),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1302),
.B(n_73),
.Y(n_1489)
);

CKINVDCx20_ASAP7_75t_R g1490 ( 
.A(n_1419),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1321),
.B(n_77),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1365),
.B(n_86),
.Y(n_1492)
);

INVx2_ASAP7_75t_SL g1493 ( 
.A(n_1304),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1287),
.B(n_89),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1349),
.Y(n_1495)
);

AOI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1318),
.A2(n_89),
.B1(n_90),
.B2(n_92),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1308),
.A2(n_90),
.B1(n_94),
.B2(n_1325),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1342),
.B(n_1356),
.Y(n_1498)
);

BUFx2_ASAP7_75t_L g1499 ( 
.A(n_1311),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1286),
.B(n_1342),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1344),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1361),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1320),
.Y(n_1503)
);

BUFx12f_ASAP7_75t_L g1504 ( 
.A(n_1340),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1344),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1347),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1366),
.A2(n_1387),
.B1(n_1358),
.B2(n_1316),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1358),
.B(n_1380),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1354),
.B(n_1380),
.Y(n_1509)
);

A2O1A1Ixp33_ASAP7_75t_L g1510 ( 
.A1(n_1285),
.A2(n_1393),
.B(n_1289),
.C(n_1332),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1357),
.B(n_1392),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_1282),
.Y(n_1512)
);

BUFx3_ASAP7_75t_L g1513 ( 
.A(n_1328),
.Y(n_1513)
);

OAI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1288),
.A2(n_1382),
.B1(n_1377),
.B2(n_1395),
.Y(n_1514)
);

AOI21xp33_ASAP7_75t_L g1515 ( 
.A1(n_1409),
.A2(n_1352),
.B(n_1296),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1293),
.B(n_1294),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1368),
.A2(n_1401),
.B1(n_1378),
.B2(n_1414),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1414),
.A2(n_1339),
.B1(n_1306),
.B2(n_1370),
.Y(n_1518)
);

AO22x2_ASAP7_75t_L g1519 ( 
.A1(n_1369),
.A2(n_1363),
.B1(n_1264),
.B2(n_1314),
.Y(n_1519)
);

NAND2x1p5_ASAP7_75t_L g1520 ( 
.A(n_1359),
.B(n_1288),
.Y(n_1520)
);

AND2x4_ASAP7_75t_L g1521 ( 
.A(n_1293),
.B(n_1310),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1327),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1327),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1414),
.A2(n_1306),
.B1(n_1288),
.B2(n_1391),
.Y(n_1524)
);

INVx4_ASAP7_75t_SL g1525 ( 
.A(n_1384),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1335),
.Y(n_1526)
);

INVx4_ASAP7_75t_L g1527 ( 
.A(n_1328),
.Y(n_1527)
);

CKINVDCx8_ASAP7_75t_R g1528 ( 
.A(n_1382),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1364),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1412),
.A2(n_1367),
.B1(n_1324),
.B2(n_1353),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1394),
.B(n_1314),
.Y(n_1531)
);

AO21x2_ASAP7_75t_L g1532 ( 
.A1(n_1363),
.A2(n_1416),
.B(n_1299),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1389),
.Y(n_1533)
);

CKINVDCx8_ASAP7_75t_R g1534 ( 
.A(n_1310),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_1340),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_1326),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1394),
.A2(n_1403),
.B1(n_1303),
.B2(n_1329),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_SL g1538 ( 
.A1(n_1329),
.A2(n_1348),
.B1(n_1298),
.B2(n_1403),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1396),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1407),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1346),
.A2(n_1377),
.B1(n_1386),
.B2(n_1319),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1381),
.A2(n_1383),
.B1(n_1359),
.B2(n_1326),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1383),
.A2(n_1359),
.B1(n_1398),
.B2(n_1405),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1371),
.Y(n_1544)
);

OAI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1273),
.A2(n_1350),
.B1(n_1383),
.B2(n_1421),
.Y(n_1545)
);

BUFx2_ASAP7_75t_L g1546 ( 
.A(n_1388),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1388),
.Y(n_1547)
);

AOI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1329),
.A2(n_1385),
.B1(n_1388),
.B2(n_1374),
.Y(n_1548)
);

OA21x2_ASAP7_75t_L g1549 ( 
.A1(n_1312),
.A2(n_1299),
.B(n_1292),
.Y(n_1549)
);

INVx8_ASAP7_75t_L g1550 ( 
.A(n_1272),
.Y(n_1550)
);

AOI21x1_ASAP7_75t_L g1551 ( 
.A1(n_1410),
.A2(n_1379),
.B(n_1312),
.Y(n_1551)
);

CKINVDCx16_ASAP7_75t_R g1552 ( 
.A(n_1273),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1310),
.B(n_1350),
.Y(n_1553)
);

INVx6_ASAP7_75t_L g1554 ( 
.A(n_1310),
.Y(n_1554)
);

OAI222xp33_ASAP7_75t_L g1555 ( 
.A1(n_1371),
.A2(n_1421),
.B1(n_1405),
.B2(n_1398),
.C1(n_1273),
.C2(n_1350),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1272),
.B(n_1276),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1403),
.A2(n_1406),
.B1(n_1404),
.B2(n_1307),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1345),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1384),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1360),
.B(n_1384),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1345),
.Y(n_1561)
);

CKINVDCx20_ASAP7_75t_R g1562 ( 
.A(n_1374),
.Y(n_1562)
);

BUFx2_ASAP7_75t_L g1563 ( 
.A(n_1374),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1384),
.Y(n_1564)
);

OAI221xp5_ASAP7_75t_L g1565 ( 
.A1(n_1385),
.A2(n_1415),
.B1(n_1270),
.B2(n_1258),
.C(n_1374),
.Y(n_1565)
);

AO21x1_ASAP7_75t_L g1566 ( 
.A1(n_1404),
.A2(n_1406),
.B(n_1307),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1384),
.B(n_1360),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1300),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1360),
.B(n_1313),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1360),
.B(n_1313),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1360),
.B(n_1300),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1272),
.B(n_1276),
.Y(n_1572)
);

NAND3xp33_ASAP7_75t_L g1573 ( 
.A(n_1275),
.B(n_1276),
.C(n_1300),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1313),
.B(n_1330),
.Y(n_1574)
);

INVx2_ASAP7_75t_SL g1575 ( 
.A(n_1275),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1275),
.B(n_1276),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1300),
.Y(n_1577)
);

OAI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1275),
.A2(n_1276),
.B1(n_1300),
.B2(n_1415),
.Y(n_1578)
);

OAI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1275),
.A2(n_1415),
.B1(n_1270),
.B2(n_1313),
.Y(n_1579)
);

AOI221xp5_ASAP7_75t_L g1580 ( 
.A1(n_1418),
.A2(n_1411),
.B1(n_1313),
.B2(n_1330),
.C(n_1402),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1411),
.A2(n_1418),
.B1(n_1270),
.B2(n_1291),
.Y(n_1581)
);

AND2x6_ASAP7_75t_L g1582 ( 
.A(n_1418),
.B(n_1411),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1330),
.Y(n_1583)
);

AOI221xp5_ASAP7_75t_L g1584 ( 
.A1(n_1497),
.A2(n_1492),
.B1(n_1510),
.B2(n_1515),
.C(n_1487),
.Y(n_1584)
);

OAI221xp5_ASAP7_75t_L g1585 ( 
.A1(n_1497),
.A2(n_1411),
.B1(n_1418),
.B2(n_1330),
.C(n_1402),
.Y(n_1585)
);

CKINVDCx6p67_ASAP7_75t_R g1586 ( 
.A(n_1481),
.Y(n_1586)
);

AOI221xp5_ASAP7_75t_L g1587 ( 
.A1(n_1492),
.A2(n_1418),
.B1(n_1411),
.B2(n_1330),
.C(n_1390),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1510),
.A2(n_1373),
.B1(n_1375),
.B2(n_1351),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1509),
.B(n_1309),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1443),
.A2(n_1373),
.B(n_1375),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1500),
.B(n_1430),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1441),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1487),
.A2(n_1291),
.B1(n_1390),
.B2(n_1290),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1449),
.Y(n_1594)
);

AO21x2_ASAP7_75t_L g1595 ( 
.A1(n_1480),
.A2(n_1292),
.B(n_1410),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1496),
.A2(n_1290),
.B1(n_1284),
.B2(n_1281),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1486),
.A2(n_1281),
.B1(n_1284),
.B2(n_1351),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1508),
.B(n_1309),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1486),
.A2(n_1279),
.B1(n_1256),
.B2(n_1269),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1429),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1514),
.A2(n_1279),
.B1(n_1256),
.B2(n_1269),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1491),
.A2(n_1489),
.B1(n_1447),
.B2(n_1464),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1511),
.B(n_1254),
.Y(n_1603)
);

AOI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1507),
.A2(n_1490),
.B1(n_1541),
.B2(n_1530),
.Y(n_1604)
);

CKINVDCx20_ASAP7_75t_R g1605 ( 
.A(n_1490),
.Y(n_1605)
);

AOI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1424),
.A2(n_1379),
.B(n_1338),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1498),
.B(n_1317),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1508),
.B(n_1317),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1434),
.A2(n_1254),
.B1(n_1271),
.B2(n_1331),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1508),
.B(n_1323),
.Y(n_1610)
);

AOI222xp33_ASAP7_75t_L g1611 ( 
.A1(n_1434),
.A2(n_1323),
.B1(n_1271),
.B2(n_1331),
.C1(n_1341),
.C2(n_1343),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1530),
.A2(n_1341),
.B1(n_1343),
.B2(n_1338),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_SL g1613 ( 
.A1(n_1582),
.A2(n_1488),
.B1(n_1516),
.B2(n_1478),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1582),
.A2(n_1471),
.B1(n_1456),
.B2(n_1440),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1582),
.A2(n_1422),
.B1(n_1427),
.B2(n_1431),
.Y(n_1615)
);

INVx3_ASAP7_75t_L g1616 ( 
.A(n_1521),
.Y(n_1616)
);

OR2x2_ASAP7_75t_SL g1617 ( 
.A(n_1446),
.B(n_1494),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1531),
.B(n_1426),
.Y(n_1618)
);

OAI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1466),
.A2(n_1528),
.B1(n_1501),
.B2(n_1505),
.Y(n_1619)
);

AO221x2_ASAP7_75t_L g1620 ( 
.A1(n_1475),
.A2(n_1559),
.B1(n_1564),
.B2(n_1582),
.C(n_1567),
.Y(n_1620)
);

AOI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1466),
.A2(n_1501),
.B1(n_1505),
.B2(n_1423),
.Y(n_1621)
);

BUFx12f_ASAP7_75t_L g1622 ( 
.A(n_1474),
.Y(n_1622)
);

AOI222xp33_ASAP7_75t_SL g1623 ( 
.A1(n_1582),
.A2(n_1482),
.B1(n_1499),
.B2(n_1437),
.C1(n_1506),
.C2(n_1495),
.Y(n_1623)
);

OAI22xp33_ASAP7_75t_L g1624 ( 
.A1(n_1528),
.A2(n_1481),
.B1(n_1493),
.B2(n_1423),
.Y(n_1624)
);

AO21x2_ASAP7_75t_L g1625 ( 
.A1(n_1452),
.A2(n_1566),
.B(n_1551),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1448),
.B(n_1454),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1432),
.A2(n_1518),
.B1(n_1467),
.B2(n_1454),
.Y(n_1627)
);

AOI211xp5_ASAP7_75t_L g1628 ( 
.A1(n_1425),
.A2(n_1542),
.B(n_1565),
.C(n_1436),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1518),
.A2(n_1485),
.B1(n_1504),
.B2(n_1524),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1502),
.Y(n_1630)
);

AOI211xp5_ASAP7_75t_L g1631 ( 
.A1(n_1545),
.A2(n_1580),
.B(n_1459),
.C(n_1535),
.Y(n_1631)
);

OAI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1517),
.A2(n_1435),
.B(n_1524),
.Y(n_1632)
);

AOI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1457),
.A2(n_1555),
.B(n_1537),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1534),
.A2(n_1460),
.B1(n_1536),
.B2(n_1562),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1534),
.A2(n_1460),
.B1(n_1536),
.B2(n_1562),
.Y(n_1635)
);

OAI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1460),
.A2(n_1444),
.B1(n_1439),
.B2(n_1465),
.Y(n_1636)
);

OAI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1535),
.A2(n_1512),
.B1(n_1504),
.B2(n_1444),
.Y(n_1637)
);

AOI221xp5_ASAP7_75t_L g1638 ( 
.A1(n_1517),
.A2(n_1484),
.B1(n_1462),
.B2(n_1463),
.C(n_1519),
.Y(n_1638)
);

AOI221xp5_ASAP7_75t_L g1639 ( 
.A1(n_1462),
.A2(n_1463),
.B1(n_1519),
.B2(n_1581),
.C(n_1438),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1473),
.B(n_1483),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1476),
.B(n_1563),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1547),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1474),
.A2(n_1483),
.B1(n_1473),
.B2(n_1540),
.Y(n_1643)
);

AOI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1512),
.A2(n_1474),
.B1(n_1521),
.B2(n_1473),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1529),
.Y(n_1645)
);

AO21x2_ASAP7_75t_L g1646 ( 
.A1(n_1532),
.A2(n_1579),
.B(n_1558),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1439),
.A2(n_1470),
.B1(n_1548),
.B2(n_1520),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1533),
.B(n_1539),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_SL g1649 ( 
.A1(n_1469),
.A2(n_1554),
.B1(n_1520),
.B2(n_1519),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1537),
.A2(n_1433),
.B1(n_1552),
.B2(n_1554),
.Y(n_1650)
);

OAI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1538),
.A2(n_1438),
.B(n_1543),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1546),
.B(n_1521),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1544),
.A2(n_1560),
.B1(n_1583),
.B2(n_1433),
.Y(n_1653)
);

INVx6_ASAP7_75t_L g1654 ( 
.A(n_1453),
.Y(n_1654)
);

INVxp33_ASAP7_75t_L g1655 ( 
.A(n_1556),
.Y(n_1655)
);

OAI221xp5_ASAP7_75t_L g1656 ( 
.A1(n_1457),
.A2(n_1557),
.B1(n_1461),
.B2(n_1573),
.C(n_1581),
.Y(n_1656)
);

AOI321xp33_ASAP7_75t_L g1657 ( 
.A1(n_1570),
.A2(n_1574),
.A3(n_1569),
.B1(n_1571),
.B2(n_1450),
.C(n_1445),
.Y(n_1657)
);

AOI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1469),
.A2(n_1428),
.B1(n_1451),
.B2(n_1453),
.Y(n_1658)
);

INVx2_ASAP7_75t_SL g1659 ( 
.A(n_1453),
.Y(n_1659)
);

AOI221xp5_ASAP7_75t_L g1660 ( 
.A1(n_1578),
.A2(n_1523),
.B1(n_1442),
.B2(n_1445),
.C(n_1450),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1525),
.A2(n_1472),
.B1(n_1442),
.B2(n_1523),
.Y(n_1661)
);

AOI21xp33_ASAP7_75t_L g1662 ( 
.A1(n_1532),
.A2(n_1577),
.B(n_1568),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1525),
.A2(n_1526),
.B1(n_1503),
.B2(n_1455),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1428),
.B(n_1451),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1525),
.A2(n_1526),
.B1(n_1503),
.B2(n_1455),
.Y(n_1665)
);

INVx4_ASAP7_75t_L g1666 ( 
.A(n_1554),
.Y(n_1666)
);

OAI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1513),
.A2(n_1527),
.B1(n_1477),
.B2(n_1428),
.C(n_1451),
.Y(n_1667)
);

AOI221xp5_ASAP7_75t_L g1668 ( 
.A1(n_1458),
.A2(n_1522),
.B1(n_1558),
.B2(n_1561),
.C(n_1513),
.Y(n_1668)
);

OAI21xp33_ASAP7_75t_L g1669 ( 
.A1(n_1522),
.A2(n_1575),
.B(n_1553),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1477),
.A2(n_1527),
.B1(n_1553),
.B2(n_1576),
.Y(n_1670)
);

OAI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1572),
.A2(n_1576),
.B(n_1549),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1477),
.A2(n_1527),
.B1(n_1479),
.B2(n_1468),
.Y(n_1672)
);

AOI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1468),
.A2(n_1479),
.B1(n_1550),
.B2(n_1549),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_SL g1674 ( 
.A1(n_1468),
.A2(n_1479),
.B(n_1549),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1468),
.B(n_1479),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1550),
.Y(n_1676)
);

OAI221xp5_ASAP7_75t_L g1677 ( 
.A1(n_1550),
.A2(n_1001),
.B1(n_940),
.B2(n_865),
.C(n_733),
.Y(n_1677)
);

OAI221xp5_ASAP7_75t_L g1678 ( 
.A1(n_1497),
.A2(n_1001),
.B1(n_940),
.B2(n_865),
.C(n_733),
.Y(n_1678)
);

BUFx3_ASAP7_75t_L g1679 ( 
.A(n_1439),
.Y(n_1679)
);

AOI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1487),
.A2(n_1001),
.B1(n_733),
.B2(n_940),
.Y(n_1680)
);

AO21x2_ASAP7_75t_L g1681 ( 
.A1(n_1480),
.A2(n_1363),
.B(n_1443),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1497),
.A2(n_1001),
.B1(n_1400),
.B2(n_1399),
.Y(n_1682)
);

OAI221xp5_ASAP7_75t_SL g1683 ( 
.A1(n_1497),
.A2(n_632),
.B1(n_797),
.B2(n_1053),
.C(n_1013),
.Y(n_1683)
);

OAI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1510),
.A2(n_1001),
.B1(n_1127),
.B2(n_1274),
.Y(n_1684)
);

BUFx6f_ASAP7_75t_L g1685 ( 
.A(n_1534),
.Y(n_1685)
);

BUFx3_ASAP7_75t_L g1686 ( 
.A(n_1439),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1509),
.B(n_1508),
.Y(n_1687)
);

OAI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1510),
.A2(n_1001),
.B1(n_1127),
.B2(n_1274),
.Y(n_1688)
);

NAND3xp33_ASAP7_75t_L g1689 ( 
.A(n_1497),
.B(n_833),
.C(n_1001),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1487),
.A2(n_1001),
.B1(n_733),
.B2(n_940),
.Y(n_1690)
);

BUFx6f_ASAP7_75t_L g1691 ( 
.A(n_1534),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1510),
.A2(n_1001),
.B1(n_1127),
.B2(n_1274),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1498),
.B(n_1531),
.Y(n_1693)
);

BUFx6f_ASAP7_75t_L g1694 ( 
.A(n_1534),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1509),
.B(n_1508),
.Y(n_1695)
);

AOI21xp33_ASAP7_75t_L g1696 ( 
.A1(n_1487),
.A2(n_833),
.B(n_1001),
.Y(n_1696)
);

OAI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1510),
.A2(n_1001),
.B1(n_1127),
.B2(n_1274),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1487),
.B(n_1217),
.Y(n_1698)
);

OAI221xp5_ASAP7_75t_L g1699 ( 
.A1(n_1497),
.A2(n_1001),
.B1(n_940),
.B2(n_865),
.C(n_733),
.Y(n_1699)
);

AOI221xp5_ASAP7_75t_L g1700 ( 
.A1(n_1497),
.A2(n_481),
.B1(n_451),
.B2(n_419),
.C(n_420),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1497),
.A2(n_1001),
.B1(n_1400),
.B2(n_1399),
.Y(n_1701)
);

AOI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1497),
.A2(n_1001),
.B1(n_1400),
.B2(n_1399),
.Y(n_1702)
);

AO31x2_ASAP7_75t_L g1703 ( 
.A1(n_1566),
.A2(n_1308),
.A3(n_1579),
.B(n_1510),
.Y(n_1703)
);

BUFx6f_ASAP7_75t_L g1704 ( 
.A(n_1534),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1498),
.B(n_1531),
.Y(n_1705)
);

OAI211xp5_ASAP7_75t_L g1706 ( 
.A1(n_1496),
.A2(n_797),
.B(n_632),
.C(n_1497),
.Y(n_1706)
);

NOR2x1p5_ASAP7_75t_L g1707 ( 
.A(n_1423),
.B(n_1326),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1497),
.A2(n_1001),
.B1(n_1400),
.B2(n_1399),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1500),
.B(n_1430),
.Y(n_1709)
);

OAI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1510),
.A2(n_1001),
.B1(n_1127),
.B2(n_1274),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1497),
.A2(n_1001),
.B1(n_1400),
.B2(n_1399),
.Y(n_1711)
);

OAI21xp33_ASAP7_75t_L g1712 ( 
.A1(n_1497),
.A2(n_833),
.B(n_1001),
.Y(n_1712)
);

AOI221xp5_ASAP7_75t_L g1713 ( 
.A1(n_1497),
.A2(n_481),
.B1(n_451),
.B2(n_419),
.C(n_420),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1620),
.B(n_1615),
.Y(n_1714)
);

OAI211xp5_ASAP7_75t_SL g1715 ( 
.A1(n_1680),
.A2(n_1690),
.B(n_1700),
.C(n_1713),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1600),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1620),
.B(n_1615),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1630),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1600),
.Y(n_1719)
);

INVxp67_ASAP7_75t_SL g1720 ( 
.A(n_1603),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1671),
.B(n_1640),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1645),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1592),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1594),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1591),
.B(n_1709),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1620),
.B(n_1703),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1607),
.Y(n_1727)
);

INVx3_ASAP7_75t_L g1728 ( 
.A(n_1664),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1703),
.B(n_1614),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1598),
.B(n_1608),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1698),
.B(n_1614),
.Y(n_1731)
);

OR2x6_ASAP7_75t_L g1732 ( 
.A(n_1633),
.B(n_1590),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1610),
.B(n_1589),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1698),
.B(n_1602),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1703),
.B(n_1653),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1703),
.B(n_1653),
.Y(n_1736)
);

BUFx3_ASAP7_75t_L g1737 ( 
.A(n_1679),
.Y(n_1737)
);

OAI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1689),
.A2(n_1678),
.B1(n_1699),
.B2(n_1604),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1602),
.B(n_1693),
.Y(n_1739)
);

AO21x2_ASAP7_75t_L g1740 ( 
.A1(n_1632),
.A2(n_1606),
.B(n_1651),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1646),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1646),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1648),
.Y(n_1743)
);

NAND3xp33_ASAP7_75t_L g1744 ( 
.A(n_1696),
.B(n_1584),
.C(n_1683),
.Y(n_1744)
);

BUFx2_ASAP7_75t_L g1745 ( 
.A(n_1642),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1625),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1639),
.B(n_1595),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1625),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1595),
.B(n_1618),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1705),
.B(n_1627),
.Y(n_1750)
);

HB1xp67_ASAP7_75t_L g1751 ( 
.A(n_1681),
.Y(n_1751)
);

AND2x4_ASAP7_75t_SL g1752 ( 
.A(n_1685),
.B(n_1691),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1609),
.B(n_1638),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1609),
.B(n_1681),
.Y(n_1754)
);

OAI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1682),
.A2(n_1711),
.B1(n_1708),
.B2(n_1702),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1611),
.B(n_1593),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1673),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1656),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1585),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1657),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1627),
.B(n_1587),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1588),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1660),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1628),
.B(n_1631),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1674),
.Y(n_1765)
);

OR2x6_ASAP7_75t_L g1766 ( 
.A(n_1650),
.B(n_1647),
.Y(n_1766)
);

AOI21xp5_ASAP7_75t_SL g1767 ( 
.A1(n_1712),
.A2(n_1677),
.B(n_1710),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1662),
.B(n_1593),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1641),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1597),
.B(n_1599),
.Y(n_1770)
);

INVx2_ASAP7_75t_SL g1771 ( 
.A(n_1686),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1629),
.B(n_1663),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1629),
.B(n_1661),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1661),
.Y(n_1774)
);

INVx2_ASAP7_75t_SL g1775 ( 
.A(n_1686),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1597),
.B(n_1599),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1663),
.B(n_1665),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1733),
.B(n_1655),
.Y(n_1778)
);

OAI211xp5_ASAP7_75t_L g1779 ( 
.A1(n_1744),
.A2(n_1706),
.B(n_1708),
.C(n_1711),
.Y(n_1779)
);

AOI221xp5_ASAP7_75t_L g1780 ( 
.A1(n_1715),
.A2(n_1697),
.B1(n_1692),
.B2(n_1688),
.C(n_1684),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1716),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1718),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1725),
.B(n_1626),
.Y(n_1783)
);

AOI33xp33_ASAP7_75t_L g1784 ( 
.A1(n_1758),
.A2(n_1738),
.A3(n_1760),
.B1(n_1701),
.B2(n_1682),
.B3(n_1702),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1718),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1722),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1755),
.A2(n_1701),
.B1(n_1621),
.B2(n_1613),
.Y(n_1787)
);

OAI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1755),
.A2(n_1619),
.B1(n_1643),
.B2(n_1605),
.Y(n_1788)
);

OAI21xp33_ASAP7_75t_L g1789 ( 
.A1(n_1744),
.A2(n_1715),
.B(n_1764),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1764),
.B(n_1624),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1733),
.B(n_1655),
.Y(n_1791)
);

AOI221xp5_ASAP7_75t_L g1792 ( 
.A1(n_1738),
.A2(n_1637),
.B1(n_1636),
.B2(n_1635),
.C(n_1634),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1716),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1722),
.Y(n_1794)
);

AOI22xp33_ASAP7_75t_L g1795 ( 
.A1(n_1760),
.A2(n_1643),
.B1(n_1622),
.B2(n_1586),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1723),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1749),
.B(n_1727),
.Y(n_1797)
);

AOI211xp5_ASAP7_75t_L g1798 ( 
.A1(n_1767),
.A2(n_1667),
.B(n_1669),
.C(n_1644),
.Y(n_1798)
);

INVxp67_ASAP7_75t_L g1799 ( 
.A(n_1745),
.Y(n_1799)
);

AND2x4_ASAP7_75t_L g1800 ( 
.A(n_1721),
.B(n_1658),
.Y(n_1800)
);

AOI222xp33_ASAP7_75t_L g1801 ( 
.A1(n_1734),
.A2(n_1622),
.B1(n_1605),
.B2(n_1707),
.C1(n_1687),
.C2(n_1695),
.Y(n_1801)
);

BUFx6f_ASAP7_75t_L g1802 ( 
.A(n_1737),
.Y(n_1802)
);

BUFx2_ASAP7_75t_L g1803 ( 
.A(n_1721),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1725),
.B(n_1652),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1733),
.B(n_1649),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1723),
.Y(n_1806)
);

BUFx2_ASAP7_75t_L g1807 ( 
.A(n_1721),
.Y(n_1807)
);

AOI221xp5_ASAP7_75t_L g1808 ( 
.A1(n_1758),
.A2(n_1668),
.B1(n_1665),
.B2(n_1676),
.C(n_1596),
.Y(n_1808)
);

OAI33xp33_ASAP7_75t_L g1809 ( 
.A1(n_1734),
.A2(n_1731),
.A3(n_1761),
.B1(n_1759),
.B2(n_1750),
.B3(n_1739),
.Y(n_1809)
);

OAI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1731),
.A2(n_1617),
.B1(n_1670),
.B2(n_1691),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1761),
.A2(n_1616),
.B1(n_1670),
.B2(n_1691),
.Y(n_1811)
);

AND2x4_ASAP7_75t_L g1812 ( 
.A(n_1721),
.B(n_1616),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1739),
.B(n_1654),
.Y(n_1813)
);

OAI211xp5_ASAP7_75t_L g1814 ( 
.A1(n_1753),
.A2(n_1596),
.B(n_1601),
.C(n_1623),
.Y(n_1814)
);

OAI221xp5_ASAP7_75t_L g1815 ( 
.A1(n_1732),
.A2(n_1659),
.B1(n_1672),
.B2(n_1654),
.C(n_1666),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1743),
.B(n_1675),
.Y(n_1816)
);

AO21x2_ASAP7_75t_L g1817 ( 
.A1(n_1746),
.A2(n_1675),
.B(n_1601),
.Y(n_1817)
);

OAI22xp33_ASAP7_75t_L g1818 ( 
.A1(n_1766),
.A2(n_1685),
.B1(n_1691),
.B2(n_1694),
.Y(n_1818)
);

OAI33xp33_ASAP7_75t_L g1819 ( 
.A1(n_1759),
.A2(n_1654),
.A3(n_1666),
.B1(n_1612),
.B2(n_1685),
.B3(n_1694),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1733),
.B(n_1612),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1733),
.B(n_1685),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_R g1822 ( 
.A(n_1737),
.B(n_1694),
.Y(n_1822)
);

NAND2xp33_ASAP7_75t_R g1823 ( 
.A(n_1728),
.B(n_1694),
.Y(n_1823)
);

INVxp67_ASAP7_75t_SL g1824 ( 
.A(n_1720),
.Y(n_1824)
);

AOI221xp5_ASAP7_75t_L g1825 ( 
.A1(n_1753),
.A2(n_1666),
.B1(n_1704),
.B2(n_1714),
.C(n_1717),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1749),
.B(n_1704),
.Y(n_1826)
);

OAI322xp33_ASAP7_75t_L g1827 ( 
.A1(n_1763),
.A2(n_1704),
.A3(n_1750),
.B1(n_1726),
.B2(n_1717),
.C1(n_1714),
.C2(n_1729),
.Y(n_1827)
);

CKINVDCx20_ASAP7_75t_R g1828 ( 
.A(n_1769),
.Y(n_1828)
);

AOI211xp5_ASAP7_75t_SL g1829 ( 
.A1(n_1747),
.A2(n_1704),
.B(n_1753),
.C(n_1756),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1724),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1730),
.B(n_1721),
.Y(n_1831)
);

NAND4xp25_ASAP7_75t_SL g1832 ( 
.A(n_1714),
.B(n_1717),
.C(n_1726),
.D(n_1729),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1719),
.Y(n_1833)
);

OA21x2_ASAP7_75t_L g1834 ( 
.A1(n_1742),
.A2(n_1748),
.B(n_1746),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1740),
.A2(n_1766),
.B1(n_1756),
.B2(n_1770),
.Y(n_1835)
);

AOI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1740),
.A2(n_1766),
.B1(n_1756),
.B2(n_1772),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1803),
.B(n_1726),
.Y(n_1837)
);

OAI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1779),
.A2(n_1763),
.B(n_1766),
.Y(n_1838)
);

AOI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1789),
.A2(n_1740),
.B1(n_1766),
.B2(n_1776),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1782),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1803),
.B(n_1729),
.Y(n_1841)
);

NAND4xp25_ASAP7_75t_L g1842 ( 
.A(n_1784),
.B(n_1735),
.C(n_1736),
.D(n_1747),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1807),
.B(n_1831),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1834),
.Y(n_1844)
);

OR2x6_ASAP7_75t_L g1845 ( 
.A(n_1807),
.B(n_1732),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_SL g1846 ( 
.A(n_1836),
.B(n_1771),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1831),
.B(n_1754),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1797),
.B(n_1749),
.Y(n_1848)
);

BUFx3_ASAP7_75t_L g1849 ( 
.A(n_1802),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1824),
.B(n_1720),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1820),
.B(n_1754),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1797),
.B(n_1727),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1820),
.B(n_1778),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1778),
.B(n_1754),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1782),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1791),
.B(n_1732),
.Y(n_1856)
);

INVx3_ASAP7_75t_L g1857 ( 
.A(n_1834),
.Y(n_1857)
);

INVx1_ASAP7_75t_SL g1858 ( 
.A(n_1826),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1785),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1791),
.B(n_1817),
.Y(n_1860)
);

OR2x2_ASAP7_75t_L g1861 ( 
.A(n_1781),
.B(n_1745),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1834),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1817),
.B(n_1732),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1785),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1834),
.Y(n_1865)
);

BUFx2_ASAP7_75t_L g1866 ( 
.A(n_1812),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1817),
.B(n_1732),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1786),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1786),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1781),
.B(n_1732),
.Y(n_1870)
);

OR2x6_ASAP7_75t_L g1871 ( 
.A(n_1800),
.B(n_1765),
.Y(n_1871)
);

INVxp67_ASAP7_75t_L g1872 ( 
.A(n_1826),
.Y(n_1872)
);

OR2x2_ASAP7_75t_L g1873 ( 
.A(n_1793),
.B(n_1762),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1812),
.B(n_1747),
.Y(n_1874)
);

BUFx3_ASAP7_75t_L g1875 ( 
.A(n_1802),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1812),
.B(n_1736),
.Y(n_1876)
);

OR2x6_ASAP7_75t_L g1877 ( 
.A(n_1800),
.B(n_1765),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1800),
.B(n_1736),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1794),
.B(n_1740),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1793),
.B(n_1762),
.Y(n_1880)
);

AOI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1780),
.A2(n_1766),
.B1(n_1776),
.B2(n_1770),
.Y(n_1881)
);

INVx1_ASAP7_75t_SL g1882 ( 
.A(n_1828),
.Y(n_1882)
);

INVx2_ASAP7_75t_SL g1883 ( 
.A(n_1833),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1794),
.B(n_1735),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1833),
.B(n_1735),
.Y(n_1885)
);

INVx1_ASAP7_75t_SL g1886 ( 
.A(n_1828),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1796),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1884),
.B(n_1796),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1859),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1859),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1884),
.B(n_1806),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1851),
.B(n_1806),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1851),
.B(n_1830),
.Y(n_1893)
);

INVxp67_ASAP7_75t_L g1894 ( 
.A(n_1846),
.Y(n_1894)
);

OR2x2_ASAP7_75t_L g1895 ( 
.A(n_1848),
.B(n_1799),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1851),
.B(n_1830),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1848),
.B(n_1832),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1885),
.B(n_1816),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1859),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1864),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1885),
.B(n_1835),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1860),
.B(n_1805),
.Y(n_1902)
);

NOR3xp33_ASAP7_75t_L g1903 ( 
.A(n_1838),
.B(n_1809),
.C(n_1787),
.Y(n_1903)
);

OAI21xp33_ASAP7_75t_L g1904 ( 
.A1(n_1842),
.A2(n_1881),
.B(n_1838),
.Y(n_1904)
);

INVx2_ASAP7_75t_SL g1905 ( 
.A(n_1849),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1866),
.B(n_1805),
.Y(n_1906)
);

AOI22x1_ASAP7_75t_L g1907 ( 
.A1(n_1882),
.A2(n_1829),
.B1(n_1801),
.B2(n_1768),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1864),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1866),
.B(n_1821),
.Y(n_1909)
);

OAI22xp5_ASAP7_75t_L g1910 ( 
.A1(n_1881),
.A2(n_1814),
.B1(n_1788),
.B2(n_1798),
.Y(n_1910)
);

OR2x6_ASAP7_75t_L g1911 ( 
.A(n_1845),
.B(n_1765),
.Y(n_1911)
);

AND2x4_ASAP7_75t_L g1912 ( 
.A(n_1866),
.B(n_1821),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1844),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1874),
.B(n_1802),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_L g1915 ( 
.A(n_1882),
.B(n_1790),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1844),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1844),
.Y(n_1917)
);

HB1xp67_ASAP7_75t_L g1918 ( 
.A(n_1864),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1874),
.B(n_1802),
.Y(n_1919)
);

AOI222xp33_ASAP7_75t_L g1920 ( 
.A1(n_1839),
.A2(n_1792),
.B1(n_1810),
.B2(n_1825),
.C1(n_1773),
.C2(n_1772),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1844),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1887),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1874),
.B(n_1802),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1887),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1887),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1876),
.B(n_1728),
.Y(n_1926)
);

INVx1_ASAP7_75t_SL g1927 ( 
.A(n_1886),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1840),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1860),
.B(n_1741),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1918),
.Y(n_1930)
);

OAI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1907),
.A2(n_1839),
.B1(n_1910),
.B2(n_1903),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1902),
.B(n_1876),
.Y(n_1932)
);

NOR3xp33_ASAP7_75t_L g1933 ( 
.A(n_1910),
.B(n_1842),
.C(n_1846),
.Y(n_1933)
);

NAND4xp25_ASAP7_75t_L g1934 ( 
.A(n_1903),
.B(n_1863),
.C(n_1867),
.D(n_1795),
.Y(n_1934)
);

OAI211xp5_ASAP7_75t_L g1935 ( 
.A1(n_1904),
.A2(n_1863),
.B(n_1867),
.C(n_1879),
.Y(n_1935)
);

INVxp67_ASAP7_75t_L g1936 ( 
.A(n_1915),
.Y(n_1936)
);

BUFx2_ASAP7_75t_L g1937 ( 
.A(n_1906),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1918),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1904),
.B(n_1878),
.Y(n_1939)
);

O2A1O1Ixp33_ASAP7_75t_L g1940 ( 
.A1(n_1894),
.A2(n_1886),
.B(n_1867),
.C(n_1863),
.Y(n_1940)
);

NAND4xp25_ASAP7_75t_L g1941 ( 
.A(n_1920),
.B(n_1808),
.C(n_1813),
.D(n_1811),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1902),
.B(n_1876),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1902),
.B(n_1853),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1901),
.B(n_1848),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1927),
.B(n_1878),
.Y(n_1945)
);

OR2x2_ASAP7_75t_L g1946 ( 
.A(n_1901),
.B(n_1879),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1928),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1928),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1927),
.B(n_1878),
.Y(n_1949)
);

NAND4xp25_ASAP7_75t_L g1950 ( 
.A(n_1920),
.B(n_1815),
.C(n_1757),
.D(n_1850),
.Y(n_1950)
);

NOR2xp33_ASAP7_75t_L g1951 ( 
.A(n_1894),
.B(n_1872),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1889),
.Y(n_1952)
);

OR2x4_ASAP7_75t_L g1953 ( 
.A(n_1897),
.B(n_1870),
.Y(n_1953)
);

INVx2_ASAP7_75t_SL g1954 ( 
.A(n_1905),
.Y(n_1954)
);

NOR2x1_ASAP7_75t_SL g1955 ( 
.A(n_1897),
.B(n_1871),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1898),
.B(n_1872),
.Y(n_1956)
);

NAND4xp25_ASAP7_75t_L g1957 ( 
.A(n_1906),
.B(n_1757),
.C(n_1850),
.D(n_1870),
.Y(n_1957)
);

AOI221xp5_ASAP7_75t_L g1958 ( 
.A1(n_1892),
.A2(n_1827),
.B1(n_1860),
.B2(n_1819),
.C(n_1858),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1898),
.B(n_1853),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1914),
.B(n_1853),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1914),
.B(n_1847),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1892),
.B(n_1852),
.Y(n_1962)
);

BUFx2_ASAP7_75t_L g1963 ( 
.A(n_1905),
.Y(n_1963)
);

CKINVDCx16_ASAP7_75t_R g1964 ( 
.A(n_1919),
.Y(n_1964)
);

AOI221xp5_ASAP7_75t_L g1965 ( 
.A1(n_1893),
.A2(n_1858),
.B1(n_1783),
.B2(n_1841),
.C(n_1770),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1893),
.B(n_1854),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1896),
.B(n_1854),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1889),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1919),
.B(n_1847),
.Y(n_1969)
);

INVx4_ASAP7_75t_L g1970 ( 
.A(n_1905),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1890),
.Y(n_1971)
);

AND2x4_ASAP7_75t_L g1972 ( 
.A(n_1912),
.B(n_1845),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1896),
.B(n_1854),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1923),
.B(n_1847),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1933),
.B(n_1936),
.Y(n_1975)
);

OAI22xp33_ASAP7_75t_L g1976 ( 
.A1(n_1931),
.A2(n_1907),
.B1(n_1773),
.B2(n_1818),
.Y(n_1976)
);

OAI22xp5_ASAP7_75t_L g1977 ( 
.A1(n_1964),
.A2(n_1937),
.B1(n_1939),
.B2(n_1935),
.Y(n_1977)
);

AND2x4_ASAP7_75t_L g1978 ( 
.A(n_1937),
.B(n_1912),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1947),
.Y(n_1979)
);

AOI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1934),
.A2(n_1845),
.B1(n_1911),
.B2(n_1923),
.Y(n_1980)
);

OAI22xp33_ASAP7_75t_L g1981 ( 
.A1(n_1941),
.A2(n_1950),
.B1(n_1953),
.B2(n_1957),
.Y(n_1981)
);

NAND3x2_ASAP7_75t_L g1982 ( 
.A(n_1946),
.B(n_1870),
.C(n_1929),
.Y(n_1982)
);

INVxp67_ASAP7_75t_L g1983 ( 
.A(n_1951),
.Y(n_1983)
);

OAI31xp33_ASAP7_75t_L g1984 ( 
.A1(n_1940),
.A2(n_1912),
.A3(n_1856),
.B(n_1929),
.Y(n_1984)
);

OAI21xp5_ASAP7_75t_L g1985 ( 
.A1(n_1958),
.A2(n_1911),
.B(n_1856),
.Y(n_1985)
);

AOI21xp5_ASAP7_75t_SL g1986 ( 
.A1(n_1955),
.A2(n_1911),
.B(n_1849),
.Y(n_1986)
);

OAI22xp5_ASAP7_75t_L g1987 ( 
.A1(n_1953),
.A2(n_1845),
.B1(n_1877),
.B2(n_1871),
.Y(n_1987)
);

AOI21xp33_ASAP7_75t_L g1988 ( 
.A1(n_1946),
.A2(n_1954),
.B(n_1944),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1960),
.B(n_1943),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1945),
.B(n_1949),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1948),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1960),
.B(n_1909),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1943),
.B(n_1909),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1965),
.B(n_1912),
.Y(n_1994)
);

AOI21xp5_ASAP7_75t_L g1995 ( 
.A1(n_1955),
.A2(n_1911),
.B(n_1845),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1952),
.Y(n_1996)
);

HB1xp67_ASAP7_75t_L g1997 ( 
.A(n_1963),
.Y(n_1997)
);

AOI22xp5_ASAP7_75t_L g1998 ( 
.A1(n_1972),
.A2(n_1845),
.B1(n_1911),
.B2(n_1871),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1930),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1932),
.B(n_1895),
.Y(n_2000)
);

A2O1A1Ixp33_ASAP7_75t_L g2001 ( 
.A1(n_1944),
.A2(n_1776),
.B(n_1768),
.C(n_1777),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1932),
.B(n_1895),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1942),
.B(n_1926),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1938),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1968),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1968),
.Y(n_2006)
);

OAI22xp33_ASAP7_75t_L g2007 ( 
.A1(n_1953),
.A2(n_1845),
.B1(n_1768),
.B2(n_1777),
.Y(n_2007)
);

INVxp67_ASAP7_75t_L g2008 ( 
.A(n_1963),
.Y(n_2008)
);

OAI22xp33_ASAP7_75t_L g2009 ( 
.A1(n_1974),
.A2(n_1777),
.B1(n_1823),
.B2(n_1871),
.Y(n_2009)
);

OR2x2_ASAP7_75t_L g2010 ( 
.A(n_1959),
.B(n_1888),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1971),
.Y(n_2011)
);

OAI22xp5_ASAP7_75t_L g2012 ( 
.A1(n_1976),
.A2(n_1972),
.B1(n_1942),
.B2(n_1956),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1997),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1997),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1978),
.Y(n_2015)
);

OAI22xp33_ASAP7_75t_L g2016 ( 
.A1(n_1976),
.A2(n_1981),
.B1(n_1975),
.B2(n_1977),
.Y(n_2016)
);

AOI222xp33_ASAP7_75t_L g2017 ( 
.A1(n_1985),
.A2(n_1929),
.B1(n_1972),
.B2(n_1961),
.C1(n_1969),
.C2(n_1967),
.Y(n_2017)
);

AOI22xp5_ASAP7_75t_L g2018 ( 
.A1(n_1981),
.A2(n_1911),
.B1(n_1961),
.B2(n_1969),
.Y(n_2018)
);

AOI21xp33_ASAP7_75t_L g2019 ( 
.A1(n_1983),
.A2(n_1954),
.B(n_1970),
.Y(n_2019)
);

INVx1_ASAP7_75t_SL g2020 ( 
.A(n_1978),
.Y(n_2020)
);

OR2x2_ASAP7_75t_L g2021 ( 
.A(n_2000),
.B(n_1962),
.Y(n_2021)
);

OAI221xp5_ASAP7_75t_L g2022 ( 
.A1(n_1984),
.A2(n_1970),
.B1(n_1962),
.B2(n_1973),
.C(n_1966),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1992),
.B(n_1926),
.Y(n_2023)
);

AOI22xp5_ASAP7_75t_L g2024 ( 
.A1(n_1980),
.A2(n_1871),
.B1(n_1877),
.B2(n_1970),
.Y(n_2024)
);

INVx2_ASAP7_75t_SL g2025 ( 
.A(n_1989),
.Y(n_2025)
);

OA22x2_ASAP7_75t_L g2026 ( 
.A1(n_1986),
.A2(n_1971),
.B1(n_1925),
.B2(n_1924),
.Y(n_2026)
);

INVxp67_ASAP7_75t_SL g2027 ( 
.A(n_2008),
.Y(n_2027)
);

OAI21xp33_ASAP7_75t_SL g2028 ( 
.A1(n_1994),
.A2(n_1843),
.B(n_1891),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1996),
.Y(n_2029)
);

AOI21xp5_ASAP7_75t_SL g2030 ( 
.A1(n_2001),
.A2(n_1875),
.B(n_1849),
.Y(n_2030)
);

O2A1O1Ixp33_ASAP7_75t_L g2031 ( 
.A1(n_2001),
.A2(n_1849),
.B(n_1875),
.C(n_1857),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1979),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1999),
.B(n_1888),
.Y(n_2033)
);

AOI322xp5_ASAP7_75t_L g2034 ( 
.A1(n_2007),
.A2(n_2009),
.A3(n_1988),
.B1(n_1993),
.B2(n_2002),
.C1(n_1990),
.C2(n_2004),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_2005),
.Y(n_2035)
);

OAI221xp5_ASAP7_75t_L g2036 ( 
.A1(n_1998),
.A2(n_1875),
.B1(n_1877),
.B2(n_1871),
.C(n_1891),
.Y(n_2036)
);

INVxp67_ASAP7_75t_L g2037 ( 
.A(n_1991),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_2007),
.B(n_1837),
.Y(n_2038)
);

AOI311xp33_ASAP7_75t_L g2039 ( 
.A1(n_2016),
.A2(n_2009),
.A3(n_1987),
.B(n_1995),
.C(n_2011),
.Y(n_2039)
);

OAI22xp33_ASAP7_75t_L g2040 ( 
.A1(n_2016),
.A2(n_1875),
.B1(n_1877),
.B2(n_1871),
.Y(n_2040)
);

NOR2xp33_ASAP7_75t_SL g2041 ( 
.A(n_2020),
.B(n_2006),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_2027),
.B(n_2003),
.Y(n_2042)
);

CKINVDCx5p33_ASAP7_75t_R g2043 ( 
.A(n_2027),
.Y(n_2043)
);

AND2x4_ASAP7_75t_L g2044 ( 
.A(n_2015),
.B(n_2010),
.Y(n_2044)
);

NAND2xp33_ASAP7_75t_SL g2045 ( 
.A(n_2012),
.B(n_1822),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2013),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_2015),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2014),
.Y(n_2048)
);

AOI222xp33_ASAP7_75t_L g2049 ( 
.A1(n_2028),
.A2(n_1982),
.B1(n_1841),
.B2(n_1837),
.C1(n_1857),
.C2(n_1862),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_2035),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2035),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2029),
.Y(n_2052)
);

NOR2x1p5_ASAP7_75t_SL g2053 ( 
.A(n_2032),
.B(n_1913),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_2025),
.B(n_1837),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_2023),
.B(n_2018),
.Y(n_2055)
);

NOR3xp33_ASAP7_75t_SL g2056 ( 
.A(n_2019),
.B(n_1804),
.C(n_1852),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_2037),
.Y(n_2057)
);

OAI21xp33_ASAP7_75t_L g2058 ( 
.A1(n_2034),
.A2(n_1877),
.B(n_1856),
.Y(n_2058)
);

NOR2xp33_ASAP7_75t_L g2059 ( 
.A(n_2037),
.B(n_1890),
.Y(n_2059)
);

NOR4xp25_ASAP7_75t_L g2060 ( 
.A(n_2039),
.B(n_2031),
.C(n_2022),
.D(n_2038),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_SL g2061 ( 
.A(n_2043),
.B(n_2026),
.Y(n_2061)
);

INVxp67_ASAP7_75t_SL g2062 ( 
.A(n_2041),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_2047),
.Y(n_2063)
);

AOI222xp33_ASAP7_75t_L g2064 ( 
.A1(n_2058),
.A2(n_2045),
.B1(n_2040),
.B2(n_2057),
.C1(n_2042),
.C2(n_2046),
.Y(n_2064)
);

AOI21xp5_ASAP7_75t_L g2065 ( 
.A1(n_2045),
.A2(n_2030),
.B(n_2026),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_2047),
.Y(n_2066)
);

OR2x2_ASAP7_75t_L g2067 ( 
.A(n_2044),
.B(n_2021),
.Y(n_2067)
);

NOR3xp33_ASAP7_75t_L g2068 ( 
.A(n_2048),
.B(n_2036),
.C(n_2024),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2050),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2051),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_2055),
.B(n_2017),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_2067),
.Y(n_2072)
);

O2A1O1Ixp33_ASAP7_75t_L g2073 ( 
.A1(n_2061),
.A2(n_2040),
.B(n_2052),
.C(n_2056),
.Y(n_2073)
);

INVxp67_ASAP7_75t_L g2074 ( 
.A(n_2062),
.Y(n_2074)
);

AOI221xp5_ASAP7_75t_L g2075 ( 
.A1(n_2060),
.A2(n_2044),
.B1(n_2059),
.B2(n_2054),
.C(n_2033),
.Y(n_2075)
);

AOI21xp5_ASAP7_75t_L g2076 ( 
.A1(n_2061),
.A2(n_2065),
.B(n_2071),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2063),
.Y(n_2077)
);

AOI322xp5_ASAP7_75t_L g2078 ( 
.A1(n_2071),
.A2(n_2059),
.A3(n_2044),
.B1(n_2049),
.B2(n_1841),
.C1(n_2053),
.C2(n_1857),
.Y(n_2078)
);

NOR4xp25_ASAP7_75t_L g2079 ( 
.A(n_2066),
.B(n_1917),
.C(n_1913),
.D(n_1916),
.Y(n_2079)
);

AOI22xp33_ASAP7_75t_L g2080 ( 
.A1(n_2068),
.A2(n_1877),
.B1(n_1774),
.B2(n_1751),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2064),
.B(n_1899),
.Y(n_2081)
);

OAI221xp5_ASAP7_75t_SL g2082 ( 
.A1(n_2070),
.A2(n_1877),
.B1(n_1913),
.B2(n_1921),
.C(n_1917),
.Y(n_2082)
);

INVxp67_ASAP7_75t_L g2083 ( 
.A(n_2072),
.Y(n_2083)
);

NAND3xp33_ASAP7_75t_L g2084 ( 
.A(n_2076),
.B(n_2063),
.C(n_2069),
.Y(n_2084)
);

INVx5_ASAP7_75t_L g2085 ( 
.A(n_2074),
.Y(n_2085)
);

OAI321xp33_ASAP7_75t_L g2086 ( 
.A1(n_2081),
.A2(n_1771),
.A3(n_1775),
.B1(n_1916),
.B2(n_1917),
.C(n_1921),
.Y(n_2086)
);

NOR2xp67_ASAP7_75t_L g2087 ( 
.A(n_2077),
.B(n_1899),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2075),
.Y(n_2088)
);

OAI211xp5_ASAP7_75t_L g2089 ( 
.A1(n_2088),
.A2(n_2073),
.B(n_2078),
.C(n_2080),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_2085),
.B(n_2073),
.Y(n_2090)
);

OAI22xp5_ASAP7_75t_L g2091 ( 
.A1(n_2083),
.A2(n_2085),
.B1(n_2084),
.B2(n_2082),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_2087),
.B(n_2079),
.Y(n_2092)
);

HB1xp67_ASAP7_75t_L g2093 ( 
.A(n_2086),
.Y(n_2093)
);

NOR3xp33_ASAP7_75t_L g2094 ( 
.A(n_2088),
.B(n_1916),
.C(n_1921),
.Y(n_2094)
);

AOI332xp33_ASAP7_75t_L g2095 ( 
.A1(n_2088),
.A2(n_1925),
.A3(n_1900),
.B1(n_1908),
.B2(n_1922),
.B3(n_1924),
.C1(n_1857),
.C2(n_1862),
.Y(n_2095)
);

OAI221xp5_ASAP7_75t_SL g2096 ( 
.A1(n_2089),
.A2(n_1861),
.B1(n_1857),
.B2(n_1843),
.C(n_1862),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_2090),
.Y(n_2097)
);

NOR2x1_ASAP7_75t_L g2098 ( 
.A(n_2091),
.B(n_1900),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_2093),
.B(n_1908),
.Y(n_2099)
);

OAI222xp33_ASAP7_75t_L g2100 ( 
.A1(n_2092),
.A2(n_1861),
.B1(n_1922),
.B2(n_1862),
.C1(n_1865),
.C2(n_1775),
.Y(n_2100)
);

XNOR2xp5_ASAP7_75t_L g2101 ( 
.A(n_2094),
.B(n_1752),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2097),
.B(n_2095),
.Y(n_2102)
);

NOR2xp33_ASAP7_75t_L g2103 ( 
.A(n_2099),
.B(n_1861),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2098),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_SL g2105 ( 
.A(n_2101),
.B(n_2096),
.Y(n_2105)
);

AOI21xp5_ASAP7_75t_L g2106 ( 
.A1(n_2105),
.A2(n_2100),
.B(n_1865),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_SL g2107 ( 
.A(n_2106),
.B(n_2104),
.Y(n_2107)
);

NOR3xp33_ASAP7_75t_L g2108 ( 
.A(n_2107),
.B(n_2102),
.C(n_2103),
.Y(n_2108)
);

INVx1_ASAP7_75t_SL g2109 ( 
.A(n_2107),
.Y(n_2109)
);

OAI21xp5_ASAP7_75t_SL g2110 ( 
.A1(n_2109),
.A2(n_1752),
.B(n_1843),
.Y(n_2110)
);

AOI221xp5_ASAP7_75t_L g2111 ( 
.A1(n_2108),
.A2(n_1865),
.B1(n_1883),
.B2(n_1869),
.C(n_1855),
.Y(n_2111)
);

AOI21xp5_ASAP7_75t_L g2112 ( 
.A1(n_2110),
.A2(n_1865),
.B(n_1883),
.Y(n_2112)
);

OAI21x1_ASAP7_75t_SL g2113 ( 
.A1(n_2111),
.A2(n_1771),
.B(n_1775),
.Y(n_2113)
);

INVxp67_ASAP7_75t_L g2114 ( 
.A(n_2113),
.Y(n_2114)
);

OAI221xp5_ASAP7_75t_R g2115 ( 
.A1(n_2114),
.A2(n_2112),
.B1(n_1883),
.B2(n_1873),
.C(n_1880),
.Y(n_2115)
);

AOI211xp5_ASAP7_75t_L g2116 ( 
.A1(n_2115),
.A2(n_1880),
.B(n_1873),
.C(n_1868),
.Y(n_2116)
);


endmodule