module fake_jpeg_20179_n_205 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_205);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_6),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_11),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_17),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_14),
.B1(n_17),
.B2(n_13),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_32),
.B1(n_24),
.B2(n_30),
.Y(n_44)
);

HAxp5_ASAP7_75t_SL g39 ( 
.A(n_26),
.B(n_20),
.CON(n_39),
.SN(n_39)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_18),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_17),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_52),
.B1(n_57),
.B2(n_59),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_27),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_45),
.B(n_46),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_28),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_54),
.C(n_35),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_20),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_20),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_25),
.B1(n_31),
.B2(n_14),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_55),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_25),
.C(n_31),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_37),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_30),
.B1(n_31),
.B2(n_29),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_34),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_35),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_30),
.B1(n_29),
.B2(n_28),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_29),
.B1(n_28),
.B2(n_18),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_43),
.B1(n_37),
.B2(n_34),
.Y(n_66)
);

NOR2x1p5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_35),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_68),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_64),
.A2(n_76),
.B(n_47),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_71),
.B1(n_72),
.B2(n_44),
.Y(n_86)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_74),
.Y(n_80)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_43),
.B1(n_37),
.B2(n_34),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_43),
.B1(n_37),
.B2(n_33),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_60),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_78),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_37),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_71),
.Y(n_90)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_43),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_65),
.B(n_48),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_81),
.B(n_87),
.Y(n_102)
);

AO21x1_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_64),
.B(n_76),
.Y(n_100)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_89),
.B1(n_93),
.B2(n_70),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_79),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_88),
.A2(n_90),
.B(n_62),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_47),
.B1(n_59),
.B2(n_46),
.Y(n_89)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_92),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_46),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_45),
.B1(n_50),
.B2(n_33),
.Y(n_93)
);

AND2x6_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_41),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_93),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_35),
.C(n_41),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_18),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_96),
.Y(n_105)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_106),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_64),
.B1(n_69),
.B2(n_72),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_101),
.A2(n_16),
.B1(n_13),
.B2(n_15),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_103),
.A2(n_9),
.B(n_11),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_104),
.B(n_110),
.Y(n_132)
);

OA21x2_ASAP7_75t_L g107 ( 
.A1(n_83),
.A2(n_70),
.B(n_67),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_116),
.Y(n_120)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_108),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_61),
.B1(n_21),
.B2(n_16),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_111),
.B(n_113),
.Y(n_137)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

AOI221xp5_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_88),
.B1(n_97),
.B2(n_89),
.C(n_90),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_61),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_115),
.B(n_117),
.Y(n_119)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_81),
.B(n_22),
.Y(n_117)
);

AOI322xp5_ASAP7_75t_L g146 ( 
.A1(n_122),
.A2(n_123),
.A3(n_109),
.B1(n_99),
.B2(n_100),
.C1(n_104),
.C2(n_8),
.Y(n_146)
);

AOI322xp5_ASAP7_75t_L g123 ( 
.A1(n_112),
.A2(n_97),
.A3(n_92),
.B1(n_86),
.B2(n_95),
.C1(n_21),
.C2(n_16),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_117),
.B(n_15),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_124),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_130),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_21),
.Y(n_126)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_127),
.A2(n_133),
.B1(n_136),
.B2(n_12),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_L g128 ( 
.A1(n_102),
.A2(n_13),
.B(n_15),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_113),
.A2(n_116),
.B1(n_111),
.B2(n_98),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_129),
.A2(n_138),
.B1(n_105),
.B2(n_98),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_102),
.B(n_7),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_107),
.A2(n_22),
.B1(n_12),
.B2(n_2),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_101),
.A2(n_22),
.B1(n_12),
.B2(n_2),
.Y(n_136)
);

MAJx2_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_7),
.C(n_11),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_118),
.C(n_106),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_141),
.C(n_148),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_140),
.B(n_151),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_118),
.C(n_107),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_142),
.B(n_136),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_104),
.B1(n_100),
.B2(n_108),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_144),
.A2(n_154),
.B1(n_127),
.B2(n_126),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_153),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_129),
.C(n_120),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_137),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_152),
.Y(n_159)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_144),
.A2(n_131),
.B(n_135),
.Y(n_156)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_158),
.A2(n_5),
.B1(n_9),
.B2(n_8),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_125),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_145),
.C(n_154),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_150),
.A2(n_135),
.B(n_126),
.Y(n_164)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_164),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_139),
.A2(n_130),
.B1(n_119),
.B2(n_138),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_165),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

INVx11_ASAP7_75t_L g170 ( 
.A(n_166),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_161),
.A2(n_141),
.B(n_142),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_163),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_157),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_155),
.A2(n_145),
.B1(n_143),
.B2(n_140),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_155),
.A2(n_5),
.B1(n_9),
.B2(n_8),
.Y(n_173)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_174),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_169),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_182),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_175),
.B(n_166),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_181),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_162),
.Y(n_180)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_180),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_160),
.C(n_159),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_159),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_176),
.A2(n_5),
.B(n_10),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_185),
.C(n_174),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_167),
.A2(n_0),
.B(n_1),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_189),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_188),
.B(n_190),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_172),
.C(n_173),
.Y(n_189)
);

OR2x6_ASAP7_75t_SL g190 ( 
.A(n_178),
.B(n_170),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_183),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_195),
.Y(n_199)
);

NOR2xp67_ASAP7_75t_L g194 ( 
.A(n_190),
.B(n_0),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_196),
.C(n_187),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_192),
.B(n_1),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_3),
.C(n_4),
.Y(n_196)
);

BUFx24_ASAP7_75t_SL g203 ( 
.A(n_200),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_3),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_197),
.Y(n_202)
);

AO21x1_ASAP7_75t_L g204 ( 
.A1(n_202),
.A2(n_199),
.B(n_4),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_203),
.Y(n_205)
);


endmodule