module fake_netlist_1_46_n_21 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_21);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_21;
wire n_20;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
INVx2_ASAP7_75t_L g9 ( .A(n_1), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_1), .Y(n_10) );
INVx2_ASAP7_75t_SL g11 ( .A(n_3), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
AOI22xp5_ASAP7_75t_L g13 ( .A1(n_8), .A2(n_0), .B1(n_6), .B2(n_5), .Y(n_13) );
OAI21x1_ASAP7_75t_L g14 ( .A1(n_12), .A2(n_2), .B(n_7), .Y(n_14) );
INVx3_ASAP7_75t_SL g15 ( .A(n_11), .Y(n_15) );
AND2x4_ASAP7_75t_L g16 ( .A(n_14), .B(n_10), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_16), .B(n_15), .Y(n_17) );
NOR2xp33_ASAP7_75t_L g18 ( .A(n_17), .B(n_15), .Y(n_18) );
AND3x2_ASAP7_75t_L g19 ( .A(n_18), .B(n_10), .C(n_9), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_20), .B(n_13), .Y(n_21) );
endmodule