module fake_ariane_1194_n_2932 (n_295, n_356, n_556, n_170, n_190, n_698, n_695, n_160, n_64, n_180, n_730, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_830, n_176, n_691, n_34, n_404, n_172, n_678, n_651, n_347, n_423, n_183, n_469, n_479, n_726, n_603, n_373, n_299, n_836, n_541, n_499, n_789, n_788, n_12, n_771, n_564, n_133, n_610, n_66, n_205, n_752, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_760, n_20, n_690, n_416, n_283, n_50, n_187, n_525, n_806, n_367, n_713, n_649, n_598, n_345, n_374, n_318, n_817, n_103, n_244, n_643, n_679, n_226, n_781, n_220, n_261, n_682, n_36, n_663, n_370, n_706, n_189, n_717, n_819, n_72, n_286, n_443, n_586, n_57, n_686, n_605, n_776, n_424, n_528, n_584, n_387, n_406, n_826, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_756, n_346, n_214, n_764, n_348, n_552, n_2, n_462, n_607, n_670, n_32, n_410, n_379, n_445, n_515, n_807, n_138, n_162, n_765, n_264, n_737, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_766, n_372, n_377, n_15, n_396, n_802, n_631, n_23, n_399, n_554, n_520, n_87, n_714, n_279, n_702, n_207, n_790, n_363, n_720, n_354, n_41, n_813, n_140, n_725, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_801, n_202, n_145, n_193, n_733, n_761, n_818, n_500, n_665, n_59, n_336, n_731, n_754, n_779, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_829, n_8, n_668, n_339, n_738, n_758, n_833, n_672, n_487, n_740, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_784, n_269, n_597, n_816, n_75, n_158, n_69, n_259, n_835, n_95, n_808, n_446, n_553, n_143, n_753, n_566, n_814, n_578, n_701, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_822, n_344, n_381, n_795, n_426, n_433, n_481, n_600, n_721, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_770, n_218, n_821, n_79, n_839, n_3, n_271, n_465, n_486, n_507, n_759, n_247, n_569, n_567, n_825, n_732, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_787, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_703, n_748, n_786, n_510, n_831, n_256, n_326, n_681, n_778, n_227, n_48, n_188, n_323, n_550, n_635, n_707, n_330, n_400, n_689, n_694, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_699, n_727, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_823, n_620, n_228, n_325, n_276, n_93, n_688, n_636, n_427, n_108, n_587, n_497, n_693, n_303, n_671, n_442, n_777, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_729, n_661, n_488, n_775, n_667, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_684, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_728, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_715, n_579, n_459, n_685, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_838, n_237, n_780, n_175, n_711, n_453, n_734, n_74, n_491, n_810, n_19, n_40, n_181, n_723, n_616, n_617, n_658, n_630, n_705, n_570, n_53, n_260, n_362, n_543, n_310, n_709, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_809, n_461, n_209, n_262, n_490, n_743, n_17, n_225, n_235, n_660, n_464, n_735, n_575, n_546, n_297, n_662, n_641, n_503, n_700, n_290, n_527, n_46, n_741, n_747, n_772, n_84, n_371, n_199, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_708, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_680, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_755, n_710, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_652, n_451, n_613, n_745, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_716, n_102, n_742, n_182, n_696, n_674, n_482, n_316, n_196, n_125, n_798, n_769, n_820, n_43, n_577, n_407, n_774, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_832, n_55, n_535, n_231, n_366, n_744, n_762, n_656, n_555, n_234, n_492, n_574, n_804, n_280, n_215, n_252, n_629, n_664, n_161, n_454, n_298, n_532, n_68, n_415, n_794, n_763, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_692, n_5, n_599, n_768, n_514, n_418, n_537, n_223, n_403, n_25, n_750, n_834, n_83, n_389, n_800, n_657, n_513, n_837, n_288, n_179, n_812, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_659, n_67, n_509, n_583, n_724, n_306, n_666, n_313, n_92, n_430, n_626, n_493, n_722, n_203, n_378, n_436, n_150, n_98, n_757, n_375, n_113, n_114, n_33, n_324, n_585, n_669, n_785, n_827, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_697, n_472, n_296, n_265, n_746, n_208, n_456, n_156, n_292, n_793, n_174, n_275, n_100, n_704, n_132, n_147, n_204, n_751, n_615, n_521, n_51, n_496, n_739, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_792, n_824, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_719, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_773, n_165, n_144, n_317, n_101, n_243, n_803, n_134, n_329, n_718, n_185, n_340, n_749, n_289, n_9, n_112, n_45, n_542, n_548, n_815, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_782, n_425, n_431, n_811, n_508, n_624, n_118, n_121, n_791, n_618, n_411, n_484, n_712, n_353, n_22, n_736, n_767, n_241, n_29, n_357, n_412, n_687, n_447, n_191, n_382, n_797, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_828, n_595, n_322, n_251, n_506, n_602, n_799, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_796, n_805, n_127, n_531, n_783, n_675, n_2932);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_698;
input n_695;
input n_160;
input n_64;
input n_180;
input n_730;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_830;
input n_176;
input n_691;
input n_34;
input n_404;
input n_172;
input n_678;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_726;
input n_603;
input n_373;
input n_299;
input n_836;
input n_541;
input n_499;
input n_789;
input n_788;
input n_12;
input n_771;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_752;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_760;
input n_20;
input n_690;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_806;
input n_367;
input n_713;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_817;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_781;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_706;
input n_189;
input n_717;
input n_819;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_686;
input n_605;
input n_776;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_826;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_756;
input n_346;
input n_214;
input n_764;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_807;
input n_138;
input n_162;
input n_765;
input n_264;
input n_737;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_766;
input n_372;
input n_377;
input n_15;
input n_396;
input n_802;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_714;
input n_279;
input n_702;
input n_207;
input n_790;
input n_363;
input n_720;
input n_354;
input n_41;
input n_813;
input n_140;
input n_725;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_801;
input n_202;
input n_145;
input n_193;
input n_733;
input n_761;
input n_818;
input n_500;
input n_665;
input n_59;
input n_336;
input n_731;
input n_754;
input n_779;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_829;
input n_8;
input n_668;
input n_339;
input n_738;
input n_758;
input n_833;
input n_672;
input n_487;
input n_740;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_784;
input n_269;
input n_597;
input n_816;
input n_75;
input n_158;
input n_69;
input n_259;
input n_835;
input n_95;
input n_808;
input n_446;
input n_553;
input n_143;
input n_753;
input n_566;
input n_814;
input n_578;
input n_701;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_822;
input n_344;
input n_381;
input n_795;
input n_426;
input n_433;
input n_481;
input n_600;
input n_721;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_770;
input n_218;
input n_821;
input n_79;
input n_839;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_759;
input n_247;
input n_569;
input n_567;
input n_825;
input n_732;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_787;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_703;
input n_748;
input n_786;
input n_510;
input n_831;
input n_256;
input n_326;
input n_681;
input n_778;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_707;
input n_330;
input n_400;
input n_689;
input n_694;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_699;
input n_727;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_823;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_693;
input n_303;
input n_671;
input n_442;
input n_777;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_729;
input n_661;
input n_488;
input n_775;
input n_667;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_728;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_715;
input n_579;
input n_459;
input n_685;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_838;
input n_237;
input n_780;
input n_175;
input n_711;
input n_453;
input n_734;
input n_74;
input n_491;
input n_810;
input n_19;
input n_40;
input n_181;
input n_723;
input n_616;
input n_617;
input n_658;
input n_630;
input n_705;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_709;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_809;
input n_461;
input n_209;
input n_262;
input n_490;
input n_743;
input n_17;
input n_225;
input n_235;
input n_660;
input n_464;
input n_735;
input n_575;
input n_546;
input n_297;
input n_662;
input n_641;
input n_503;
input n_700;
input n_290;
input n_527;
input n_46;
input n_741;
input n_747;
input n_772;
input n_84;
input n_371;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_708;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_755;
input n_710;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_652;
input n_451;
input n_613;
input n_745;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_716;
input n_102;
input n_742;
input n_182;
input n_696;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_798;
input n_769;
input n_820;
input n_43;
input n_577;
input n_407;
input n_774;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_832;
input n_55;
input n_535;
input n_231;
input n_366;
input n_744;
input n_762;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_804;
input n_280;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_794;
input n_763;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_692;
input n_5;
input n_599;
input n_768;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_750;
input n_834;
input n_83;
input n_389;
input n_800;
input n_657;
input n_513;
input n_837;
input n_288;
input n_179;
input n_812;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_659;
input n_67;
input n_509;
input n_583;
input n_724;
input n_306;
input n_666;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_722;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_757;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_669;
input n_785;
input n_827;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_697;
input n_472;
input n_296;
input n_265;
input n_746;
input n_208;
input n_456;
input n_156;
input n_292;
input n_793;
input n_174;
input n_275;
input n_100;
input n_704;
input n_132;
input n_147;
input n_204;
input n_751;
input n_615;
input n_521;
input n_51;
input n_496;
input n_739;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_792;
input n_824;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_719;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_773;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_803;
input n_134;
input n_329;
input n_718;
input n_185;
input n_340;
input n_749;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_815;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_782;
input n_425;
input n_431;
input n_811;
input n_508;
input n_624;
input n_118;
input n_121;
input n_791;
input n_618;
input n_411;
input n_484;
input n_712;
input n_353;
input n_22;
input n_736;
input n_767;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_191;
input n_382;
input n_797;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_828;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_799;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_796;
input n_805;
input n_127;
input n_531;
input n_783;
input n_675;

output n_2932;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_2484;
wire n_2866;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_1353;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_850;
wire n_1916;
wire n_2879;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_2818;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_1837;
wire n_924;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_2731;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_2646;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_2873;
wire n_1366;
wire n_2084;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_870;
wire n_2547;
wire n_1453;
wire n_958;
wire n_945;
wire n_2554;
wire n_2248;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_1761;
wire n_1062;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_2634;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_1944;
wire n_2233;
wire n_2370;
wire n_2663;
wire n_2914;
wire n_1988;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2782;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_2847;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_1900;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2332;
wire n_2391;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_2867;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_2739;
wire n_1597;
wire n_1771;
wire n_2902;
wire n_1544;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_2349;
wire n_1918;
wire n_2788;
wire n_1443;
wire n_1021;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_2909;
wire n_1461;
wire n_2717;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_1216;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_2038;
wire n_2263;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_1935;
wire n_2806;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_1819;
wire n_947;
wire n_2134;
wire n_1260;
wire n_930;
wire n_1179;
wire n_2703;
wire n_1442;
wire n_2926;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_1468;
wire n_1253;
wire n_1661;
wire n_2791;
wire n_2683;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_2015;
wire n_1972;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_2922;
wire n_2871;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_931;
wire n_1491;
wire n_2628;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_2659;
wire n_1139;
wire n_2836;
wire n_2439;
wire n_2864;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_2388;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_2898;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_976;
wire n_909;
wire n_1392;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_2895;
wire n_2903;
wire n_974;
wire n_1731;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_2467;
wire n_2768;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_2924;
wire n_1209;
wire n_1563;
wire n_1020;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_1483;
wire n_1363;
wire n_2681;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_2120;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_2860;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_2312;
wire n_2677;
wire n_1826;
wire n_2834;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_1592;
wire n_2812;
wire n_2662;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_2811;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_1365;
wire n_2476;
wire n_2814;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_1609;
wire n_1053;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_983;
wire n_2783;
wire n_2599;
wire n_1726;
wire n_2075;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_2418;
wire n_2496;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_2853;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2861;
wire n_2780;
wire n_1120;
wire n_1202;
wire n_2254;
wire n_1498;
wire n_1188;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_1402;
wire n_957;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_1005;
wire n_2379;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_845;
wire n_888;
wire n_2894;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_1919;
wire n_2508;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_890;
wire n_842;
wire n_1898;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_1895;
wire n_2821;
wire n_2690;
wire n_2474;
wire n_2623;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_1734;
wire n_1860;
wire n_2785;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_951;
wire n_2772;
wire n_862;
wire n_1700;
wire n_2637;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_2893;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_2737;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_2581;
wire n_1783;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_876;
wire n_1191;
wire n_2492;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_2900;
wire n_2026;
wire n_2912;
wire n_1786;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_1405;
wire n_2684;
wire n_2726;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_1499;
wire n_1318;
wire n_854;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_1526;
wire n_1305;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_1733;
wire n_1476;
wire n_1524;
wire n_1856;
wire n_2016;
wire n_2667;
wire n_2723;
wire n_2725;
wire n_2928;
wire n_943;
wire n_1118;
wire n_2905;
wire n_2884;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_1657;
wire n_878;
wire n_2857;
wire n_1784;
wire n_1321;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_1561;
wire n_2412;
wire n_2720;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_1154;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_2890;
wire n_2911;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_1151;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_2170;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_883;
wire n_1852;
wire n_1286;
wire n_2612;
wire n_1685;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_2892;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_858;
wire n_2796;
wire n_1185;
wire n_2475;
wire n_2804;
wire n_2173;
wire n_2715;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_1291;
wire n_2020;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_988;
wire n_914;
wire n_1116;
wire n_1958;
wire n_2747;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_1197;
wire n_2820;
wire n_2613;
wire n_1165;
wire n_1641;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_843;
wire n_2647;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_2666;
wire n_1370;
wire n_1603;
wire n_2401;
wire n_889;
wire n_1549;
wire n_1066;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2886;
wire n_2478;
wire n_911;
wire n_2658;
wire n_2608;
wire n_2920;
wire n_1712;
wire n_1403;
wire n_1534;
wire n_1065;
wire n_1948;
wire n_2767;
wire n_1290;
wire n_1959;
wire n_2396;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_2692;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_1194;
wire n_2862;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_918;
wire n_1968;
wire n_1885;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_1193;
wire n_1345;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2882;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_1612;
wire n_2498;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_2189;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_2204;
wire n_2931;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_875;
wire n_1617;
wire n_2455;
wire n_2600;
wire n_2231;
wire n_2828;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_2114;
wire n_2927;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_1221;
wire n_1785;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_1579;
wire n_2809;
wire n_2181;
wire n_2014;
wire n_975;
wire n_923;
wire n_1645;
wire n_1381;
wire n_1124;
wire n_2870;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2910;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2586;
wire n_1360;
wire n_973;
wire n_2858;
wire n_972;
wire n_2251;
wire n_2923;
wire n_2843;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2872;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_1411;
wire n_1359;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_1024;
wire n_2291;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_1775;
wire n_908;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_2630;
wire n_2794;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2901;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_1630;
wire n_1720;
wire n_2409;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_956;
wire n_1930;
wire n_1809;
wire n_2787;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_2395;
wire n_917;
wire n_2868;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_2212;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_2734;
wire n_2569;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_2897;
wire n_1322;
wire n_2583;
wire n_2918;
wire n_1473;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_1094;
wire n_1459;
wire n_840;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_1754;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_2775;
wire n_1212;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_2290;
wire n_2856;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1600;
wire n_1190;
wire n_1144;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_1915;
wire n_2360;
wire n_1393;
wire n_2240;
wire n_1369;
wire n_2846;
wire n_1781;
wire n_2917;
wire n_2544;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_2430;
wire n_2504;
wire n_910;
wire n_1410;
wire n_939;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_2587;
wire n_1347;
wire n_2839;
wire n_860;
wire n_1043;
wire n_2869;
wire n_1923;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_2644;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_2562;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_2673;
wire n_1591;
wire n_2585;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_2875;
wire n_1639;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_1581;
wire n_1928;
wire n_946;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_2081;
wire n_1474;
wire n_937;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1368;
wire n_1211;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_2880;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_2798;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_1871;
wire n_2514;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_2915;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_1308;
wire n_2851;
wire n_2823;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_734),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_325),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_565),
.Y(n_842)
);

CKINVDCx16_ASAP7_75t_R g843 ( 
.A(n_583),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_45),
.Y(n_844)
);

INVx1_ASAP7_75t_SL g845 ( 
.A(n_568),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_576),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_585),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_808),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_755),
.Y(n_849)
);

CKINVDCx20_ASAP7_75t_R g850 ( 
.A(n_503),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_161),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_60),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_574),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_598),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_229),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_208),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_558),
.Y(n_857)
);

CKINVDCx20_ASAP7_75t_R g858 ( 
.A(n_78),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_169),
.Y(n_859)
);

BUFx2_ASAP7_75t_L g860 ( 
.A(n_242),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_731),
.Y(n_861)
);

BUFx5_ASAP7_75t_L g862 ( 
.A(n_760),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_269),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_253),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_812),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_554),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_429),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_522),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_188),
.Y(n_869)
);

CKINVDCx20_ASAP7_75t_R g870 ( 
.A(n_743),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_22),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_561),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_555),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_33),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_468),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_279),
.Y(n_876)
);

INVx1_ASAP7_75t_SL g877 ( 
.A(n_741),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_738),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_297),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_778),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_776),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_580),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_307),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_337),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_60),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_189),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_703),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_99),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_439),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_554),
.Y(n_890)
);

CKINVDCx20_ASAP7_75t_R g891 ( 
.A(n_364),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_507),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_567),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_720),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_254),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_369),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_405),
.Y(n_897)
);

BUFx10_ASAP7_75t_L g898 ( 
.A(n_323),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_795),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_411),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_822),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_532),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_395),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_547),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_675),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_577),
.Y(n_906)
);

BUFx10_ASAP7_75t_L g907 ( 
.A(n_394),
.Y(n_907)
);

BUFx10_ASAP7_75t_L g908 ( 
.A(n_613),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_465),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_337),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_796),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_243),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_814),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_727),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_506),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_807),
.Y(n_916)
);

BUFx8_ASAP7_75t_SL g917 ( 
.A(n_695),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_684),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_763),
.Y(n_919)
);

BUFx10_ASAP7_75t_L g920 ( 
.A(n_357),
.Y(n_920)
);

CKINVDCx20_ASAP7_75t_R g921 ( 
.A(n_138),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_775),
.Y(n_922)
);

BUFx2_ASAP7_75t_SL g923 ( 
.A(n_544),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_833),
.Y(n_924)
);

INVx1_ASAP7_75t_SL g925 ( 
.A(n_794),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_427),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_747),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_384),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_603),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_793),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_379),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_135),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_185),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_246),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_737),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_552),
.Y(n_936)
);

BUFx2_ASAP7_75t_SL g937 ( 
.A(n_823),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_641),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_756),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_801),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_810),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_739),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_55),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_275),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_541),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_271),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_44),
.Y(n_947)
);

CKINVDCx14_ASAP7_75t_R g948 ( 
.A(n_203),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_522),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_798),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_815),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_767),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_38),
.Y(n_953)
);

BUFx10_ASAP7_75t_L g954 ( 
.A(n_706),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_186),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_402),
.Y(n_956)
);

BUFx10_ASAP7_75t_L g957 ( 
.A(n_331),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_148),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_612),
.Y(n_959)
);

CKINVDCx16_ASAP7_75t_R g960 ( 
.A(n_156),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_748),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_339),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_7),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_826),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_212),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_217),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_645),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_167),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_253),
.Y(n_969)
);

CKINVDCx16_ASAP7_75t_R g970 ( 
.A(n_714),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_732),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_305),
.Y(n_972)
);

CKINVDCx12_ASAP7_75t_R g973 ( 
.A(n_828),
.Y(n_973)
);

INVx1_ASAP7_75t_SL g974 ( 
.A(n_77),
.Y(n_974)
);

INVx1_ASAP7_75t_SL g975 ( 
.A(n_513),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_593),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_771),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_317),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_834),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_412),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_487),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_606),
.Y(n_982)
);

INVx2_ASAP7_75t_SL g983 ( 
.A(n_650),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_102),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_134),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_35),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_782),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_664),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_248),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_336),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_744),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_460),
.Y(n_992)
);

CKINVDCx20_ASAP7_75t_R g993 ( 
.A(n_686),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_103),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_518),
.Y(n_995)
);

INVx1_ASAP7_75t_SL g996 ( 
.A(n_451),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_434),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_555),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_259),
.Y(n_999)
);

BUFx5_ASAP7_75t_L g1000 ( 
.A(n_785),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_525),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_120),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_799),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_716),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_761),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_728),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_423),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_751),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_779),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_85),
.Y(n_1010)
);

CKINVDCx20_ASAP7_75t_R g1011 ( 
.A(n_811),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_236),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_9),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_173),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_560),
.Y(n_1015)
);

INVx2_ASAP7_75t_SL g1016 ( 
.A(n_514),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_676),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_569),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_240),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_708),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_84),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_772),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_750),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_777),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_547),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_511),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_248),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_363),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_35),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_757),
.Y(n_1030)
);

INVx1_ASAP7_75t_SL g1031 ( 
.A(n_316),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_699),
.Y(n_1032)
);

CKINVDCx20_ASAP7_75t_R g1033 ( 
.A(n_470),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_515),
.Y(n_1034)
);

BUFx8_ASAP7_75t_SL g1035 ( 
.A(n_832),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_789),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_595),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_500),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_176),
.Y(n_1039)
);

INVx1_ASAP7_75t_SL g1040 ( 
.A(n_169),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_397),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_781),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_153),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_384),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_273),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_802),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_759),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_752),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_210),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_770),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_725),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_797),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_350),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_552),
.Y(n_1054)
);

BUFx2_ASAP7_75t_L g1055 ( 
.A(n_216),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_246),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_49),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_800),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_280),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_194),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_533),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_820),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_484),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_232),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_510),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_477),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_669),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_193),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_590),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_238),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_109),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_620),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_573),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_717),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_11),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_13),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_400),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_99),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_339),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_34),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_586),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_657),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_766),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_719),
.Y(n_1084)
);

CKINVDCx20_ASAP7_75t_R g1085 ( 
.A(n_658),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_792),
.Y(n_1086)
);

INVx1_ASAP7_75t_SL g1087 ( 
.A(n_293),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_430),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_784),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_804),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_312),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_558),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_422),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_87),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_774),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_289),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_449),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_704),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_614),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_21),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_301),
.Y(n_1101)
);

INVx1_ASAP7_75t_SL g1102 ( 
.A(n_765),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_41),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_174),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_838),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_488),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_236),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_839),
.Y(n_1108)
);

CKINVDCx20_ASAP7_75t_R g1109 ( 
.A(n_553),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_340),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_564),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_482),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_666),
.Y(n_1113)
);

CKINVDCx16_ASAP7_75t_R g1114 ( 
.A(n_780),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_819),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_255),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_730),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_140),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_301),
.Y(n_1119)
);

CKINVDCx16_ASAP7_75t_R g1120 ( 
.A(n_296),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_813),
.Y(n_1121)
);

BUFx8_ASAP7_75t_SL g1122 ( 
.A(n_831),
.Y(n_1122)
);

CKINVDCx20_ASAP7_75t_R g1123 ( 
.A(n_721),
.Y(n_1123)
);

BUFx2_ASAP7_75t_SL g1124 ( 
.A(n_577),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_516),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_425),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_660),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_830),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_575),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_392),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_490),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_740),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_729),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_305),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_571),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_102),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_132),
.Y(n_1137)
);

CKINVDCx20_ASAP7_75t_R g1138 ( 
.A(n_16),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_489),
.Y(n_1139)
);

INVx2_ASAP7_75t_SL g1140 ( 
.A(n_722),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_566),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_758),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_821),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_803),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_397),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_540),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_733),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_682),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_616),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_86),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_790),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_476),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_570),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_326),
.Y(n_1154)
);

BUFx5_ASAP7_75t_L g1155 ( 
.A(n_563),
.Y(n_1155)
);

CKINVDCx20_ASAP7_75t_R g1156 ( 
.A(n_825),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_296),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_631),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_478),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_835),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_670),
.Y(n_1161)
);

CKINVDCx20_ASAP7_75t_R g1162 ( 
.A(n_334),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_809),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_226),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_242),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_764),
.Y(n_1166)
);

CKINVDCx20_ASAP7_75t_R g1167 ( 
.A(n_570),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_749),
.Y(n_1168)
);

CKINVDCx16_ASAP7_75t_R g1169 ( 
.A(n_818),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_594),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_597),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_306),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_736),
.Y(n_1173)
);

CKINVDCx20_ASAP7_75t_R g1174 ( 
.A(n_635),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_85),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_642),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_312),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_121),
.Y(n_1178)
);

CKINVDCx20_ASAP7_75t_R g1179 ( 
.A(n_723),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_506),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_410),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_566),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_285),
.Y(n_1183)
);

CKINVDCx20_ASAP7_75t_R g1184 ( 
.A(n_211),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_420),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_791),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_726),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_222),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_220),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_754),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_355),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_474),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_495),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_816),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_145),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_735),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_120),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_324),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_295),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_783),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_502),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_539),
.Y(n_1202)
);

CKINVDCx20_ASAP7_75t_R g1203 ( 
.A(n_604),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_559),
.Y(n_1204)
);

INVxp33_ASAP7_75t_SL g1205 ( 
.A(n_377),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_805),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_742),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_538),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_486),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_462),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_37),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_436),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_557),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_542),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_806),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_166),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_401),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_368),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_636),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_746),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_836),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_437),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_677),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_551),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_576),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_104),
.Y(n_1226)
);

INVx1_ASAP7_75t_SL g1227 ( 
.A(n_15),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_17),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_82),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_100),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_108),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_786),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_654),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_180),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_140),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_724),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_827),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_399),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_68),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_753),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_78),
.Y(n_1241)
);

CKINVDCx20_ASAP7_75t_R g1242 ( 
.A(n_683),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_82),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_318),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_829),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_787),
.Y(n_1246)
);

BUFx5_ASAP7_75t_L g1247 ( 
.A(n_629),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_181),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_773),
.Y(n_1249)
);

CKINVDCx11_ASAP7_75t_R g1250 ( 
.A(n_718),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_79),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_745),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_769),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_151),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_587),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_817),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_435),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_162),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_281),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_459),
.Y(n_1260)
);

CKINVDCx16_ASAP7_75t_R g1261 ( 
.A(n_762),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_562),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_23),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_611),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_359),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_442),
.Y(n_1266)
);

INVx1_ASAP7_75t_SL g1267 ( 
.A(n_581),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_443),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_662),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_768),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_112),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_369),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_837),
.Y(n_1273)
);

INVx2_ASAP7_75t_SL g1274 ( 
.A(n_556),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_572),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_550),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_788),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_493),
.Y(n_1278)
);

INVx1_ASAP7_75t_SL g1279 ( 
.A(n_396),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_184),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_824),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_50),
.Y(n_1282)
);

CKINVDCx20_ASAP7_75t_R g1283 ( 
.A(n_948),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_917),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1155),
.Y(n_1285)
);

CKINVDCx20_ASAP7_75t_R g1286 ( 
.A(n_870),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1155),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1155),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_R g1289 ( 
.A(n_993),
.B(n_578),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_1035),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_1122),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1250),
.Y(n_1292)
);

INVxp67_ASAP7_75t_L g1293 ( 
.A(n_860),
.Y(n_1293)
);

CKINVDCx20_ASAP7_75t_R g1294 ( 
.A(n_1011),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1155),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1155),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_960),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1120),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_841),
.Y(n_1299)
);

CKINVDCx14_ASAP7_75t_R g1300 ( 
.A(n_908),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_842),
.Y(n_1301)
);

CKINVDCx16_ASAP7_75t_R g1302 ( 
.A(n_843),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_855),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1085),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_866),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_875),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_884),
.Y(n_1307)
);

HB1xp67_ASAP7_75t_L g1308 ( 
.A(n_1045),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_892),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_902),
.Y(n_1310)
);

BUFx3_ASAP7_75t_L g1311 ( 
.A(n_1160),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1123),
.Y(n_1312)
);

CKINVDCx20_ASAP7_75t_R g1313 ( 
.A(n_1156),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_1174),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1179),
.Y(n_1315)
);

CKINVDCx20_ASAP7_75t_R g1316 ( 
.A(n_1203),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_1242),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1205),
.B(n_1),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1206),
.B(n_0),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_908),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_906),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1245),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_1255),
.Y(n_1323)
);

BUFx3_ASAP7_75t_L g1324 ( 
.A(n_954),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_1270),
.Y(n_1325)
);

CKINVDCx20_ASAP7_75t_R g1326 ( 
.A(n_850),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_844),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_909),
.Y(n_1328)
);

CKINVDCx20_ASAP7_75t_R g1329 ( 
.A(n_858),
.Y(n_1329)
);

INVxp67_ASAP7_75t_L g1330 ( 
.A(n_986),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_943),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_944),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_846),
.Y(n_1333)
);

INVxp33_ASAP7_75t_SL g1334 ( 
.A(n_1055),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_851),
.Y(n_1335)
);

INVx3_ASAP7_75t_L g1336 ( 
.A(n_1071),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_946),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_852),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_947),
.Y(n_1339)
);

CKINVDCx16_ASAP7_75t_R g1340 ( 
.A(n_970),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_956),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_958),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_969),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_978),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_927),
.B(n_0),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_984),
.Y(n_1346)
);

BUFx2_ASAP7_75t_L g1347 ( 
.A(n_1112),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_853),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_856),
.Y(n_1349)
);

CKINVDCx20_ASAP7_75t_R g1350 ( 
.A(n_890),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_857),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1285),
.Y(n_1352)
);

CKINVDCx8_ASAP7_75t_R g1353 ( 
.A(n_1284),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1287),
.Y(n_1354)
);

INVx3_ASAP7_75t_L g1355 ( 
.A(n_1336),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1297),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1288),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1295),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1296),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1300),
.B(n_959),
.Y(n_1360)
);

BUFx6f_ASAP7_75t_L g1361 ( 
.A(n_1320),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_1324),
.B(n_1101),
.Y(n_1362)
);

AND2x4_ASAP7_75t_L g1363 ( 
.A(n_1311),
.B(n_1150),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1299),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1301),
.A2(n_1170),
.B(n_878),
.Y(n_1365)
);

INVx1_ASAP7_75t_SL g1366 ( 
.A(n_1304),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1336),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1303),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1305),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1306),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1307),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1309),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1310),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1321),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1328),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1302),
.B(n_1114),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1298),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1331),
.Y(n_1378)
);

NAND3xp33_ASAP7_75t_L g1379 ( 
.A(n_1293),
.B(n_863),
.C(n_859),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1332),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1337),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1339),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1341),
.Y(n_1383)
);

INVxp67_ASAP7_75t_L g1384 ( 
.A(n_1347),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1340),
.B(n_1169),
.Y(n_1385)
);

INVx3_ASAP7_75t_L g1386 ( 
.A(n_1342),
.Y(n_1386)
);

INVxp67_ASAP7_75t_L g1387 ( 
.A(n_1308),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1343),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1344),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1346),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1345),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1319),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1330),
.B(n_893),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1327),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1333),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_SL g1396 ( 
.A(n_1335),
.B(n_1261),
.Y(n_1396)
);

BUFx6f_ASAP7_75t_L g1397 ( 
.A(n_1338),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1348),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1349),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1351),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1292),
.Y(n_1401)
);

NAND2xp33_ASAP7_75t_R g1402 ( 
.A(n_1334),
.B(n_864),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_1318),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1289),
.B(n_1161),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1283),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1290),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_SL g1407 ( 
.A1(n_1326),
.A2(n_896),
.B1(n_921),
.B2(n_891),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1291),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1312),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_SL g1410 ( 
.A1(n_1407),
.A2(n_1315),
.B1(n_1317),
.B2(n_1314),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1384),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1357),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1374),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1391),
.B(n_1200),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1361),
.B(n_1286),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1387),
.Y(n_1416)
);

INVx1_ASAP7_75t_SL g1417 ( 
.A(n_1366),
.Y(n_1417)
);

AND2x6_ASAP7_75t_L g1418 ( 
.A(n_1397),
.B(n_845),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1361),
.B(n_1294),
.Y(n_1419)
);

BUFx10_ASAP7_75t_L g1420 ( 
.A(n_1397),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1380),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1404),
.B(n_1322),
.Y(n_1422)
);

INVxp67_ASAP7_75t_SL g1423 ( 
.A(n_1355),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1383),
.Y(n_1424)
);

INVx1_ASAP7_75t_SL g1425 ( 
.A(n_1376),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1385),
.B(n_1323),
.Y(n_1426)
);

CKINVDCx20_ASAP7_75t_R g1427 ( 
.A(n_1409),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1392),
.A2(n_1274),
.B1(n_1016),
.B2(n_933),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1403),
.A2(n_867),
.B1(n_869),
.B2(n_868),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1367),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1354),
.B(n_1358),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1393),
.A2(n_1018),
.B1(n_1118),
.B2(n_900),
.Y(n_1432)
);

AO22x2_ASAP7_75t_L g1433 ( 
.A1(n_1405),
.A2(n_1350),
.B1(n_1329),
.B2(n_1313),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1364),
.Y(n_1434)
);

INVx6_ASAP7_75t_L g1435 ( 
.A(n_1363),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1386),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_1353),
.Y(n_1437)
);

BUFx2_ASAP7_75t_L g1438 ( 
.A(n_1356),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1368),
.Y(n_1439)
);

OR2x6_ASAP7_75t_L g1440 ( 
.A(n_1401),
.B(n_1406),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1359),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1369),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1370),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1371),
.Y(n_1444)
);

BUFx6f_ASAP7_75t_L g1445 ( 
.A(n_1365),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1403),
.B(n_1325),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1377),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1360),
.B(n_1215),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1372),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_SL g1450 ( 
.A(n_1395),
.B(n_871),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_SL g1451 ( 
.A(n_1398),
.B(n_872),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1373),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_SL g1453 ( 
.A(n_1394),
.B(n_873),
.Y(n_1453)
);

INVx5_ASAP7_75t_L g1454 ( 
.A(n_1362),
.Y(n_1454)
);

INVx4_ASAP7_75t_L g1455 ( 
.A(n_1393),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1375),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_1378),
.Y(n_1457)
);

AOI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1402),
.A2(n_1279),
.B1(n_975),
.B2(n_996),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1399),
.B(n_1316),
.Y(n_1459)
);

INVx5_ASAP7_75t_L g1460 ( 
.A(n_1408),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1400),
.B(n_1273),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1381),
.Y(n_1462)
);

INVx3_ASAP7_75t_L g1463 ( 
.A(n_1382),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1388),
.B(n_1033),
.Y(n_1464)
);

AND2x4_ASAP7_75t_L g1465 ( 
.A(n_1389),
.B(n_1109),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1390),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1379),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1396),
.B(n_1281),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1352),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1355),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1374),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1374),
.Y(n_1472)
);

AND2x4_ASAP7_75t_L g1473 ( 
.A(n_1361),
.B(n_1138),
.Y(n_1473)
);

INVx4_ASAP7_75t_L g1474 ( 
.A(n_1397),
.Y(n_1474)
);

INVx2_ASAP7_75t_SL g1475 ( 
.A(n_1397),
.Y(n_1475)
);

INVx2_ASAP7_75t_SL g1476 ( 
.A(n_1397),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_SL g1477 ( 
.A(n_1404),
.B(n_874),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_SL g1478 ( 
.A(n_1404),
.B(n_876),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1434),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1461),
.B(n_877),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1417),
.B(n_974),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1439),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1442),
.Y(n_1483)
);

OR2x6_ASAP7_75t_L g1484 ( 
.A(n_1475),
.B(n_923),
.Y(n_1484)
);

AOI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1468),
.A2(n_1167),
.B1(n_1184),
.B2(n_1162),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1443),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1413),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1444),
.Y(n_1488)
);

AND2x2_ASAP7_75t_SL g1489 ( 
.A(n_1438),
.B(n_1136),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1449),
.Y(n_1490)
);

OR2x2_ASAP7_75t_SL g1491 ( 
.A(n_1411),
.B(n_1193),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1421),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1456),
.Y(n_1493)
);

AO22x2_ASAP7_75t_L g1494 ( 
.A1(n_1425),
.A2(n_1040),
.B1(n_1087),
.B2(n_1031),
.Y(n_1494)
);

NAND2x1p5_ASAP7_75t_L g1495 ( 
.A(n_1474),
.B(n_1227),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1412),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1469),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1430),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1424),
.Y(n_1499)
);

INVx2_ASAP7_75t_SL g1500 ( 
.A(n_1420),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1471),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1472),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1462),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1452),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1466),
.Y(n_1505)
);

AO22x2_ASAP7_75t_L g1506 ( 
.A1(n_1464),
.A2(n_1465),
.B1(n_1459),
.B2(n_1419),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1452),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1463),
.Y(n_1508)
);

OAI221xp5_ASAP7_75t_L g1509 ( 
.A1(n_1428),
.A2(n_998),
.B1(n_999),
.B2(n_997),
.C(n_985),
.Y(n_1509)
);

NAND2x1p5_ASAP7_75t_L g1510 ( 
.A(n_1476),
.B(n_925),
.Y(n_1510)
);

AO22x2_ASAP7_75t_L g1511 ( 
.A1(n_1415),
.A2(n_1124),
.B1(n_1012),
.B2(n_1013),
.Y(n_1511)
);

AO22x2_ASAP7_75t_L g1512 ( 
.A1(n_1426),
.A2(n_1473),
.B1(n_1433),
.B2(n_1422),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1416),
.Y(n_1513)
);

NAND2xp33_ASAP7_75t_L g1514 ( 
.A(n_1445),
.B(n_879),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1437),
.B(n_1007),
.Y(n_1515)
);

AO22x2_ASAP7_75t_L g1516 ( 
.A1(n_1410),
.A2(n_1448),
.B1(n_1455),
.B2(n_1446),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1431),
.Y(n_1517)
);

AO22x2_ASAP7_75t_L g1518 ( 
.A1(n_1429),
.A2(n_1015),
.B1(n_1019),
.B2(n_1014),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1457),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1467),
.B(n_1282),
.Y(n_1520)
);

INVx3_ASAP7_75t_L g1521 ( 
.A(n_1435),
.Y(n_1521)
);

AOI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1457),
.A2(n_983),
.B1(n_1140),
.B2(n_1050),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1441),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1441),
.A2(n_1148),
.B1(n_937),
.B2(n_887),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1436),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1423),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1470),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1414),
.B(n_1477),
.Y(n_1528)
);

OAI221xp5_ASAP7_75t_L g1529 ( 
.A1(n_1432),
.A2(n_1276),
.B1(n_1280),
.B2(n_1275),
.C(n_1272),
.Y(n_1529)
);

AND2x6_ASAP7_75t_L g1530 ( 
.A(n_1445),
.B(n_1170),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1450),
.Y(n_1531)
);

INVx3_ASAP7_75t_R g1532 ( 
.A(n_1447),
.Y(n_1532)
);

NAND2x1p5_ASAP7_75t_L g1533 ( 
.A(n_1454),
.B(n_1102),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1451),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_1427),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1453),
.Y(n_1536)
);

AO22x2_ASAP7_75t_L g1537 ( 
.A1(n_1458),
.A2(n_1025),
.B1(n_1026),
.B2(n_1021),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1478),
.A2(n_894),
.B1(n_899),
.B2(n_865),
.Y(n_1538)
);

NAND2x1p5_ASAP7_75t_L g1539 ( 
.A(n_1454),
.B(n_1267),
.Y(n_1539)
);

OAI221xp5_ASAP7_75t_L g1540 ( 
.A1(n_1460),
.A2(n_1056),
.B1(n_1057),
.B2(n_1054),
.C(n_1034),
.Y(n_1540)
);

INVx2_ASAP7_75t_SL g1541 ( 
.A(n_1440),
.Y(n_1541)
);

AND2x4_ASAP7_75t_L g1542 ( 
.A(n_1418),
.B(n_1063),
.Y(n_1542)
);

AO22x2_ASAP7_75t_L g1543 ( 
.A1(n_1418),
.A2(n_1068),
.B1(n_1073),
.B2(n_1064),
.Y(n_1543)
);

OAI221xp5_ASAP7_75t_L g1544 ( 
.A1(n_1468),
.A2(n_1092),
.B1(n_1096),
.B2(n_1088),
.C(n_1078),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1416),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1461),
.B(n_949),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1434),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1434),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1434),
.Y(n_1549)
);

AO22x2_ASAP7_75t_L g1550 ( 
.A1(n_1417),
.A2(n_1104),
.B1(n_1106),
.B2(n_1100),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1417),
.B(n_1110),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1417),
.B(n_1119),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1434),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1413),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1416),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1434),
.Y(n_1556)
);

AOI22x1_ASAP7_75t_SL g1557 ( 
.A1(n_1437),
.A2(n_885),
.B1(n_886),
.B2(n_883),
.Y(n_1557)
);

CKINVDCx20_ASAP7_75t_R g1558 ( 
.A(n_1437),
.Y(n_1558)
);

CKINVDCx16_ASAP7_75t_R g1559 ( 
.A(n_1420),
.Y(n_1559)
);

AO22x2_ASAP7_75t_L g1560 ( 
.A1(n_1417),
.A2(n_1129),
.B1(n_1134),
.B2(n_1126),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1434),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1434),
.Y(n_1562)
);

INVxp67_ASAP7_75t_L g1563 ( 
.A(n_1416),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1461),
.B(n_949),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1434),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_L g1566 ( 
.A(n_1417),
.B(n_1260),
.Y(n_1566)
);

NAND2x1p5_ASAP7_75t_L g1567 ( 
.A(n_1474),
.B(n_1146),
.Y(n_1567)
);

OAI221xp5_ASAP7_75t_L g1568 ( 
.A1(n_1468),
.A2(n_1157),
.B1(n_1178),
.B2(n_1159),
.C(n_1153),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1420),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1413),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1417),
.B(n_898),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1434),
.Y(n_1572)
);

AO22x2_ASAP7_75t_L g1573 ( 
.A1(n_1417),
.A2(n_1182),
.B1(n_1195),
.B2(n_1183),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1417),
.B(n_1271),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1434),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1461),
.B(n_949),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1417),
.B(n_898),
.Y(n_1577)
);

AND2x2_ASAP7_75t_SL g1578 ( 
.A(n_1438),
.B(n_1145),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1434),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1434),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1434),
.Y(n_1581)
);

CKINVDCx16_ASAP7_75t_R g1582 ( 
.A(n_1420),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1413),
.Y(n_1583)
);

OAI221xp5_ASAP7_75t_L g1584 ( 
.A1(n_1468),
.A2(n_1208),
.B1(n_1213),
.B2(n_1198),
.C(n_1197),
.Y(n_1584)
);

INVxp67_ASAP7_75t_L g1585 ( 
.A(n_1416),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1413),
.Y(n_1586)
);

AO22x2_ASAP7_75t_L g1587 ( 
.A1(n_1417),
.A2(n_1224),
.B1(n_1234),
.B2(n_1228),
.Y(n_1587)
);

AOI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1468),
.A2(n_929),
.B1(n_935),
.B2(n_918),
.Y(n_1588)
);

AO22x2_ASAP7_75t_L g1589 ( 
.A1(n_1417),
.A2(n_1259),
.B1(n_1238),
.B2(n_1210),
.Y(n_1589)
);

INVxp67_ASAP7_75t_L g1590 ( 
.A(n_1416),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1461),
.B(n_1152),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1434),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1434),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1434),
.Y(n_1594)
);

AO22x2_ASAP7_75t_L g1595 ( 
.A1(n_1417),
.A2(n_1216),
.B1(n_1217),
.B2(n_1202),
.Y(n_1595)
);

AO22x2_ASAP7_75t_L g1596 ( 
.A1(n_1417),
.A2(n_907),
.B1(n_957),
.B2(n_920),
.Y(n_1596)
);

NAND2x1p5_ASAP7_75t_L g1597 ( 
.A(n_1474),
.B(n_1048),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1434),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1416),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_SL g1600 ( 
.A1(n_1418),
.A2(n_920),
.B1(n_907),
.B2(n_957),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1461),
.B(n_1152),
.Y(n_1601)
);

NAND2xp33_ASAP7_75t_SL g1602 ( 
.A(n_1532),
.B(n_888),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1489),
.B(n_889),
.Y(n_1603)
);

NAND2xp33_ASAP7_75t_SL g1604 ( 
.A(n_1500),
.B(n_895),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_SL g1605 ( 
.A(n_1585),
.B(n_897),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1590),
.B(n_903),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_SL g1607 ( 
.A(n_1578),
.B(n_904),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1517),
.B(n_910),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1480),
.B(n_912),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_SL g1610 ( 
.A(n_1528),
.B(n_915),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_SL g1611 ( 
.A(n_1513),
.B(n_926),
.Y(n_1611)
);

NAND2xp33_ASAP7_75t_SL g1612 ( 
.A(n_1569),
.B(n_928),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_SL g1613 ( 
.A(n_1545),
.B(n_931),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1555),
.B(n_932),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_SL g1615 ( 
.A(n_1599),
.B(n_934),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_SL g1616 ( 
.A(n_1559),
.B(n_936),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1541),
.B(n_941),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_SL g1618 ( 
.A(n_1582),
.B(n_945),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1526),
.B(n_953),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1481),
.B(n_955),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1504),
.B(n_950),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1566),
.B(n_962),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1574),
.B(n_1508),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_SL g1624 ( 
.A(n_1507),
.B(n_963),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_SL g1625 ( 
.A(n_1523),
.B(n_965),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_SL g1626 ( 
.A(n_1519),
.B(n_966),
.Y(n_1626)
);

XNOR2x2_ASAP7_75t_L g1627 ( 
.A(n_1485),
.B(n_951),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_SL g1628 ( 
.A(n_1536),
.B(n_968),
.Y(n_1628)
);

NAND2xp33_ASAP7_75t_SL g1629 ( 
.A(n_1558),
.B(n_972),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_SL g1630 ( 
.A(n_1531),
.B(n_980),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_SL g1631 ( 
.A(n_1534),
.B(n_1520),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_SL g1632 ( 
.A(n_1479),
.B(n_981),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_SL g1633 ( 
.A(n_1482),
.B(n_989),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1483),
.B(n_990),
.Y(n_1634)
);

NAND2xp33_ASAP7_75t_SL g1635 ( 
.A(n_1486),
.B(n_992),
.Y(n_1635)
);

NAND2xp33_ASAP7_75t_SL g1636 ( 
.A(n_1488),
.B(n_994),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_SL g1637 ( 
.A(n_1490),
.B(n_995),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1493),
.B(n_1001),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1547),
.B(n_1002),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_SL g1640 ( 
.A(n_1548),
.B(n_1010),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1571),
.B(n_1027),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_SL g1642 ( 
.A(n_1549),
.B(n_1028),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_L g1643 ( 
.A(n_1577),
.B(n_1029),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_SL g1644 ( 
.A(n_1553),
.B(n_1038),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_SL g1645 ( 
.A(n_1556),
.B(n_1039),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1561),
.B(n_1041),
.Y(n_1646)
);

NAND2xp33_ASAP7_75t_SL g1647 ( 
.A(n_1562),
.B(n_1043),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_SL g1648 ( 
.A(n_1565),
.B(n_1044),
.Y(n_1648)
);

NAND2xp33_ASAP7_75t_SL g1649 ( 
.A(n_1572),
.B(n_1049),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_SL g1650 ( 
.A(n_1575),
.B(n_1053),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_SL g1651 ( 
.A(n_1579),
.B(n_1059),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1535),
.B(n_1060),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_SL g1653 ( 
.A(n_1580),
.B(n_1061),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1581),
.B(n_1065),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1592),
.B(n_1066),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_SL g1656 ( 
.A(n_1593),
.B(n_1070),
.Y(n_1656)
);

NAND2xp33_ASAP7_75t_SL g1657 ( 
.A(n_1594),
.B(n_1598),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_SL g1658 ( 
.A(n_1588),
.B(n_1075),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1546),
.B(n_1076),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_SL g1660 ( 
.A(n_1601),
.B(n_1077),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_SL g1661 ( 
.A(n_1564),
.B(n_1079),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1576),
.B(n_1080),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_SL g1663 ( 
.A(n_1591),
.B(n_1524),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_SL g1664 ( 
.A(n_1538),
.B(n_1091),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_SL g1665 ( 
.A(n_1527),
.B(n_1093),
.Y(n_1665)
);

NAND2xp33_ASAP7_75t_SL g1666 ( 
.A(n_1525),
.B(n_1094),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_SL g1667 ( 
.A(n_1515),
.B(n_1097),
.Y(n_1667)
);

NAND2xp33_ASAP7_75t_SL g1668 ( 
.A(n_1503),
.B(n_1103),
.Y(n_1668)
);

NAND2xp33_ASAP7_75t_SL g1669 ( 
.A(n_1505),
.B(n_1107),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1551),
.B(n_1111),
.Y(n_1670)
);

NAND2xp33_ASAP7_75t_SL g1671 ( 
.A(n_1499),
.B(n_1116),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_SL g1672 ( 
.A(n_1495),
.B(n_1125),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_SL g1673 ( 
.A(n_1567),
.B(n_1130),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_SL g1674 ( 
.A(n_1522),
.B(n_1131),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1501),
.B(n_1135),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_SL g1676 ( 
.A(n_1510),
.B(n_1502),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_SL g1677 ( 
.A(n_1533),
.B(n_1137),
.Y(n_1677)
);

NAND2xp33_ASAP7_75t_SL g1678 ( 
.A(n_1498),
.B(n_1139),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1539),
.B(n_1141),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1552),
.B(n_1154),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_SL g1681 ( 
.A(n_1600),
.B(n_1164),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_SL g1682 ( 
.A(n_1521),
.B(n_1165),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_SL g1683 ( 
.A(n_1597),
.B(n_1172),
.Y(n_1683)
);

NAND2xp33_ASAP7_75t_SL g1684 ( 
.A(n_1514),
.B(n_1177),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1487),
.B(n_1180),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_SL g1686 ( 
.A(n_1542),
.B(n_1181),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1550),
.B(n_1185),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1492),
.B(n_1188),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_SL g1689 ( 
.A(n_1496),
.B(n_1189),
.Y(n_1689)
);

NAND2xp33_ASAP7_75t_SL g1690 ( 
.A(n_1497),
.B(n_1191),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1554),
.B(n_1192),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1570),
.B(n_1199),
.Y(n_1692)
);

NAND2xp33_ASAP7_75t_SL g1693 ( 
.A(n_1583),
.B(n_1201),
.Y(n_1693)
);

NAND2xp33_ASAP7_75t_SL g1694 ( 
.A(n_1586),
.B(n_1204),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1530),
.B(n_1209),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_SL g1696 ( 
.A(n_1516),
.B(n_1211),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1530),
.B(n_1212),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_SL g1698 ( 
.A(n_1484),
.B(n_1214),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_SL g1699 ( 
.A(n_1518),
.B(n_1218),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_SL g1700 ( 
.A(n_1506),
.B(n_1222),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_SL g1701 ( 
.A(n_1543),
.B(n_1225),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1512),
.B(n_976),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_SL g1703 ( 
.A(n_1544),
.B(n_1226),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_SL g1704 ( 
.A(n_1568),
.B(n_1229),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_SL g1705 ( 
.A(n_1584),
.B(n_1230),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_SL g1706 ( 
.A(n_1540),
.B(n_1231),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_SL g1707 ( 
.A(n_1491),
.B(n_1235),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1595),
.B(n_1239),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1537),
.B(n_1241),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_SL g1710 ( 
.A(n_1557),
.B(n_1243),
.Y(n_1710)
);

NAND2xp33_ASAP7_75t_SL g1711 ( 
.A(n_1511),
.B(n_1244),
.Y(n_1711)
);

NAND2xp33_ASAP7_75t_SL g1712 ( 
.A(n_1509),
.B(n_1248),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_SL g1713 ( 
.A(n_1589),
.B(n_1251),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1560),
.B(n_1254),
.Y(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1573),
.B(n_982),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_SL g1716 ( 
.A(n_1587),
.B(n_1257),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_SL g1717 ( 
.A(n_1596),
.B(n_1258),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_SL g1718 ( 
.A(n_1529),
.B(n_1262),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_SL g1719 ( 
.A(n_1494),
.B(n_1263),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_SL g1720 ( 
.A(n_1563),
.B(n_1265),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_SL g1721 ( 
.A(n_1563),
.B(n_1266),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1517),
.B(n_1268),
.Y(n_1722)
);

NAND2xp33_ASAP7_75t_SL g1723 ( 
.A(n_1532),
.B(n_1175),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1489),
.B(n_1175),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1513),
.B(n_1278),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_SL g1726 ( 
.A(n_1563),
.B(n_1278),
.Y(n_1726)
);

AND2x6_ASAP7_75t_L g1727 ( 
.A(n_1517),
.B(n_847),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1563),
.B(n_840),
.Y(n_1728)
);

NAND2xp33_ASAP7_75t_SL g1729 ( 
.A(n_1532),
.B(n_1249),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1563),
.B(n_848),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_SL g1731 ( 
.A(n_1563),
.B(n_849),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1517),
.B(n_988),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_SL g1733 ( 
.A(n_1563),
.B(n_854),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_SL g1734 ( 
.A(n_1563),
.B(n_861),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1489),
.B(n_1),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1569),
.B(n_1004),
.Y(n_1736)
);

NAND2xp33_ASAP7_75t_SL g1737 ( 
.A(n_1532),
.B(n_1253),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_SL g1738 ( 
.A(n_1563),
.B(n_880),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_SL g1739 ( 
.A(n_1563),
.B(n_881),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_SL g1740 ( 
.A(n_1563),
.B(n_901),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_SL g1741 ( 
.A(n_1563),
.B(n_911),
.Y(n_1741)
);

XNOR2x2_ASAP7_75t_L g1742 ( 
.A(n_1485),
.B(n_1005),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1517),
.B(n_1221),
.Y(n_1743)
);

NAND2xp33_ASAP7_75t_SL g1744 ( 
.A(n_1532),
.B(n_1252),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_SL g1745 ( 
.A(n_1563),
.B(n_913),
.Y(n_1745)
);

NAND2xp33_ASAP7_75t_R g1746 ( 
.A(n_1535),
.B(n_914),
.Y(n_1746)
);

NAND2xp33_ASAP7_75t_SL g1747 ( 
.A(n_1532),
.B(n_1269),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_SL g1748 ( 
.A(n_1563),
.B(n_916),
.Y(n_1748)
);

NAND2xp33_ASAP7_75t_SL g1749 ( 
.A(n_1532),
.B(n_1236),
.Y(n_1749)
);

NAND2xp33_ASAP7_75t_SL g1750 ( 
.A(n_1532),
.B(n_1237),
.Y(n_1750)
);

NAND2xp33_ASAP7_75t_SL g1751 ( 
.A(n_1532),
.B(n_1240),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_SL g1752 ( 
.A(n_1563),
.B(n_919),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1517),
.B(n_1008),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_SL g1754 ( 
.A(n_1563),
.B(n_922),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1517),
.B(n_1022),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1517),
.B(n_1024),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_SL g1757 ( 
.A(n_1563),
.B(n_924),
.Y(n_1757)
);

NAND2xp33_ASAP7_75t_SL g1758 ( 
.A(n_1532),
.B(n_1232),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_SL g1759 ( 
.A(n_1563),
.B(n_930),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_SL g1760 ( 
.A(n_1563),
.B(n_938),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_SL g1761 ( 
.A(n_1563),
.B(n_939),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1517),
.B(n_1207),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_SL g1763 ( 
.A(n_1563),
.B(n_940),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_SL g1764 ( 
.A(n_1563),
.B(n_942),
.Y(n_1764)
);

NAND2xp33_ASAP7_75t_SL g1765 ( 
.A(n_1532),
.B(n_952),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_SL g1766 ( 
.A(n_1563),
.B(n_961),
.Y(n_1766)
);

NAND2xp33_ASAP7_75t_SL g1767 ( 
.A(n_1532),
.B(n_1246),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1563),
.B(n_1030),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1489),
.B(n_2),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1489),
.B(n_2),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_SL g1771 ( 
.A(n_1563),
.B(n_964),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1489),
.B(n_3),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_SL g1773 ( 
.A(n_1563),
.B(n_967),
.Y(n_1773)
);

O2A1O1Ixp5_ASAP7_75t_L g1774 ( 
.A1(n_1657),
.A2(n_1051),
.B(n_1052),
.C(n_1042),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1620),
.B(n_1603),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1643),
.B(n_4),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1621),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1641),
.B(n_4),
.Y(n_1778)
);

OAI21x1_ASAP7_75t_L g1779 ( 
.A1(n_1663),
.A2(n_1082),
.B(n_1062),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1609),
.B(n_5),
.Y(n_1780)
);

AOI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1610),
.A2(n_1117),
.B(n_1113),
.Y(n_1781)
);

OAI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1608),
.A2(n_1722),
.B1(n_1743),
.B2(n_1732),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1680),
.B(n_5),
.Y(n_1783)
);

AO21x1_ASAP7_75t_L g1784 ( 
.A1(n_1696),
.A2(n_1144),
.B(n_1132),
.Y(n_1784)
);

AOI211x1_ASAP7_75t_L g1785 ( 
.A1(n_1632),
.A2(n_1171),
.B(n_1190),
.C(n_1166),
.Y(n_1785)
);

BUFx6f_ASAP7_75t_L g1786 ( 
.A(n_1736),
.Y(n_1786)
);

OAI21x1_ASAP7_75t_L g1787 ( 
.A1(n_1753),
.A2(n_1223),
.B(n_1196),
.Y(n_1787)
);

AOI21xp5_ASAP7_75t_SL g1788 ( 
.A1(n_1755),
.A2(n_1058),
.B(n_882),
.Y(n_1788)
);

NAND3xp33_ASAP7_75t_L g1789 ( 
.A(n_1768),
.B(n_1233),
.C(n_1036),
.Y(n_1789)
);

OAI21xp5_ASAP7_75t_L g1790 ( 
.A1(n_1756),
.A2(n_1264),
.B(n_1219),
.Y(n_1790)
);

BUFx6f_ASAP7_75t_L g1791 ( 
.A(n_1736),
.Y(n_1791)
);

AO31x2_ASAP7_75t_L g1792 ( 
.A1(n_1762),
.A2(n_1194),
.A3(n_905),
.B(n_1000),
.Y(n_1792)
);

OAI21xp5_ASAP7_75t_SL g1793 ( 
.A1(n_1652),
.A2(n_6),
.B(n_7),
.Y(n_1793)
);

OAI21x1_ASAP7_75t_L g1794 ( 
.A1(n_1676),
.A2(n_1689),
.B(n_1688),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1685),
.Y(n_1795)
);

AO31x2_ASAP7_75t_L g1796 ( 
.A1(n_1708),
.A2(n_862),
.A3(n_1247),
.B(n_1000),
.Y(n_1796)
);

OAI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1623),
.A2(n_1646),
.B(n_1634),
.Y(n_1797)
);

AO21x2_ASAP7_75t_L g1798 ( 
.A1(n_1659),
.A2(n_973),
.B(n_862),
.Y(n_1798)
);

AOI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1660),
.A2(n_1662),
.B(n_1661),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1654),
.Y(n_1800)
);

A2O1A1Ixp33_ASAP7_75t_L g1801 ( 
.A1(n_1712),
.A2(n_1046),
.B(n_1074),
.C(n_1003),
.Y(n_1801)
);

OAI21x1_ASAP7_75t_SL g1802 ( 
.A1(n_1695),
.A2(n_8),
.B(n_9),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1631),
.B(n_971),
.Y(n_1803)
);

BUFx10_ASAP7_75t_L g1804 ( 
.A(n_1617),
.Y(n_1804)
);

NAND3xp33_ASAP7_75t_L g1805 ( 
.A(n_1622),
.B(n_979),
.C(n_977),
.Y(n_1805)
);

OAI21x1_ASAP7_75t_L g1806 ( 
.A1(n_1691),
.A2(n_1000),
.B(n_862),
.Y(n_1806)
);

AND2x6_ASAP7_75t_L g1807 ( 
.A(n_1735),
.B(n_847),
.Y(n_1807)
);

OAI21x1_ASAP7_75t_L g1808 ( 
.A1(n_1692),
.A2(n_1000),
.B(n_862),
.Y(n_1808)
);

NAND2x1p5_ASAP7_75t_L g1809 ( 
.A(n_1715),
.B(n_847),
.Y(n_1809)
);

AND2x4_ASAP7_75t_L g1810 ( 
.A(n_1724),
.B(n_10),
.Y(n_1810)
);

AOI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1628),
.A2(n_1256),
.B(n_1220),
.Y(n_1811)
);

AOI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1769),
.A2(n_1770),
.B1(n_1772),
.B2(n_1746),
.Y(n_1812)
);

OAI21xp5_ASAP7_75t_L g1813 ( 
.A1(n_1655),
.A2(n_1006),
.B(n_991),
.Y(n_1813)
);

AND2x4_ASAP7_75t_L g1814 ( 
.A(n_1617),
.B(n_10),
.Y(n_1814)
);

AOI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1630),
.A2(n_1017),
.B(n_1009),
.Y(n_1815)
);

OAI21x1_ASAP7_75t_L g1816 ( 
.A1(n_1624),
.A2(n_1000),
.B(n_862),
.Y(n_1816)
);

BUFx10_ASAP7_75t_L g1817 ( 
.A(n_1715),
.Y(n_1817)
);

OAI21x1_ASAP7_75t_L g1818 ( 
.A1(n_1625),
.A2(n_1247),
.B(n_582),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_SL g1819 ( 
.A(n_1635),
.B(n_1149),
.Y(n_1819)
);

OAI21x1_ASAP7_75t_L g1820 ( 
.A1(n_1626),
.A2(n_1247),
.B(n_584),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1675),
.B(n_1607),
.Y(n_1821)
);

AOI21xp5_ASAP7_75t_L g1822 ( 
.A1(n_1619),
.A2(n_1163),
.B(n_1158),
.Y(n_1822)
);

BUFx2_ASAP7_75t_R g1823 ( 
.A(n_1707),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1702),
.B(n_11),
.Y(n_1824)
);

AOI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1633),
.A2(n_1176),
.B(n_1173),
.Y(n_1825)
);

AOI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1637),
.A2(n_1277),
.B(n_1032),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1702),
.B(n_12),
.Y(n_1827)
);

OAI21x1_ASAP7_75t_SL g1828 ( 
.A1(n_1697),
.A2(n_1742),
.B(n_1627),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1725),
.Y(n_1829)
);

AOI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1638),
.A2(n_1037),
.B(n_1023),
.Y(n_1830)
);

NOR2xp67_ASAP7_75t_L g1831 ( 
.A(n_1670),
.B(n_1047),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1703),
.B(n_12),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1704),
.B(n_1705),
.Y(n_1833)
);

OA22x2_ASAP7_75t_L g1834 ( 
.A1(n_1699),
.A2(n_1098),
.B1(n_1115),
.B2(n_1072),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1636),
.B(n_1128),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1639),
.Y(n_1836)
);

AO21x1_ASAP7_75t_L g1837 ( 
.A1(n_1711),
.A2(n_1247),
.B(n_987),
.Y(n_1837)
);

AOI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1640),
.A2(n_1142),
.B(n_1133),
.Y(n_1838)
);

OAI21x1_ASAP7_75t_L g1839 ( 
.A1(n_1665),
.A2(n_1247),
.B(n_588),
.Y(n_1839)
);

BUFx2_ASAP7_75t_SL g1840 ( 
.A(n_1616),
.Y(n_1840)
);

AOI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1642),
.A2(n_1168),
.B(n_1151),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1718),
.B(n_13),
.Y(n_1842)
);

INVx2_ASAP7_75t_SL g1843 ( 
.A(n_1682),
.Y(n_1843)
);

BUFx6f_ASAP7_75t_L g1844 ( 
.A(n_1677),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1687),
.B(n_14),
.Y(n_1845)
);

AOI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1644),
.A2(n_1069),
.B(n_1067),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1645),
.Y(n_1847)
);

AOI22xp5_ASAP7_75t_L g1848 ( 
.A1(n_1647),
.A2(n_1083),
.B1(n_1084),
.B2(n_1081),
.Y(n_1848)
);

AOI21x1_ASAP7_75t_L g1849 ( 
.A1(n_1648),
.A2(n_987),
.B(n_882),
.Y(n_1849)
);

AO31x2_ASAP7_75t_L g1850 ( 
.A1(n_1714),
.A2(n_987),
.A3(n_1020),
.B(n_882),
.Y(n_1850)
);

AO31x2_ASAP7_75t_L g1851 ( 
.A1(n_1709),
.A2(n_1186),
.A3(n_1187),
.B(n_1020),
.Y(n_1851)
);

NOR2x1_ASAP7_75t_L g1852 ( 
.A(n_1679),
.B(n_1020),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1650),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1651),
.Y(n_1854)
);

OAI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1653),
.A2(n_1127),
.B1(n_1090),
.B2(n_1089),
.Y(n_1855)
);

AOI22xp5_ASAP7_75t_L g1856 ( 
.A1(n_1649),
.A2(n_1095),
.B1(n_1099),
.B2(n_1086),
.Y(n_1856)
);

BUFx6f_ASAP7_75t_L g1857 ( 
.A(n_1672),
.Y(n_1857)
);

OAI21x1_ASAP7_75t_L g1858 ( 
.A1(n_1656),
.A2(n_589),
.B(n_579),
.Y(n_1858)
);

AOI21xp5_ASAP7_75t_L g1859 ( 
.A1(n_1671),
.A2(n_1730),
.B(n_1728),
.Y(n_1859)
);

OAI21x1_ASAP7_75t_L g1860 ( 
.A1(n_1683),
.A2(n_592),
.B(n_591),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1701),
.B(n_14),
.Y(n_1861)
);

OAI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1731),
.A2(n_1143),
.B1(n_1108),
.B2(n_1121),
.Y(n_1862)
);

BUFx3_ASAP7_75t_L g1863 ( 
.A(n_1727),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1658),
.B(n_15),
.Y(n_1864)
);

OA21x2_ASAP7_75t_L g1865 ( 
.A1(n_1726),
.A2(n_1147),
.B(n_1105),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1706),
.B(n_16),
.Y(n_1866)
);

AOI21xp5_ASAP7_75t_L g1867 ( 
.A1(n_1733),
.A2(n_1187),
.B(n_1186),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1668),
.Y(n_1868)
);

A2O1A1Ixp33_ASAP7_75t_L g1869 ( 
.A1(n_1669),
.A2(n_1187),
.B(n_19),
.C(n_17),
.Y(n_1869)
);

OA21x2_ASAP7_75t_L g1870 ( 
.A1(n_1713),
.A2(n_599),
.B(n_596),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1698),
.B(n_18),
.Y(n_1871)
);

OAI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1734),
.A2(n_18),
.B(n_19),
.Y(n_1872)
);

AOI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1738),
.A2(n_601),
.B(n_600),
.Y(n_1873)
);

OAI21xp5_ASAP7_75t_L g1874 ( 
.A1(n_1739),
.A2(n_20),
.B(n_21),
.Y(n_1874)
);

OA21x2_ASAP7_75t_L g1875 ( 
.A1(n_1700),
.A2(n_605),
.B(n_602),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1667),
.B(n_22),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1727),
.Y(n_1877)
);

NOR2xp33_ASAP7_75t_L g1878 ( 
.A(n_1686),
.B(n_23),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1716),
.B(n_24),
.Y(n_1879)
);

AOI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1740),
.A2(n_608),
.B(n_607),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1673),
.B(n_24),
.Y(n_1881)
);

INVx2_ASAP7_75t_SL g1882 ( 
.A(n_1618),
.Y(n_1882)
);

OAI21x1_ASAP7_75t_L g1883 ( 
.A1(n_1674),
.A2(n_610),
.B(n_609),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1664),
.B(n_25),
.Y(n_1884)
);

OAI21x1_ASAP7_75t_L g1885 ( 
.A1(n_1741),
.A2(n_617),
.B(n_615),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_SL g1886 ( 
.A(n_1612),
.B(n_25),
.Y(n_1886)
);

AOI21xp5_ASAP7_75t_L g1887 ( 
.A1(n_1745),
.A2(n_619),
.B(n_618),
.Y(n_1887)
);

OAI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1748),
.A2(n_1754),
.B1(n_1757),
.B2(n_1752),
.Y(n_1888)
);

OAI21x1_ASAP7_75t_L g1889 ( 
.A1(n_1759),
.A2(n_622),
.B(n_621),
.Y(n_1889)
);

AOI21xp5_ASAP7_75t_L g1890 ( 
.A1(n_1760),
.A2(n_624),
.B(n_623),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1773),
.B(n_26),
.Y(n_1891)
);

AO22x2_ASAP7_75t_L g1892 ( 
.A1(n_1719),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1771),
.B(n_28),
.Y(n_1893)
);

AOI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1761),
.A2(n_626),
.B(n_625),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1717),
.B(n_1611),
.Y(n_1895)
);

AO31x2_ASAP7_75t_L g1896 ( 
.A1(n_1678),
.A2(n_628),
.A3(n_630),
.B(n_627),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1763),
.B(n_29),
.Y(n_1897)
);

AOI21xp5_ASAP7_75t_L g1898 ( 
.A1(n_1764),
.A2(n_1766),
.B(n_1666),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1605),
.B(n_1606),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1720),
.B(n_29),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_SL g1901 ( 
.A(n_1602),
.B(n_30),
.Y(n_1901)
);

AND2x6_ASAP7_75t_L g1902 ( 
.A(n_1863),
.B(n_1723),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1775),
.B(n_1681),
.Y(n_1903)
);

OA21x2_ASAP7_75t_L g1904 ( 
.A1(n_1779),
.A2(n_1721),
.B(n_1614),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1800),
.B(n_1613),
.Y(n_1905)
);

OAI21x1_ASAP7_75t_L g1906 ( 
.A1(n_1806),
.A2(n_1615),
.B(n_1710),
.Y(n_1906)
);

CKINVDCx20_ASAP7_75t_R g1907 ( 
.A(n_1812),
.Y(n_1907)
);

BUFx8_ASAP7_75t_L g1908 ( 
.A(n_1786),
.Y(n_1908)
);

OAI21x1_ASAP7_75t_L g1909 ( 
.A1(n_1808),
.A2(n_1693),
.B(n_1690),
.Y(n_1909)
);

OAI21x1_ASAP7_75t_L g1910 ( 
.A1(n_1816),
.A2(n_1694),
.B(n_1684),
.Y(n_1910)
);

NAND2x1p5_ASAP7_75t_L g1911 ( 
.A(n_1786),
.B(n_1791),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1777),
.Y(n_1912)
);

OAI21x1_ASAP7_75t_L g1913 ( 
.A1(n_1818),
.A2(n_633),
.B(n_632),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1795),
.Y(n_1914)
);

OR2x6_ASAP7_75t_L g1915 ( 
.A(n_1809),
.B(n_1791),
.Y(n_1915)
);

OAI21x1_ASAP7_75t_L g1916 ( 
.A1(n_1839),
.A2(n_1820),
.B(n_1787),
.Y(n_1916)
);

AOI22xp33_ASAP7_75t_L g1917 ( 
.A1(n_1807),
.A2(n_1629),
.B1(n_1737),
.B2(n_1729),
.Y(n_1917)
);

CKINVDCx5p33_ASAP7_75t_R g1918 ( 
.A(n_1840),
.Y(n_1918)
);

AOI21xp5_ASAP7_75t_L g1919 ( 
.A1(n_1797),
.A2(n_1776),
.B(n_1799),
.Y(n_1919)
);

AOI21xp5_ASAP7_75t_L g1920 ( 
.A1(n_1821),
.A2(n_1604),
.B(n_1744),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1794),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1832),
.Y(n_1922)
);

O2A1O1Ixp33_ASAP7_75t_L g1923 ( 
.A1(n_1793),
.A2(n_1749),
.B(n_1750),
.C(n_1747),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1866),
.Y(n_1924)
);

CKINVDCx5p33_ASAP7_75t_R g1925 ( 
.A(n_1857),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1807),
.B(n_1751),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1814),
.B(n_30),
.Y(n_1927)
);

OAI21x1_ASAP7_75t_SL g1928 ( 
.A1(n_1872),
.A2(n_33),
.B(n_32),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1842),
.Y(n_1929)
);

OAI21x1_ASAP7_75t_L g1930 ( 
.A1(n_1849),
.A2(n_637),
.B(n_634),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1829),
.B(n_1810),
.Y(n_1931)
);

OAI21xp5_ASAP7_75t_L g1932 ( 
.A1(n_1774),
.A2(n_1765),
.B(n_1758),
.Y(n_1932)
);

OR2x2_ASAP7_75t_L g1933 ( 
.A(n_1778),
.B(n_1767),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_SL g1934 ( 
.A(n_1868),
.B(n_1824),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1836),
.Y(n_1935)
);

AOI21xp5_ASAP7_75t_R g1936 ( 
.A1(n_1888),
.A2(n_31),
.B(n_32),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1847),
.Y(n_1937)
);

AND2x6_ASAP7_75t_L g1938 ( 
.A(n_1877),
.B(n_638),
.Y(n_1938)
);

AO21x2_ASAP7_75t_L g1939 ( 
.A1(n_1790),
.A2(n_640),
.B(n_639),
.Y(n_1939)
);

INVx3_ASAP7_75t_L g1940 ( 
.A(n_1804),
.Y(n_1940)
);

OAI21x1_ASAP7_75t_L g1941 ( 
.A1(n_1858),
.A2(n_644),
.B(n_643),
.Y(n_1941)
);

AOI22xp5_ASAP7_75t_L g1942 ( 
.A1(n_1876),
.A2(n_37),
.B1(n_34),
.B2(n_36),
.Y(n_1942)
);

OR2x2_ASAP7_75t_L g1943 ( 
.A(n_1827),
.B(n_36),
.Y(n_1943)
);

OAI21x1_ASAP7_75t_L g1944 ( 
.A1(n_1883),
.A2(n_647),
.B(n_646),
.Y(n_1944)
);

OAI21x1_ASAP7_75t_L g1945 ( 
.A1(n_1885),
.A2(n_649),
.B(n_648),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1884),
.Y(n_1946)
);

NAND3xp33_ASAP7_75t_L g1947 ( 
.A(n_1869),
.B(n_39),
.C(n_40),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_SL g1948 ( 
.A(n_1813),
.B(n_39),
.Y(n_1948)
);

AOI22xp33_ASAP7_75t_L g1949 ( 
.A1(n_1817),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1853),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1854),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1783),
.B(n_43),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1803),
.B(n_44),
.Y(n_1953)
);

O2A1O1Ixp33_ASAP7_75t_L g1954 ( 
.A1(n_1780),
.A2(n_47),
.B(n_45),
.C(n_46),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1882),
.B(n_46),
.Y(n_1955)
);

HB1xp67_ASAP7_75t_L g1956 ( 
.A(n_1864),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1831),
.B(n_47),
.Y(n_1957)
);

AND2x4_ASAP7_75t_L g1958 ( 
.A(n_1844),
.B(n_651),
.Y(n_1958)
);

AOI22xp33_ASAP7_75t_L g1959 ( 
.A1(n_1828),
.A2(n_51),
.B1(n_48),
.B2(n_49),
.Y(n_1959)
);

INVx3_ASAP7_75t_L g1960 ( 
.A(n_1843),
.Y(n_1960)
);

OR2x2_ASAP7_75t_L g1961 ( 
.A(n_1899),
.B(n_48),
.Y(n_1961)
);

AOI222xp33_ASAP7_75t_L g1962 ( 
.A1(n_1845),
.A2(n_53),
.B1(n_55),
.B2(n_51),
.C1(n_52),
.C2(n_54),
.Y(n_1962)
);

OAI21x1_ASAP7_75t_L g1963 ( 
.A1(n_1889),
.A2(n_653),
.B(n_652),
.Y(n_1963)
);

OAI22xp5_ASAP7_75t_L g1964 ( 
.A1(n_1805),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_1964)
);

HB1xp67_ASAP7_75t_L g1965 ( 
.A(n_1833),
.Y(n_1965)
);

HB1xp67_ASAP7_75t_L g1966 ( 
.A(n_1861),
.Y(n_1966)
);

OAI22xp5_ASAP7_75t_L g1967 ( 
.A1(n_1859),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_1967)
);

A2O1A1Ixp33_ASAP7_75t_L g1968 ( 
.A1(n_1878),
.A2(n_1898),
.B(n_1789),
.C(n_1874),
.Y(n_1968)
);

NOR3xp33_ASAP7_75t_L g1969 ( 
.A(n_1886),
.B(n_57),
.C(n_59),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1879),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1900),
.Y(n_1971)
);

OAI21x1_ASAP7_75t_L g1972 ( 
.A1(n_1860),
.A2(n_656),
.B(n_655),
.Y(n_1972)
);

NOR2xp67_ASAP7_75t_L g1973 ( 
.A(n_1819),
.B(n_1835),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1892),
.B(n_59),
.Y(n_1974)
);

INVxp67_ASAP7_75t_L g1975 ( 
.A(n_1871),
.Y(n_1975)
);

HB1xp67_ASAP7_75t_L g1976 ( 
.A(n_1895),
.Y(n_1976)
);

OAI21x1_ASAP7_75t_L g1977 ( 
.A1(n_1867),
.A2(n_661),
.B(n_659),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1796),
.Y(n_1978)
);

AND2x4_ASAP7_75t_L g1979 ( 
.A(n_1852),
.B(n_663),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1796),
.Y(n_1980)
);

OAI21x1_ASAP7_75t_L g1981 ( 
.A1(n_1873),
.A2(n_667),
.B(n_665),
.Y(n_1981)
);

AOI222xp33_ASAP7_75t_L g1982 ( 
.A1(n_1892),
.A2(n_63),
.B1(n_65),
.B2(n_61),
.C1(n_62),
.C2(n_64),
.Y(n_1982)
);

BUFx8_ASAP7_75t_L g1983 ( 
.A(n_1823),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1891),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1870),
.Y(n_1985)
);

BUFx3_ASAP7_75t_L g1986 ( 
.A(n_1893),
.Y(n_1986)
);

INVxp33_ASAP7_75t_SL g1987 ( 
.A(n_1834),
.Y(n_1987)
);

BUFx12f_ASAP7_75t_L g1988 ( 
.A(n_1802),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1897),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1881),
.B(n_64),
.Y(n_1990)
);

OAI21xp5_ASAP7_75t_L g1991 ( 
.A1(n_1801),
.A2(n_65),
.B(n_66),
.Y(n_1991)
);

NAND2x1p5_ASAP7_75t_L g1992 ( 
.A(n_1901),
.B(n_668),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1784),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1851),
.Y(n_1994)
);

HB1xp67_ASAP7_75t_L g1995 ( 
.A(n_1875),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1848),
.B(n_66),
.Y(n_1996)
);

INVx3_ASAP7_75t_L g1997 ( 
.A(n_1865),
.Y(n_1997)
);

O2A1O1Ixp33_ASAP7_75t_SL g1998 ( 
.A1(n_1880),
.A2(n_69),
.B(n_67),
.C(n_68),
.Y(n_1998)
);

INVx1_ASAP7_75t_SL g1999 ( 
.A(n_1798),
.Y(n_1999)
);

INVx3_ASAP7_75t_L g2000 ( 
.A(n_1851),
.Y(n_2000)
);

NOR2xp33_ASAP7_75t_L g2001 ( 
.A(n_1856),
.B(n_1862),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1785),
.Y(n_2002)
);

OAI21x1_ASAP7_75t_SL g2003 ( 
.A1(n_1887),
.A2(n_70),
.B(n_69),
.Y(n_2003)
);

AO21x2_ASAP7_75t_L g2004 ( 
.A1(n_1781),
.A2(n_672),
.B(n_671),
.Y(n_2004)
);

NAND2xp33_ASAP7_75t_R g2005 ( 
.A(n_1890),
.B(n_673),
.Y(n_2005)
);

NAND2x1p5_ASAP7_75t_L g2006 ( 
.A(n_1894),
.B(n_674),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1855),
.B(n_67),
.Y(n_2007)
);

OR2x6_ASAP7_75t_L g2008 ( 
.A(n_1788),
.B(n_70),
.Y(n_2008)
);

AND2x4_ASAP7_75t_L g2009 ( 
.A(n_1811),
.B(n_678),
.Y(n_2009)
);

OAI21xp5_ASAP7_75t_L g2010 ( 
.A1(n_1822),
.A2(n_71),
.B(n_72),
.Y(n_2010)
);

OAI21xp5_ASAP7_75t_L g2011 ( 
.A1(n_1825),
.A2(n_72),
.B(n_73),
.Y(n_2011)
);

OA21x2_ASAP7_75t_L g2012 ( 
.A1(n_1792),
.A2(n_1850),
.B(n_1830),
.Y(n_2012)
);

HB1xp67_ASAP7_75t_L g2013 ( 
.A(n_1792),
.Y(n_2013)
);

OA21x2_ASAP7_75t_L g2014 ( 
.A1(n_1850),
.A2(n_680),
.B(n_679),
.Y(n_2014)
);

O2A1O1Ixp33_ASAP7_75t_L g2015 ( 
.A1(n_1826),
.A2(n_75),
.B(n_73),
.C(n_74),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1896),
.Y(n_2016)
);

NOR2xp67_ASAP7_75t_L g2017 ( 
.A(n_1815),
.B(n_681),
.Y(n_2017)
);

CKINVDCx5p33_ASAP7_75t_R g2018 ( 
.A(n_1838),
.Y(n_2018)
);

OAI21xp5_ASAP7_75t_L g2019 ( 
.A1(n_1841),
.A2(n_74),
.B(n_75),
.Y(n_2019)
);

A2O1A1Ixp33_ASAP7_75t_L g2020 ( 
.A1(n_1846),
.A2(n_79),
.B(n_80),
.C(n_77),
.Y(n_2020)
);

AND2x4_ASAP7_75t_L g2021 ( 
.A(n_1896),
.B(n_685),
.Y(n_2021)
);

OA21x2_ASAP7_75t_L g2022 ( 
.A1(n_1779),
.A2(n_688),
.B(n_687),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1795),
.Y(n_2023)
);

INVx8_ASAP7_75t_L g2024 ( 
.A(n_1786),
.Y(n_2024)
);

AO31x2_ASAP7_75t_L g2025 ( 
.A1(n_1837),
.A2(n_690),
.A3(n_691),
.B(n_689),
.Y(n_2025)
);

INVx4_ASAP7_75t_L g2026 ( 
.A(n_1786),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_R g2027 ( 
.A(n_1775),
.B(n_692),
.Y(n_2027)
);

NAND2x1p5_ASAP7_75t_L g2028 ( 
.A(n_1786),
.B(n_693),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1777),
.Y(n_2029)
);

OAI21x1_ASAP7_75t_L g2030 ( 
.A1(n_1806),
.A2(n_696),
.B(n_694),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1775),
.B(n_76),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1775),
.B(n_81),
.Y(n_2032)
);

NOR2x1_ASAP7_75t_SL g2033 ( 
.A(n_1782),
.B(n_83),
.Y(n_2033)
);

OAI21x1_ASAP7_75t_L g2034 ( 
.A1(n_1916),
.A2(n_698),
.B(n_697),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1912),
.Y(n_2035)
);

OAI21x1_ASAP7_75t_L g2036 ( 
.A1(n_2000),
.A2(n_701),
.B(n_700),
.Y(n_2036)
);

OR2x6_ASAP7_75t_L g2037 ( 
.A(n_2024),
.B(n_702),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_2029),
.Y(n_2038)
);

OAI21xp33_ASAP7_75t_SL g2039 ( 
.A1(n_2001),
.A2(n_83),
.B(n_84),
.Y(n_2039)
);

CKINVDCx14_ASAP7_75t_R g2040 ( 
.A(n_1925),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_1927),
.B(n_86),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1914),
.Y(n_2042)
);

BUFx2_ASAP7_75t_L g2043 ( 
.A(n_1918),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2023),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1935),
.Y(n_2045)
);

AOI21xp5_ASAP7_75t_SL g2046 ( 
.A1(n_1968),
.A2(n_87),
.B(n_88),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1937),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_1952),
.B(n_89),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1950),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1951),
.Y(n_2050)
);

OAI21xp5_ASAP7_75t_L g2051 ( 
.A1(n_1953),
.A2(n_90),
.B(n_91),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_1970),
.Y(n_2052)
);

INVx3_ASAP7_75t_L g2053 ( 
.A(n_1908),
.Y(n_2053)
);

OAI21x1_ASAP7_75t_L g2054 ( 
.A1(n_1978),
.A2(n_707),
.B(n_705),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1946),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1922),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1965),
.Y(n_2057)
);

INVx3_ASAP7_75t_L g2058 ( 
.A(n_2026),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1924),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1956),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1929),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_1974),
.B(n_91),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1971),
.Y(n_2063)
);

INVx6_ASAP7_75t_L g2064 ( 
.A(n_1983),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1984),
.Y(n_2065)
);

OA21x2_ASAP7_75t_L g2066 ( 
.A1(n_2016),
.A2(n_1994),
.B(n_1980),
.Y(n_2066)
);

BUFx6f_ASAP7_75t_L g2067 ( 
.A(n_1911),
.Y(n_2067)
);

BUFx2_ASAP7_75t_L g2068 ( 
.A(n_1921),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1989),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_2002),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1905),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1976),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1966),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1904),
.Y(n_2074)
);

BUFx2_ASAP7_75t_L g2075 ( 
.A(n_2013),
.Y(n_2075)
);

INVx2_ASAP7_75t_SL g2076 ( 
.A(n_1940),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1934),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1960),
.Y(n_2078)
);

INVx3_ASAP7_75t_L g2079 ( 
.A(n_1915),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_1997),
.Y(n_2080)
);

HB1xp67_ASAP7_75t_L g2081 ( 
.A(n_1986),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1961),
.Y(n_2082)
);

INVx2_ASAP7_75t_L g2083 ( 
.A(n_1993),
.Y(n_2083)
);

BUFx2_ASAP7_75t_SL g2084 ( 
.A(n_1973),
.Y(n_2084)
);

OAI21x1_ASAP7_75t_L g2085 ( 
.A1(n_2030),
.A2(n_710),
.B(n_709),
.Y(n_2085)
);

INVx3_ASAP7_75t_L g2086 ( 
.A(n_1915),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1958),
.Y(n_2087)
);

AOI21x1_ASAP7_75t_L g2088 ( 
.A1(n_1995),
.A2(n_712),
.B(n_711),
.Y(n_2088)
);

HB1xp67_ASAP7_75t_L g2089 ( 
.A(n_1931),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2033),
.Y(n_2090)
);

HB1xp67_ASAP7_75t_L g2091 ( 
.A(n_1975),
.Y(n_2091)
);

AO21x1_ASAP7_75t_SL g2092 ( 
.A1(n_1991),
.A2(n_92),
.B(n_93),
.Y(n_2092)
);

INVx1_ASAP7_75t_SL g2093 ( 
.A(n_2027),
.Y(n_2093)
);

NOR2xp33_ASAP7_75t_L g2094 ( 
.A(n_1987),
.B(n_94),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1906),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_2031),
.B(n_95),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1943),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1990),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_2004),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2032),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_1928),
.Y(n_2101)
);

AND2x4_ASAP7_75t_L g2102 ( 
.A(n_1902),
.B(n_96),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_2021),
.Y(n_2103)
);

OAI21x1_ASAP7_75t_L g2104 ( 
.A1(n_1985),
.A2(n_715),
.B(n_713),
.Y(n_2104)
);

INVxp67_ASAP7_75t_L g2105 ( 
.A(n_1903),
.Y(n_2105)
);

OR2x2_ASAP7_75t_L g2106 ( 
.A(n_1933),
.B(n_97),
.Y(n_2106)
);

AOI22xp33_ASAP7_75t_SL g2107 ( 
.A1(n_1907),
.A2(n_100),
.B1(n_101),
.B2(n_98),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1919),
.Y(n_2108)
);

BUFx2_ASAP7_75t_L g2109 ( 
.A(n_1988),
.Y(n_2109)
);

INVx2_ASAP7_75t_SL g2110 ( 
.A(n_1955),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1938),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_2028),
.Y(n_2112)
);

A2O1A1Ixp33_ASAP7_75t_L g2113 ( 
.A1(n_1923),
.A2(n_1920),
.B(n_1932),
.C(n_2015),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1938),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_2012),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_2007),
.B(n_97),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1938),
.Y(n_2117)
);

INVx3_ASAP7_75t_L g2118 ( 
.A(n_1902),
.Y(n_2118)
);

AOI22xp33_ASAP7_75t_SL g2119 ( 
.A1(n_1936),
.A2(n_103),
.B1(n_104),
.B2(n_101),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1967),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1954),
.Y(n_2121)
);

XOR2xp5_ASAP7_75t_L g2122 ( 
.A(n_2040),
.B(n_2018),
.Y(n_2122)
);

AND2x4_ASAP7_75t_L g2123 ( 
.A(n_2081),
.B(n_1926),
.Y(n_2123)
);

INVxp67_ASAP7_75t_L g2124 ( 
.A(n_2089),
.Y(n_2124)
);

CKINVDCx5p33_ASAP7_75t_R g2125 ( 
.A(n_2064),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2062),
.B(n_1982),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2057),
.Y(n_2127)
);

HB1xp67_ASAP7_75t_L g2128 ( 
.A(n_2072),
.Y(n_2128)
);

BUFx3_ASAP7_75t_L g2129 ( 
.A(n_2043),
.Y(n_2129)
);

NAND2xp33_ASAP7_75t_R g2130 ( 
.A(n_2053),
.B(n_2102),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_2071),
.B(n_1962),
.Y(n_2131)
);

AND2x4_ASAP7_75t_L g2132 ( 
.A(n_2079),
.B(n_1902),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_2050),
.Y(n_2133)
);

XOR2xp5_ASAP7_75t_L g2134 ( 
.A(n_2106),
.B(n_1917),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_2105),
.B(n_1942),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_2045),
.Y(n_2136)
);

BUFx3_ASAP7_75t_L g2137 ( 
.A(n_2064),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_2047),
.Y(n_2138)
);

NAND2xp33_ASAP7_75t_R g2139 ( 
.A(n_2109),
.B(n_1957),
.Y(n_2139)
);

XNOR2xp5_ASAP7_75t_L g2140 ( 
.A(n_2093),
.B(n_1949),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_2091),
.B(n_1959),
.Y(n_2141)
);

NAND2xp33_ASAP7_75t_R g2142 ( 
.A(n_2118),
.B(n_2008),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2035),
.Y(n_2143)
);

BUFx3_ASAP7_75t_L g2144 ( 
.A(n_2076),
.Y(n_2144)
);

INVxp67_ASAP7_75t_L g2145 ( 
.A(n_2078),
.Y(n_2145)
);

BUFx3_ASAP7_75t_L g2146 ( 
.A(n_2058),
.Y(n_2146)
);

NAND2xp33_ASAP7_75t_R g2147 ( 
.A(n_2037),
.B(n_2008),
.Y(n_2147)
);

NAND2xp33_ASAP7_75t_R g2148 ( 
.A(n_2037),
.B(n_1996),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2038),
.Y(n_2149)
);

NOR2xp33_ASAP7_75t_R g2150 ( 
.A(n_2086),
.B(n_2005),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2098),
.B(n_1969),
.Y(n_2151)
);

NAND2xp33_ASAP7_75t_R g2152 ( 
.A(n_2094),
.B(n_1979),
.Y(n_2152)
);

BUFx3_ASAP7_75t_L g2153 ( 
.A(n_2067),
.Y(n_2153)
);

NOR2xp33_ASAP7_75t_R g2154 ( 
.A(n_2110),
.B(n_2009),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_2052),
.B(n_1948),
.Y(n_2155)
);

BUFx3_ASAP7_75t_L g2156 ( 
.A(n_2060),
.Y(n_2156)
);

NOR2xp33_ASAP7_75t_R g2157 ( 
.A(n_2111),
.B(n_2114),
.Y(n_2157)
);

AND2x4_ASAP7_75t_L g2158 ( 
.A(n_2103),
.B(n_1999),
.Y(n_2158)
);

AND2x4_ASAP7_75t_L g2159 ( 
.A(n_2087),
.B(n_2117),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_2055),
.B(n_1964),
.Y(n_2160)
);

XNOR2xp5_ASAP7_75t_L g2161 ( 
.A(n_2041),
.B(n_1947),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_2049),
.Y(n_2162)
);

OR2x6_ASAP7_75t_L g2163 ( 
.A(n_2084),
.B(n_1992),
.Y(n_2163)
);

AND2x4_ASAP7_75t_L g2164 ( 
.A(n_2073),
.B(n_1909),
.Y(n_2164)
);

OR2x6_ASAP7_75t_L g2165 ( 
.A(n_2046),
.B(n_2003),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_2082),
.B(n_2010),
.Y(n_2166)
);

NOR2xp33_ASAP7_75t_R g2167 ( 
.A(n_2100),
.B(n_2097),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2056),
.Y(n_2168)
);

AND2x4_ASAP7_75t_L g2169 ( 
.A(n_2112),
.B(n_2020),
.Y(n_2169)
);

NOR2xp33_ASAP7_75t_R g2170 ( 
.A(n_2090),
.B(n_98),
.Y(n_2170)
);

AND2x4_ASAP7_75t_L g2171 ( 
.A(n_2059),
.B(n_2061),
.Y(n_2171)
);

NOR2xp33_ASAP7_75t_R g2172 ( 
.A(n_2048),
.B(n_105),
.Y(n_2172)
);

AOI22xp33_ASAP7_75t_L g2173 ( 
.A1(n_2126),
.A2(n_2092),
.B1(n_2150),
.B2(n_2131),
.Y(n_2173)
);

AND2x2_ASAP7_75t_L g2174 ( 
.A(n_2156),
.B(n_2116),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2128),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_2136),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2143),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_2129),
.B(n_2075),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_2138),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_2127),
.B(n_2075),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_2166),
.B(n_2077),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_2162),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2149),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2168),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2171),
.Y(n_2185)
);

OR2x6_ASAP7_75t_L g2186 ( 
.A(n_2163),
.B(n_2132),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2133),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2164),
.Y(n_2188)
);

HB1xp67_ASAP7_75t_L g2189 ( 
.A(n_2123),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2155),
.Y(n_2190)
);

NOR2x1_ASAP7_75t_L g2191 ( 
.A(n_2144),
.B(n_2113),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_2167),
.B(n_2096),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2159),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_2146),
.B(n_2068),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_2151),
.B(n_2063),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2145),
.B(n_2065),
.Y(n_2196)
);

OR2x2_ASAP7_75t_L g2197 ( 
.A(n_2135),
.B(n_2068),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2158),
.Y(n_2198)
);

OR2x2_ASAP7_75t_L g2199 ( 
.A(n_2141),
.B(n_2069),
.Y(n_2199)
);

OR2x2_ASAP7_75t_L g2200 ( 
.A(n_2160),
.B(n_2083),
.Y(n_2200)
);

OR2x2_ASAP7_75t_L g2201 ( 
.A(n_2134),
.B(n_2080),
.Y(n_2201)
);

CKINVDCx11_ASAP7_75t_R g2202 ( 
.A(n_2137),
.Y(n_2202)
);

BUFx2_ASAP7_75t_L g2203 ( 
.A(n_2157),
.Y(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_2172),
.B(n_2070),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2169),
.Y(n_2205)
);

NOR2x1_ASAP7_75t_L g2206 ( 
.A(n_2122),
.B(n_2121),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2153),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_2161),
.B(n_2108),
.Y(n_2208)
);

AOI22xp33_ASAP7_75t_L g2209 ( 
.A1(n_2140),
.A2(n_2119),
.B1(n_2051),
.B2(n_2120),
.Y(n_2209)
);

INVxp67_ASAP7_75t_L g2210 ( 
.A(n_2139),
.Y(n_2210)
);

AND2x4_ASAP7_75t_L g2211 ( 
.A(n_2125),
.B(n_2042),
.Y(n_2211)
);

AOI22xp33_ASAP7_75t_L g2212 ( 
.A1(n_2154),
.A2(n_2107),
.B1(n_2011),
.B2(n_2019),
.Y(n_2212)
);

INVxp67_ASAP7_75t_SL g2213 ( 
.A(n_2148),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_2165),
.Y(n_2214)
);

AND2x4_ASAP7_75t_L g2215 ( 
.A(n_2165),
.B(n_2044),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2170),
.Y(n_2216)
);

INVxp67_ASAP7_75t_L g2217 ( 
.A(n_2130),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_2142),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_2147),
.B(n_2101),
.Y(n_2219)
);

AND2x4_ASAP7_75t_L g2220 ( 
.A(n_2152),
.B(n_2074),
.Y(n_2220)
);

AND2x4_ASAP7_75t_L g2221 ( 
.A(n_2156),
.B(n_2095),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2124),
.B(n_2039),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2177),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_2176),
.Y(n_2224)
);

BUFx2_ASAP7_75t_L g2225 ( 
.A(n_2188),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2183),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_2179),
.Y(n_2227)
);

AND2x4_ASAP7_75t_SL g2228 ( 
.A(n_2186),
.B(n_2099),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_2178),
.B(n_2174),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_2181),
.B(n_2115),
.Y(n_2230)
);

AOI22xp5_ASAP7_75t_L g2231 ( 
.A1(n_2212),
.A2(n_1998),
.B1(n_2017),
.B2(n_1939),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2190),
.B(n_2025),
.Y(n_2232)
);

AND2x2_ASAP7_75t_L g2233 ( 
.A(n_2194),
.B(n_2189),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_2182),
.Y(n_2234)
);

AND2x2_ASAP7_75t_L g2235 ( 
.A(n_2180),
.B(n_2066),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_2175),
.B(n_2066),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2184),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_2208),
.B(n_2034),
.Y(n_2238)
);

AND2x2_ASAP7_75t_L g2239 ( 
.A(n_2213),
.B(n_2025),
.Y(n_2239)
);

HB1xp67_ASAP7_75t_L g2240 ( 
.A(n_2197),
.Y(n_2240)
);

AND2x2_ASAP7_75t_L g2241 ( 
.A(n_2203),
.B(n_1910),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_2187),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_2185),
.Y(n_2243)
);

BUFx3_ASAP7_75t_L g2244 ( 
.A(n_2202),
.Y(n_2244)
);

AND2x2_ASAP7_75t_L g2245 ( 
.A(n_2203),
.B(n_2088),
.Y(n_2245)
);

HB1xp67_ASAP7_75t_L g2246 ( 
.A(n_2222),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2199),
.Y(n_2247)
);

AND2x4_ASAP7_75t_L g2248 ( 
.A(n_2221),
.B(n_2036),
.Y(n_2248)
);

NOR2xp33_ASAP7_75t_R g2249 ( 
.A(n_2216),
.B(n_105),
.Y(n_2249)
);

NOR2xp33_ASAP7_75t_L g2250 ( 
.A(n_2206),
.B(n_106),
.Y(n_2250)
);

BUFx2_ASAP7_75t_L g2251 ( 
.A(n_2214),
.Y(n_2251)
);

AND2x2_ASAP7_75t_L g2252 ( 
.A(n_2210),
.B(n_2085),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_2198),
.Y(n_2253)
);

AND2x4_ASAP7_75t_L g2254 ( 
.A(n_2205),
.B(n_2054),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_2192),
.B(n_1913),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2200),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2196),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_2193),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_2217),
.B(n_1945),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2195),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_2218),
.B(n_1963),
.Y(n_2261)
);

AND2x2_ASAP7_75t_SL g2262 ( 
.A(n_2220),
.B(n_2014),
.Y(n_2262)
);

OAI31xp33_ASAP7_75t_L g2263 ( 
.A1(n_2209),
.A2(n_2006),
.A3(n_110),
.B(n_107),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2201),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2186),
.B(n_1972),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2215),
.Y(n_2266)
);

OAI211xp5_ASAP7_75t_L g2267 ( 
.A1(n_2173),
.A2(n_114),
.B(n_111),
.C(n_113),
.Y(n_2267)
);

BUFx3_ASAP7_75t_L g2268 ( 
.A(n_2207),
.Y(n_2268)
);

AOI22xp5_ASAP7_75t_L g2269 ( 
.A1(n_2204),
.A2(n_2022),
.B1(n_2104),
.B2(n_1981),
.Y(n_2269)
);

INVx3_ASAP7_75t_L g2270 ( 
.A(n_2211),
.Y(n_2270)
);

AND2x4_ASAP7_75t_L g2271 ( 
.A(n_2178),
.B(n_1944),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2181),
.B(n_115),
.Y(n_2272)
);

OR2x2_ASAP7_75t_L g2273 ( 
.A(n_2197),
.B(n_115),
.Y(n_2273)
);

AO21x2_ASAP7_75t_L g2274 ( 
.A1(n_2219),
.A2(n_1930),
.B(n_1941),
.Y(n_2274)
);

OAI22xp5_ASAP7_75t_L g2275 ( 
.A1(n_2209),
.A2(n_118),
.B1(n_116),
.B2(n_117),
.Y(n_2275)
);

OR2x2_ASAP7_75t_L g2276 ( 
.A(n_2197),
.B(n_116),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_2176),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2181),
.B(n_118),
.Y(n_2278)
);

AND2x2_ASAP7_75t_L g2279 ( 
.A(n_2178),
.B(n_119),
.Y(n_2279)
);

OR2x2_ASAP7_75t_L g2280 ( 
.A(n_2197),
.B(n_119),
.Y(n_2280)
);

OR2x2_ASAP7_75t_L g2281 ( 
.A(n_2197),
.B(n_121),
.Y(n_2281)
);

OR2x2_ASAP7_75t_L g2282 ( 
.A(n_2197),
.B(n_122),
.Y(n_2282)
);

HB1xp67_ASAP7_75t_L g2283 ( 
.A(n_2175),
.Y(n_2283)
);

OAI21x1_ASAP7_75t_L g2284 ( 
.A1(n_2191),
.A2(n_1977),
.B(n_122),
.Y(n_2284)
);

AND2x2_ASAP7_75t_L g2285 ( 
.A(n_2178),
.B(n_123),
.Y(n_2285)
);

OR2x2_ASAP7_75t_L g2286 ( 
.A(n_2240),
.B(n_123),
.Y(n_2286)
);

INVx2_ASAP7_75t_SL g2287 ( 
.A(n_2244),
.Y(n_2287)
);

INVx2_ASAP7_75t_SL g2288 ( 
.A(n_2233),
.Y(n_2288)
);

NOR2xp33_ASAP7_75t_SL g2289 ( 
.A(n_2250),
.B(n_2268),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_2229),
.B(n_2246),
.Y(n_2290)
);

INVxp67_ASAP7_75t_L g2291 ( 
.A(n_2283),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2223),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_2270),
.B(n_124),
.Y(n_2293)
);

AOI21x1_ASAP7_75t_SL g2294 ( 
.A1(n_2252),
.A2(n_124),
.B(n_125),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_2225),
.B(n_125),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2226),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_2242),
.Y(n_2297)
);

OR2x2_ASAP7_75t_L g2298 ( 
.A(n_2230),
.B(n_126),
.Y(n_2298)
);

OR2x2_ASAP7_75t_L g2299 ( 
.A(n_2256),
.B(n_126),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_2224),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2257),
.B(n_127),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2260),
.B(n_127),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2237),
.Y(n_2303)
);

NAND2x1p5_ASAP7_75t_L g2304 ( 
.A(n_2279),
.B(n_128),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2247),
.Y(n_2305)
);

BUFx3_ASAP7_75t_L g2306 ( 
.A(n_2251),
.Y(n_2306)
);

AND2x2_ASAP7_75t_L g2307 ( 
.A(n_2241),
.B(n_128),
.Y(n_2307)
);

INVx4_ASAP7_75t_L g2308 ( 
.A(n_2285),
.Y(n_2308)
);

AND2x4_ASAP7_75t_SL g2309 ( 
.A(n_2266),
.B(n_129),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2264),
.Y(n_2310)
);

AND2x2_ASAP7_75t_L g2311 ( 
.A(n_2238),
.B(n_2251),
.Y(n_2311)
);

OR2x2_ASAP7_75t_L g2312 ( 
.A(n_2235),
.B(n_129),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2253),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2258),
.Y(n_2314)
);

HB1xp67_ASAP7_75t_L g2315 ( 
.A(n_2245),
.Y(n_2315)
);

AND2x2_ASAP7_75t_L g2316 ( 
.A(n_2255),
.B(n_130),
.Y(n_2316)
);

OR2x2_ASAP7_75t_L g2317 ( 
.A(n_2273),
.B(n_2276),
.Y(n_2317)
);

INVx2_ASAP7_75t_SL g2318 ( 
.A(n_2280),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2239),
.B(n_130),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2243),
.Y(n_2320)
);

INVx2_ASAP7_75t_L g2321 ( 
.A(n_2227),
.Y(n_2321)
);

INVx2_ASAP7_75t_SL g2322 ( 
.A(n_2281),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2234),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2277),
.Y(n_2324)
);

BUFx3_ASAP7_75t_L g2325 ( 
.A(n_2282),
.Y(n_2325)
);

AND2x6_ASAP7_75t_SL g2326 ( 
.A(n_2272),
.B(n_131),
.Y(n_2326)
);

INVx2_ASAP7_75t_SL g2327 ( 
.A(n_2249),
.Y(n_2327)
);

AND2x4_ASAP7_75t_L g2328 ( 
.A(n_2228),
.B(n_132),
.Y(n_2328)
);

OA21x2_ASAP7_75t_L g2329 ( 
.A1(n_2232),
.A2(n_133),
.B(n_134),
.Y(n_2329)
);

NAND2x1p5_ASAP7_75t_L g2330 ( 
.A(n_2265),
.B(n_133),
.Y(n_2330)
);

AND2x4_ASAP7_75t_L g2331 ( 
.A(n_2261),
.B(n_135),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_2278),
.B(n_136),
.Y(n_2332)
);

OR2x2_ASAP7_75t_L g2333 ( 
.A(n_2259),
.B(n_137),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2254),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_2271),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_2248),
.B(n_138),
.Y(n_2336)
);

NAND2x1p5_ASAP7_75t_L g2337 ( 
.A(n_2262),
.B(n_139),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2231),
.B(n_139),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2274),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2284),
.Y(n_2340)
);

AND2x4_ASAP7_75t_L g2341 ( 
.A(n_2269),
.B(n_141),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_2275),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_2267),
.B(n_142),
.Y(n_2343)
);

AND2x2_ASAP7_75t_L g2344 ( 
.A(n_2263),
.B(n_143),
.Y(n_2344)
);

AND2x2_ASAP7_75t_L g2345 ( 
.A(n_2229),
.B(n_144),
.Y(n_2345)
);

OR2x6_ASAP7_75t_L g2346 ( 
.A(n_2244),
.B(n_144),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2283),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2246),
.B(n_146),
.Y(n_2348)
);

OR2x2_ASAP7_75t_L g2349 ( 
.A(n_2240),
.B(n_147),
.Y(n_2349)
);

OR2x2_ASAP7_75t_L g2350 ( 
.A(n_2240),
.B(n_147),
.Y(n_2350)
);

HB1xp67_ASAP7_75t_L g2351 ( 
.A(n_2246),
.Y(n_2351)
);

INVxp67_ASAP7_75t_SL g2352 ( 
.A(n_2246),
.Y(n_2352)
);

AND2x2_ASAP7_75t_L g2353 ( 
.A(n_2229),
.B(n_148),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_2236),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2283),
.Y(n_2355)
);

NOR2x1_ASAP7_75t_L g2356 ( 
.A(n_2244),
.B(n_149),
.Y(n_2356)
);

NOR2xp33_ASAP7_75t_L g2357 ( 
.A(n_2244),
.B(n_150),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2283),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2283),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2283),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2283),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2283),
.Y(n_2362)
);

AND3x2_ASAP7_75t_L g2363 ( 
.A(n_2250),
.B(n_151),
.C(n_152),
.Y(n_2363)
);

HB1xp67_ASAP7_75t_L g2364 ( 
.A(n_2246),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2283),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2283),
.Y(n_2366)
);

HB1xp67_ASAP7_75t_L g2367 ( 
.A(n_2246),
.Y(n_2367)
);

NOR2xp67_ASAP7_75t_L g2368 ( 
.A(n_2246),
.B(n_152),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2283),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2283),
.Y(n_2370)
);

AND2x2_ASAP7_75t_L g2371 ( 
.A(n_2229),
.B(n_153),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2236),
.Y(n_2372)
);

NAND2xp33_ASAP7_75t_SL g2373 ( 
.A(n_2295),
.B(n_154),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_2352),
.B(n_155),
.Y(n_2374)
);

CKINVDCx5p33_ASAP7_75t_R g2375 ( 
.A(n_2287),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_SL g2376 ( 
.A(n_2306),
.B(n_157),
.Y(n_2376)
);

AO221x2_ASAP7_75t_L g2377 ( 
.A1(n_2319),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.C(n_161),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2290),
.B(n_158),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2351),
.B(n_160),
.Y(n_2379)
);

AO221x2_ASAP7_75t_L g2380 ( 
.A1(n_2348),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.C(n_165),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2364),
.B(n_163),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2292),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2367),
.B(n_164),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2291),
.B(n_167),
.Y(n_2384)
);

INVxp67_ASAP7_75t_SL g2385 ( 
.A(n_2368),
.Y(n_2385)
);

CKINVDCx16_ASAP7_75t_R g2386 ( 
.A(n_2289),
.Y(n_2386)
);

NOR2xp33_ASAP7_75t_L g2387 ( 
.A(n_2326),
.B(n_2308),
.Y(n_2387)
);

NOR2xp33_ASAP7_75t_L g2388 ( 
.A(n_2327),
.B(n_168),
.Y(n_2388)
);

OAI22xp33_ASAP7_75t_L g2389 ( 
.A1(n_2337),
.A2(n_172),
.B1(n_173),
.B2(n_171),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2347),
.B(n_170),
.Y(n_2390)
);

OAI22xp33_ASAP7_75t_L g2391 ( 
.A1(n_2338),
.A2(n_2312),
.B1(n_2333),
.B2(n_2329),
.Y(n_2391)
);

INVxp67_ASAP7_75t_L g2392 ( 
.A(n_2356),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_2355),
.B(n_175),
.Y(n_2393)
);

OR2x2_ASAP7_75t_L g2394 ( 
.A(n_2317),
.B(n_177),
.Y(n_2394)
);

AOI22xp5_ASAP7_75t_L g2395 ( 
.A1(n_2341),
.A2(n_2344),
.B1(n_2342),
.B2(n_2343),
.Y(n_2395)
);

NOR2xp33_ASAP7_75t_L g2396 ( 
.A(n_2332),
.B(n_177),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2358),
.B(n_178),
.Y(n_2397)
);

OAI22xp33_ASAP7_75t_L g2398 ( 
.A1(n_2330),
.A2(n_181),
.B1(n_182),
.B2(n_180),
.Y(n_2398)
);

AO221x2_ASAP7_75t_L g2399 ( 
.A1(n_2359),
.A2(n_2361),
.B1(n_2365),
.B2(n_2362),
.C(n_2360),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_2366),
.B(n_179),
.Y(n_2400)
);

INVx3_ASAP7_75t_L g2401 ( 
.A(n_2334),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2369),
.B(n_179),
.Y(n_2402)
);

AND2x4_ASAP7_75t_L g2403 ( 
.A(n_2325),
.B(n_182),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_2370),
.B(n_183),
.Y(n_2404)
);

NOR4xp25_ASAP7_75t_SL g2405 ( 
.A(n_2340),
.B(n_2310),
.C(n_2305),
.D(n_2296),
.Y(n_2405)
);

AND2x4_ASAP7_75t_L g2406 ( 
.A(n_2288),
.B(n_183),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_2298),
.B(n_186),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2307),
.B(n_187),
.Y(n_2408)
);

NAND2xp33_ASAP7_75t_SL g2409 ( 
.A(n_2345),
.B(n_187),
.Y(n_2409)
);

OAI22xp33_ASAP7_75t_L g2410 ( 
.A1(n_2318),
.A2(n_192),
.B1(n_193),
.B2(n_191),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_2316),
.B(n_190),
.Y(n_2411)
);

OAI22xp33_ASAP7_75t_L g2412 ( 
.A1(n_2322),
.A2(n_194),
.B1(n_195),
.B2(n_192),
.Y(n_2412)
);

AO221x2_ASAP7_75t_L g2413 ( 
.A1(n_2346),
.A2(n_196),
.B1(n_191),
.B2(n_195),
.C(n_197),
.Y(n_2413)
);

AND2x2_ASAP7_75t_L g2414 ( 
.A(n_2311),
.B(n_196),
.Y(n_2414)
);

CKINVDCx8_ASAP7_75t_R g2415 ( 
.A(n_2346),
.Y(n_2415)
);

AND2x4_ASAP7_75t_L g2416 ( 
.A(n_2331),
.B(n_198),
.Y(n_2416)
);

OAI22xp33_ASAP7_75t_L g2417 ( 
.A1(n_2286),
.A2(n_200),
.B1(n_201),
.B2(n_199),
.Y(n_2417)
);

CKINVDCx5p33_ASAP7_75t_R g2418 ( 
.A(n_2357),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_L g2419 ( 
.A(n_2303),
.B(n_2302),
.Y(n_2419)
);

AO221x2_ASAP7_75t_L g2420 ( 
.A1(n_2335),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.C(n_202),
.Y(n_2420)
);

OAI22xp33_ASAP7_75t_L g2421 ( 
.A1(n_2349),
.A2(n_204),
.B1(n_205),
.B2(n_203),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2301),
.B(n_2350),
.Y(n_2422)
);

NOR2xp33_ASAP7_75t_L g2423 ( 
.A(n_2304),
.B(n_202),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2315),
.B(n_2299),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2354),
.B(n_206),
.Y(n_2425)
);

NOR2xp33_ASAP7_75t_L g2426 ( 
.A(n_2336),
.B(n_207),
.Y(n_2426)
);

NOR2xp33_ASAP7_75t_R g2427 ( 
.A(n_2353),
.B(n_208),
.Y(n_2427)
);

INVx4_ASAP7_75t_L g2428 ( 
.A(n_2293),
.Y(n_2428)
);

INVxp67_ASAP7_75t_L g2429 ( 
.A(n_2328),
.Y(n_2429)
);

AO221x2_ASAP7_75t_L g2430 ( 
.A1(n_2372),
.A2(n_213),
.B1(n_209),
.B2(n_212),
.C(n_214),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2313),
.Y(n_2431)
);

NOR2xp33_ASAP7_75t_L g2432 ( 
.A(n_2371),
.B(n_214),
.Y(n_2432)
);

AO221x2_ASAP7_75t_L g2433 ( 
.A1(n_2294),
.A2(n_217),
.B1(n_215),
.B2(n_216),
.C(n_218),
.Y(n_2433)
);

NOR2x1_ASAP7_75t_L g2434 ( 
.A(n_2339),
.B(n_215),
.Y(n_2434)
);

HB1xp67_ASAP7_75t_L g2435 ( 
.A(n_2314),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2320),
.B(n_218),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2297),
.B(n_219),
.Y(n_2437)
);

AND2x2_ASAP7_75t_L g2438 ( 
.A(n_2309),
.B(n_220),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2323),
.B(n_221),
.Y(n_2439)
);

INVxp67_ASAP7_75t_L g2440 ( 
.A(n_2324),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2363),
.B(n_223),
.Y(n_2441)
);

AO221x2_ASAP7_75t_L g2442 ( 
.A1(n_2300),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.C(n_227),
.Y(n_2442)
);

NOR2xp33_ASAP7_75t_L g2443 ( 
.A(n_2321),
.B(n_224),
.Y(n_2443)
);

NOR2xp33_ASAP7_75t_R g2444 ( 
.A(n_2287),
.B(n_225),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2352),
.B(n_228),
.Y(n_2445)
);

NAND2xp33_ASAP7_75t_SL g2446 ( 
.A(n_2295),
.B(n_230),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2352),
.B(n_231),
.Y(n_2447)
);

BUFx12f_ASAP7_75t_L g2448 ( 
.A(n_2346),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2352),
.B(n_233),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2352),
.B(n_234),
.Y(n_2450)
);

CKINVDCx16_ASAP7_75t_R g2451 ( 
.A(n_2289),
.Y(n_2451)
);

NOR2xp33_ASAP7_75t_SL g2452 ( 
.A(n_2327),
.B(n_235),
.Y(n_2452)
);

CKINVDCx5p33_ASAP7_75t_R g2453 ( 
.A(n_2287),
.Y(n_2453)
);

BUFx3_ASAP7_75t_L g2454 ( 
.A(n_2287),
.Y(n_2454)
);

NOR4xp25_ASAP7_75t_SL g2455 ( 
.A(n_2352),
.B(n_240),
.C(n_237),
.D(n_239),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2352),
.B(n_237),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2352),
.B(n_241),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2352),
.B(n_241),
.Y(n_2458)
);

AND2x4_ASAP7_75t_L g2459 ( 
.A(n_2306),
.B(n_243),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2352),
.B(n_244),
.Y(n_2460)
);

NOR2xp67_ASAP7_75t_L g2461 ( 
.A(n_2327),
.B(n_245),
.Y(n_2461)
);

INVx2_ASAP7_75t_SL g2462 ( 
.A(n_2287),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_L g2463 ( 
.A(n_2352),
.B(n_247),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_2352),
.B(n_249),
.Y(n_2464)
);

NOR2xp33_ASAP7_75t_R g2465 ( 
.A(n_2287),
.B(n_250),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2352),
.B(n_251),
.Y(n_2466)
);

NOR2xp33_ASAP7_75t_L g2467 ( 
.A(n_2326),
.B(n_252),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_2352),
.B(n_254),
.Y(n_2468)
);

AO221x2_ASAP7_75t_L g2469 ( 
.A1(n_2319),
.A2(n_257),
.B1(n_255),
.B2(n_256),
.C(n_258),
.Y(n_2469)
);

INVx4_ASAP7_75t_L g2470 ( 
.A(n_2448),
.Y(n_2470)
);

OR2x2_ASAP7_75t_L g2471 ( 
.A(n_2419),
.B(n_256),
.Y(n_2471)
);

AND2x4_ASAP7_75t_L g2472 ( 
.A(n_2454),
.B(n_257),
.Y(n_2472)
);

BUFx3_ASAP7_75t_L g2473 ( 
.A(n_2415),
.Y(n_2473)
);

BUFx12f_ASAP7_75t_L g2474 ( 
.A(n_2375),
.Y(n_2474)
);

OR2x6_ASAP7_75t_L g2475 ( 
.A(n_2403),
.B(n_260),
.Y(n_2475)
);

AND2x2_ASAP7_75t_L g2476 ( 
.A(n_2414),
.B(n_261),
.Y(n_2476)
);

OAI22xp5_ASAP7_75t_L g2477 ( 
.A1(n_2386),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.Y(n_2477)
);

AND2x2_ASAP7_75t_L g2478 ( 
.A(n_2462),
.B(n_264),
.Y(n_2478)
);

AND2x2_ASAP7_75t_L g2479 ( 
.A(n_2378),
.B(n_265),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2431),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2435),
.Y(n_2481)
);

HB1xp67_ASAP7_75t_L g2482 ( 
.A(n_2424),
.Y(n_2482)
);

INVx1_ASAP7_75t_SL g2483 ( 
.A(n_2444),
.Y(n_2483)
);

INVxp67_ASAP7_75t_SL g2484 ( 
.A(n_2387),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_L g2485 ( 
.A(n_2391),
.B(n_266),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2440),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2437),
.Y(n_2487)
);

AND2x2_ASAP7_75t_L g2488 ( 
.A(n_2406),
.B(n_267),
.Y(n_2488)
);

OR2x6_ASAP7_75t_L g2489 ( 
.A(n_2461),
.B(n_267),
.Y(n_2489)
);

OR2x2_ASAP7_75t_L g2490 ( 
.A(n_2422),
.B(n_268),
.Y(n_2490)
);

BUFx3_ASAP7_75t_L g2491 ( 
.A(n_2453),
.Y(n_2491)
);

NOR2xp33_ASAP7_75t_SL g2492 ( 
.A(n_2451),
.B(n_270),
.Y(n_2492)
);

OR2x2_ASAP7_75t_L g2493 ( 
.A(n_2394),
.B(n_271),
.Y(n_2493)
);

AND2x2_ASAP7_75t_L g2494 ( 
.A(n_2405),
.B(n_272),
.Y(n_2494)
);

OR2x2_ASAP7_75t_L g2495 ( 
.A(n_2425),
.B(n_272),
.Y(n_2495)
);

INVx1_ASAP7_75t_SL g2496 ( 
.A(n_2465),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2439),
.Y(n_2497)
);

AO21x2_ASAP7_75t_L g2498 ( 
.A1(n_2374),
.A2(n_273),
.B(n_274),
.Y(n_2498)
);

NAND2xp33_ASAP7_75t_SL g2499 ( 
.A(n_2459),
.B(n_274),
.Y(n_2499)
);

AND2x2_ASAP7_75t_L g2500 ( 
.A(n_2429),
.B(n_276),
.Y(n_2500)
);

HB1xp67_ASAP7_75t_L g2501 ( 
.A(n_2390),
.Y(n_2501)
);

INVx4_ASAP7_75t_L g2502 ( 
.A(n_2418),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2401),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2436),
.Y(n_2504)
);

INVx1_ASAP7_75t_SL g2505 ( 
.A(n_2409),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2445),
.B(n_277),
.Y(n_2506)
);

AND2x2_ASAP7_75t_L g2507 ( 
.A(n_2393),
.B(n_278),
.Y(n_2507)
);

INVx1_ASAP7_75t_SL g2508 ( 
.A(n_2373),
.Y(n_2508)
);

BUFx3_ASAP7_75t_L g2509 ( 
.A(n_2416),
.Y(n_2509)
);

AND2x2_ASAP7_75t_L g2510 ( 
.A(n_2397),
.B(n_279),
.Y(n_2510)
);

OAI22xp5_ASAP7_75t_L g2511 ( 
.A1(n_2395),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_2511)
);

INVx2_ASAP7_75t_SL g2512 ( 
.A(n_2438),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_L g2513 ( 
.A(n_2447),
.B(n_282),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2379),
.Y(n_2514)
);

BUFx3_ASAP7_75t_L g2515 ( 
.A(n_2467),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2381),
.Y(n_2516)
);

AND2x2_ASAP7_75t_L g2517 ( 
.A(n_2400),
.B(n_2402),
.Y(n_2517)
);

INVx3_ASAP7_75t_SL g2518 ( 
.A(n_2376),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2383),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_2385),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2384),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2404),
.Y(n_2522)
);

OR2x2_ASAP7_75t_L g2523 ( 
.A(n_2449),
.B(n_283),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2450),
.B(n_284),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2456),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2457),
.B(n_286),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2458),
.Y(n_2527)
);

OAI21x1_ASAP7_75t_L g2528 ( 
.A1(n_2460),
.A2(n_286),
.B(n_287),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_2463),
.B(n_2464),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2466),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2468),
.Y(n_2531)
);

BUFx3_ASAP7_75t_L g2532 ( 
.A(n_2388),
.Y(n_2532)
);

AND2x2_ASAP7_75t_L g2533 ( 
.A(n_2426),
.B(n_287),
.Y(n_2533)
);

OR2x2_ASAP7_75t_L g2534 ( 
.A(n_2407),
.B(n_288),
.Y(n_2534)
);

NOR2xp33_ASAP7_75t_L g2535 ( 
.A(n_2452),
.B(n_288),
.Y(n_2535)
);

OR2x2_ASAP7_75t_L g2536 ( 
.A(n_2430),
.B(n_2469),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_2380),
.B(n_2443),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2420),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_2380),
.B(n_289),
.Y(n_2539)
);

AND2x2_ASAP7_75t_L g2540 ( 
.A(n_2432),
.B(n_290),
.Y(n_2540)
);

INVxp67_ASAP7_75t_L g2541 ( 
.A(n_2441),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2408),
.Y(n_2542)
);

NAND2x1_ASAP7_75t_SL g2543 ( 
.A(n_2423),
.B(n_291),
.Y(n_2543)
);

OR2x2_ASAP7_75t_L g2544 ( 
.A(n_2377),
.B(n_292),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2411),
.Y(n_2545)
);

INVx2_ASAP7_75t_SL g2546 ( 
.A(n_2413),
.Y(n_2546)
);

AND2x2_ASAP7_75t_L g2547 ( 
.A(n_2396),
.B(n_294),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2469),
.Y(n_2548)
);

INVxp67_ASAP7_75t_L g2549 ( 
.A(n_2446),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2410),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2412),
.Y(n_2551)
);

AND2x2_ASAP7_75t_L g2552 ( 
.A(n_2433),
.B(n_297),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2417),
.B(n_2421),
.Y(n_2553)
);

INVx3_ASAP7_75t_SL g2554 ( 
.A(n_2398),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2455),
.B(n_298),
.Y(n_2555)
);

OAI22xp5_ASAP7_75t_L g2556 ( 
.A1(n_2389),
.A2(n_300),
.B1(n_298),
.B2(n_299),
.Y(n_2556)
);

CKINVDCx16_ASAP7_75t_R g2557 ( 
.A(n_2386),
.Y(n_2557)
);

OR2x2_ASAP7_75t_L g2558 ( 
.A(n_2419),
.B(n_299),
.Y(n_2558)
);

AND2x4_ASAP7_75t_SL g2559 ( 
.A(n_2428),
.B(n_302),
.Y(n_2559)
);

AOI22xp33_ASAP7_75t_SL g2560 ( 
.A1(n_2442),
.A2(n_307),
.B1(n_303),
.B2(n_304),
.Y(n_2560)
);

AND2x2_ASAP7_75t_L g2561 ( 
.A(n_2399),
.B(n_308),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2382),
.Y(n_2562)
);

AND2x2_ASAP7_75t_L g2563 ( 
.A(n_2399),
.B(n_309),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2382),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2382),
.Y(n_2565)
);

NOR2xp33_ASAP7_75t_L g2566 ( 
.A(n_2392),
.B(n_310),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2382),
.Y(n_2567)
);

INVx1_ASAP7_75t_SL g2568 ( 
.A(n_2427),
.Y(n_2568)
);

OR2x6_ASAP7_75t_L g2569 ( 
.A(n_2448),
.B(n_311),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2382),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2382),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2382),
.Y(n_2572)
);

INVx1_ASAP7_75t_SL g2573 ( 
.A(n_2427),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2382),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_L g2575 ( 
.A(n_2391),
.B(n_313),
.Y(n_2575)
);

NAND2xp33_ASAP7_75t_SL g2576 ( 
.A(n_2444),
.B(n_314),
.Y(n_2576)
);

HB1xp67_ASAP7_75t_L g2577 ( 
.A(n_2382),
.Y(n_2577)
);

BUFx3_ASAP7_75t_L g2578 ( 
.A(n_2448),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2434),
.Y(n_2579)
);

AND2x2_ASAP7_75t_L g2580 ( 
.A(n_2399),
.B(n_315),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2382),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2382),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2382),
.Y(n_2583)
);

BUFx2_ASAP7_75t_L g2584 ( 
.A(n_2448),
.Y(n_2584)
);

HB1xp67_ASAP7_75t_L g2585 ( 
.A(n_2382),
.Y(n_2585)
);

NOR2xp33_ASAP7_75t_L g2586 ( 
.A(n_2392),
.B(n_317),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2391),
.B(n_319),
.Y(n_2587)
);

BUFx2_ASAP7_75t_L g2588 ( 
.A(n_2448),
.Y(n_2588)
);

AND3x1_ASAP7_75t_L g2589 ( 
.A(n_2387),
.B(n_320),
.C(n_321),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_L g2590 ( 
.A(n_2391),
.B(n_320),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2382),
.Y(n_2591)
);

INVxp67_ASAP7_75t_SL g2592 ( 
.A(n_2473),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2577),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2585),
.Y(n_2594)
);

NOR3xp33_ASAP7_75t_L g2595 ( 
.A(n_2557),
.B(n_322),
.C(n_323),
.Y(n_2595)
);

AOI322xp5_ASAP7_75t_L g2596 ( 
.A1(n_2548),
.A2(n_329),
.A3(n_328),
.B1(n_326),
.B2(n_324),
.C1(n_325),
.C2(n_327),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2501),
.B(n_2522),
.Y(n_2597)
);

INVx1_ASAP7_75t_SL g2598 ( 
.A(n_2474),
.Y(n_2598)
);

AOI21xp33_ASAP7_75t_SL g2599 ( 
.A1(n_2518),
.A2(n_338),
.B(n_328),
.Y(n_2599)
);

NOR2x1_ASAP7_75t_SL g2600 ( 
.A(n_2489),
.B(n_330),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_2584),
.Y(n_2601)
);

OAI221xp5_ASAP7_75t_L g2602 ( 
.A1(n_2536),
.A2(n_334),
.B1(n_332),
.B2(n_333),
.C(n_335),
.Y(n_2602)
);

AND2x4_ASAP7_75t_L g2603 ( 
.A(n_2520),
.B(n_333),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_SL g2604 ( 
.A(n_2561),
.B(n_335),
.Y(n_2604)
);

NOR2x1_ASAP7_75t_R g2605 ( 
.A(n_2470),
.B(n_338),
.Y(n_2605)
);

INVxp67_ASAP7_75t_L g2606 ( 
.A(n_2588),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2562),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2564),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2512),
.Y(n_2609)
);

OAI322xp33_ASAP7_75t_L g2610 ( 
.A1(n_2485),
.A2(n_346),
.A3(n_345),
.B1(n_343),
.B2(n_341),
.C1(n_342),
.C2(n_344),
.Y(n_2610)
);

AND2x2_ASAP7_75t_L g2611 ( 
.A(n_2482),
.B(n_343),
.Y(n_2611)
);

AOI222xp33_ASAP7_75t_L g2612 ( 
.A1(n_2539),
.A2(n_365),
.B1(n_352),
.B2(n_374),
.C1(n_359),
.C2(n_344),
.Y(n_2612)
);

AOI32xp33_ASAP7_75t_L g2613 ( 
.A1(n_2563),
.A2(n_348),
.A3(n_350),
.B1(n_347),
.B2(n_349),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2565),
.Y(n_2614)
);

INVxp33_ASAP7_75t_L g2615 ( 
.A(n_2492),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_2541),
.B(n_351),
.Y(n_2616)
);

INVxp67_ASAP7_75t_L g2617 ( 
.A(n_2484),
.Y(n_2617)
);

AND2x2_ASAP7_75t_L g2618 ( 
.A(n_2517),
.B(n_353),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_L g2619 ( 
.A(n_2575),
.B(n_354),
.Y(n_2619)
);

AOI21xp5_ASAP7_75t_L g2620 ( 
.A1(n_2537),
.A2(n_356),
.B(n_357),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_L g2621 ( 
.A(n_2587),
.B(n_358),
.Y(n_2621)
);

OR2x2_ASAP7_75t_L g2622 ( 
.A(n_2486),
.B(n_358),
.Y(n_2622)
);

NOR2xp33_ASAP7_75t_L g2623 ( 
.A(n_2502),
.B(n_2578),
.Y(n_2623)
);

AND2x2_ASAP7_75t_L g2624 ( 
.A(n_2580),
.B(n_360),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2567),
.Y(n_2625)
);

AOI21xp33_ASAP7_75t_L g2626 ( 
.A1(n_2494),
.A2(n_360),
.B(n_361),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2570),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_L g2628 ( 
.A(n_2590),
.B(n_361),
.Y(n_2628)
);

AOI32xp33_ASAP7_75t_L g2629 ( 
.A1(n_2552),
.A2(n_364),
.A3(n_366),
.B1(n_362),
.B2(n_365),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_L g2630 ( 
.A(n_2525),
.B(n_2527),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_L g2631 ( 
.A(n_2530),
.B(n_366),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2571),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_2531),
.B(n_367),
.Y(n_2633)
);

OAI22xp5_ASAP7_75t_L g2634 ( 
.A1(n_2546),
.A2(n_371),
.B1(n_367),
.B2(n_370),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2572),
.Y(n_2635)
);

OAI21xp5_ASAP7_75t_L g2636 ( 
.A1(n_2560),
.A2(n_370),
.B(n_371),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2574),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2581),
.Y(n_2638)
);

INVx1_ASAP7_75t_SL g2639 ( 
.A(n_2576),
.Y(n_2639)
);

AOI21xp5_ASAP7_75t_L g2640 ( 
.A1(n_2589),
.A2(n_372),
.B(n_373),
.Y(n_2640)
);

INVx1_ASAP7_75t_SL g2641 ( 
.A(n_2491),
.Y(n_2641)
);

BUFx3_ASAP7_75t_L g2642 ( 
.A(n_2569),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2582),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_2542),
.B(n_374),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2545),
.B(n_375),
.Y(n_2645)
);

NOR4xp25_ASAP7_75t_SL g2646 ( 
.A(n_2499),
.B(n_378),
.C(n_375),
.D(n_376),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2538),
.B(n_376),
.Y(n_2647)
);

AND2x2_ASAP7_75t_L g2648 ( 
.A(n_2521),
.B(n_380),
.Y(n_2648)
);

NOR2xp33_ASAP7_75t_L g2649 ( 
.A(n_2532),
.B(n_381),
.Y(n_2649)
);

NOR2xp33_ASAP7_75t_L g2650 ( 
.A(n_2505),
.B(n_382),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_L g2651 ( 
.A(n_2487),
.B(n_383),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2579),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2497),
.B(n_385),
.Y(n_2653)
);

AOI21xp5_ASAP7_75t_L g2654 ( 
.A1(n_2553),
.A2(n_385),
.B(n_386),
.Y(n_2654)
);

INVxp67_ASAP7_75t_L g2655 ( 
.A(n_2515),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2583),
.Y(n_2656)
);

A2O1A1Ixp33_ASAP7_75t_L g2657 ( 
.A1(n_2544),
.A2(n_388),
.B(n_386),
.C(n_387),
.Y(n_2657)
);

AND2x2_ASAP7_75t_L g2658 ( 
.A(n_2514),
.B(n_387),
.Y(n_2658)
);

AND2x2_ASAP7_75t_L g2659 ( 
.A(n_2516),
.B(n_389),
.Y(n_2659)
);

OAI22xp5_ASAP7_75t_L g2660 ( 
.A1(n_2554),
.A2(n_391),
.B1(n_389),
.B2(n_390),
.Y(n_2660)
);

INVx2_ASAP7_75t_SL g2661 ( 
.A(n_2509),
.Y(n_2661)
);

HB1xp67_ASAP7_75t_L g2662 ( 
.A(n_2591),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2480),
.Y(n_2663)
);

AOI21xp5_ASAP7_75t_L g2664 ( 
.A1(n_2508),
.A2(n_393),
.B(n_396),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2481),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2504),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2498),
.B(n_398),
.Y(n_2667)
);

INVxp67_ASAP7_75t_SL g2668 ( 
.A(n_2549),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_L g2669 ( 
.A(n_2519),
.B(n_403),
.Y(n_2669)
);

OR2x2_ASAP7_75t_L g2670 ( 
.A(n_2529),
.B(n_404),
.Y(n_2670)
);

AND2x2_ASAP7_75t_L g2671 ( 
.A(n_2478),
.B(n_406),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2550),
.Y(n_2672)
);

OAI22xp5_ASAP7_75t_L g2673 ( 
.A1(n_2471),
.A2(n_409),
.B1(n_407),
.B2(n_408),
.Y(n_2673)
);

OAI22xp5_ASAP7_75t_L g2674 ( 
.A1(n_2558),
.A2(n_410),
.B1(n_408),
.B2(n_409),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2551),
.Y(n_2675)
);

AND2x2_ASAP7_75t_L g2676 ( 
.A(n_2503),
.B(n_412),
.Y(n_2676)
);

OAI22xp33_ASAP7_75t_SL g2677 ( 
.A1(n_2490),
.A2(n_415),
.B1(n_413),
.B2(n_414),
.Y(n_2677)
);

AND2x2_ASAP7_75t_L g2678 ( 
.A(n_2592),
.B(n_2472),
.Y(n_2678)
);

NOR2xp33_ASAP7_75t_SL g2679 ( 
.A(n_2605),
.B(n_2568),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_L g2680 ( 
.A(n_2618),
.B(n_2540),
.Y(n_2680)
);

INVxp67_ASAP7_75t_SL g2681 ( 
.A(n_2600),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_SL g2682 ( 
.A(n_2617),
.B(n_2483),
.Y(n_2682)
);

NOR2xp33_ASAP7_75t_L g2683 ( 
.A(n_2598),
.B(n_2496),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2662),
.Y(n_2684)
);

NOR2xp33_ASAP7_75t_L g2685 ( 
.A(n_2641),
.B(n_2573),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_L g2686 ( 
.A(n_2611),
.B(n_2547),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2630),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2672),
.Y(n_2688)
);

OR2x2_ASAP7_75t_L g2689 ( 
.A(n_2597),
.B(n_2493),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_2654),
.B(n_2603),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2675),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2666),
.Y(n_2692)
);

OR2x2_ASAP7_75t_L g2693 ( 
.A(n_2668),
.B(n_2523),
.Y(n_2693)
);

NOR2xp33_ASAP7_75t_L g2694 ( 
.A(n_2606),
.B(n_2655),
.Y(n_2694)
);

AND2x2_ASAP7_75t_L g2695 ( 
.A(n_2601),
.B(n_2559),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2603),
.B(n_2507),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2648),
.B(n_2510),
.Y(n_2697)
);

CKINVDCx20_ASAP7_75t_R g2698 ( 
.A(n_2642),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_L g2699 ( 
.A(n_2658),
.B(n_2533),
.Y(n_2699)
);

AOI21xp5_ASAP7_75t_SL g2700 ( 
.A1(n_2657),
.A2(n_2535),
.B(n_2477),
.Y(n_2700)
);

CKINVDCx5p33_ASAP7_75t_R g2701 ( 
.A(n_2623),
.Y(n_2701)
);

NOR2xp33_ASAP7_75t_L g2702 ( 
.A(n_2670),
.B(n_2639),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_SL g2703 ( 
.A(n_2661),
.B(n_2566),
.Y(n_2703)
);

INVxp67_ASAP7_75t_L g2704 ( 
.A(n_2649),
.Y(n_2704)
);

AND2x2_ASAP7_75t_L g2705 ( 
.A(n_2609),
.B(n_2476),
.Y(n_2705)
);

HB1xp67_ASAP7_75t_L g2706 ( 
.A(n_2622),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_2659),
.B(n_2479),
.Y(n_2707)
);

AND2x2_ASAP7_75t_L g2708 ( 
.A(n_2624),
.B(n_2500),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2607),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2608),
.Y(n_2710)
);

AND2x4_ASAP7_75t_L g2711 ( 
.A(n_2593),
.B(n_2475),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_L g2712 ( 
.A(n_2620),
.B(n_2613),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2614),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2612),
.B(n_2586),
.Y(n_2714)
);

AOI221xp5_ASAP7_75t_L g2715 ( 
.A1(n_2626),
.A2(n_2511),
.B1(n_2555),
.B2(n_2556),
.C(n_2513),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_L g2716 ( 
.A(n_2677),
.B(n_2534),
.Y(n_2716)
);

AOI222xp33_ASAP7_75t_L g2717 ( 
.A1(n_2636),
.A2(n_2526),
.B1(n_2524),
.B2(n_2506),
.C1(n_2528),
.C2(n_2488),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2625),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_SL g2719 ( 
.A(n_2599),
.B(n_2495),
.Y(n_2719)
);

AND2x4_ASAP7_75t_L g2720 ( 
.A(n_2594),
.B(n_2475),
.Y(n_2720)
);

NOR2xp33_ASAP7_75t_L g2721 ( 
.A(n_2604),
.B(n_2543),
.Y(n_2721)
);

OR2x2_ASAP7_75t_L g2722 ( 
.A(n_2665),
.B(n_414),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2627),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2632),
.Y(n_2724)
);

NOR2xp33_ASAP7_75t_L g2725 ( 
.A(n_2615),
.B(n_416),
.Y(n_2725)
);

INVx3_ASAP7_75t_L g2726 ( 
.A(n_2676),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2635),
.Y(n_2727)
);

AND2x2_ASAP7_75t_L g2728 ( 
.A(n_2671),
.B(n_417),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2637),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2638),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2643),
.Y(n_2731)
);

AND2x2_ASAP7_75t_L g2732 ( 
.A(n_2650),
.B(n_418),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2656),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2629),
.B(n_418),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_2667),
.B(n_419),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2664),
.B(n_419),
.Y(n_2736)
);

NOR2xp33_ASAP7_75t_L g2737 ( 
.A(n_2619),
.B(n_421),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2663),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_2698),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2706),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2688),
.Y(n_2741)
);

INVx5_ASAP7_75t_SL g2742 ( 
.A(n_2711),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2691),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2735),
.Y(n_2744)
);

HB1xp67_ASAP7_75t_L g2745 ( 
.A(n_2708),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2678),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2722),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_2726),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2726),
.B(n_2595),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2709),
.Y(n_2750)
);

AND2x2_ASAP7_75t_L g2751 ( 
.A(n_2681),
.B(n_2621),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2710),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2713),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2705),
.B(n_2660),
.Y(n_2754)
);

BUFx2_ASAP7_75t_L g2755 ( 
.A(n_2701),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2718),
.Y(n_2756)
);

HB1xp67_ASAP7_75t_SL g2757 ( 
.A(n_2685),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2723),
.Y(n_2758)
);

INVx2_ASAP7_75t_L g2759 ( 
.A(n_2693),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2724),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2727),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2729),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2730),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2731),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2696),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2733),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2680),
.B(n_2644),
.Y(n_2767)
);

CKINVDCx5p33_ASAP7_75t_R g2768 ( 
.A(n_2683),
.Y(n_2768)
);

BUFx4_ASAP7_75t_SL g2769 ( 
.A(n_2684),
.Y(n_2769)
);

INVx3_ASAP7_75t_L g2770 ( 
.A(n_2711),
.Y(n_2770)
);

HB1xp67_ASAP7_75t_L g2771 ( 
.A(n_2686),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2738),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2692),
.Y(n_2773)
);

HB1xp67_ASAP7_75t_L g2774 ( 
.A(n_2707),
.Y(n_2774)
);

INVxp67_ASAP7_75t_L g2775 ( 
.A(n_2679),
.Y(n_2775)
);

HB1xp67_ASAP7_75t_L g2776 ( 
.A(n_2697),
.Y(n_2776)
);

HB1xp67_ASAP7_75t_L g2777 ( 
.A(n_2699),
.Y(n_2777)
);

CKINVDCx5p33_ASAP7_75t_R g2778 ( 
.A(n_2728),
.Y(n_2778)
);

AND2x2_ASAP7_75t_L g2779 ( 
.A(n_2695),
.B(n_2628),
.Y(n_2779)
);

INVx2_ASAP7_75t_L g2780 ( 
.A(n_2720),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_2720),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2689),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2687),
.Y(n_2783)
);

HB1xp67_ASAP7_75t_L g2784 ( 
.A(n_2694),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2725),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2736),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2734),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2682),
.Y(n_2788)
);

NOR2xp33_ASAP7_75t_L g2789 ( 
.A(n_2690),
.B(n_2645),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2732),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2716),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2737),
.Y(n_2792)
);

INVx2_ASAP7_75t_SL g2793 ( 
.A(n_2703),
.Y(n_2793)
);

INVxp67_ASAP7_75t_L g2794 ( 
.A(n_2721),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2704),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2719),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2702),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2712),
.Y(n_2798)
);

INVx3_ASAP7_75t_L g2799 ( 
.A(n_2714),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2717),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2715),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2700),
.Y(n_2802)
);

OA211x2_ASAP7_75t_L g2803 ( 
.A1(n_2775),
.A2(n_2789),
.B(n_2794),
.C(n_2749),
.Y(n_2803)
);

AND4x2_ASAP7_75t_L g2804 ( 
.A(n_2757),
.B(n_2640),
.C(n_2602),
.D(n_2596),
.Y(n_2804)
);

NAND3xp33_ASAP7_75t_SL g2805 ( 
.A(n_2802),
.B(n_2768),
.C(n_2778),
.Y(n_2805)
);

NAND4xp75_ASAP7_75t_L g2806 ( 
.A(n_2791),
.B(n_2647),
.C(n_2631),
.D(n_2633),
.Y(n_2806)
);

NOR2x1_ASAP7_75t_L g2807 ( 
.A(n_2755),
.B(n_2616),
.Y(n_2807)
);

NOR2xp33_ASAP7_75t_L g2808 ( 
.A(n_2739),
.B(n_2653),
.Y(n_2808)
);

AOI211x1_ASAP7_75t_SL g2809 ( 
.A1(n_2746),
.A2(n_2634),
.B(n_2652),
.C(n_2673),
.Y(n_2809)
);

NOR2xp33_ASAP7_75t_L g2810 ( 
.A(n_2784),
.B(n_2651),
.Y(n_2810)
);

AND2x2_ASAP7_75t_L g2811 ( 
.A(n_2742),
.B(n_2669),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_2790),
.B(n_2674),
.Y(n_2812)
);

NOR3x1_ASAP7_75t_L g2813 ( 
.A(n_2793),
.B(n_2610),
.C(n_2646),
.Y(n_2813)
);

NAND5xp2_ASAP7_75t_L g2814 ( 
.A(n_2798),
.B(n_2782),
.C(n_2788),
.D(n_2796),
.E(n_2797),
.Y(n_2814)
);

NOR3xp33_ASAP7_75t_L g2815 ( 
.A(n_2799),
.B(n_424),
.C(n_426),
.Y(n_2815)
);

NOR2xp33_ASAP7_75t_L g2816 ( 
.A(n_2770),
.B(n_424),
.Y(n_2816)
);

NOR3xp33_ASAP7_75t_L g2817 ( 
.A(n_2799),
.B(n_426),
.C(n_427),
.Y(n_2817)
);

NAND2x1_ASAP7_75t_L g2818 ( 
.A(n_2748),
.B(n_428),
.Y(n_2818)
);

NAND3xp33_ASAP7_75t_L g2819 ( 
.A(n_2801),
.B(n_431),
.C(n_432),
.Y(n_2819)
);

AOI22xp33_ASAP7_75t_L g2820 ( 
.A1(n_2800),
.A2(n_436),
.B1(n_433),
.B2(n_435),
.Y(n_2820)
);

NOR3xp33_ASAP7_75t_L g2821 ( 
.A(n_2795),
.B(n_437),
.C(n_438),
.Y(n_2821)
);

NOR2xp33_ASAP7_75t_L g2822 ( 
.A(n_2792),
.B(n_438),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_L g2823 ( 
.A(n_2776),
.B(n_439),
.Y(n_2823)
);

NOR3x1_ASAP7_75t_L g2824 ( 
.A(n_2767),
.B(n_440),
.C(n_441),
.Y(n_2824)
);

NAND4xp25_ASAP7_75t_L g2825 ( 
.A(n_2751),
.B(n_442),
.C(n_440),
.D(n_441),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2745),
.Y(n_2826)
);

NAND3xp33_ASAP7_75t_L g2827 ( 
.A(n_2786),
.B(n_443),
.C(n_444),
.Y(n_2827)
);

NOR3xp33_ASAP7_75t_L g2828 ( 
.A(n_2787),
.B(n_445),
.C(n_446),
.Y(n_2828)
);

NAND3xp33_ASAP7_75t_L g2829 ( 
.A(n_2780),
.B(n_2781),
.C(n_2759),
.Y(n_2829)
);

NOR4xp75_ASAP7_75t_L g2830 ( 
.A(n_2754),
.B(n_447),
.C(n_445),
.D(n_446),
.Y(n_2830)
);

OAI21xp33_ASAP7_75t_L g2831 ( 
.A1(n_2779),
.A2(n_448),
.B(n_449),
.Y(n_2831)
);

NOR3xp33_ASAP7_75t_SL g2832 ( 
.A(n_2740),
.B(n_450),
.C(n_451),
.Y(n_2832)
);

NOR2x1_ASAP7_75t_L g2833 ( 
.A(n_2765),
.B(n_452),
.Y(n_2833)
);

AND2x2_ASAP7_75t_L g2834 ( 
.A(n_2742),
.B(n_453),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_2774),
.B(n_454),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_L g2836 ( 
.A(n_2777),
.B(n_455),
.Y(n_2836)
);

OAI21xp5_ASAP7_75t_SL g2837 ( 
.A1(n_2771),
.A2(n_456),
.B(n_457),
.Y(n_2837)
);

INVx2_ASAP7_75t_L g2838 ( 
.A(n_2769),
.Y(n_2838)
);

INVxp67_ASAP7_75t_L g2839 ( 
.A(n_2747),
.Y(n_2839)
);

NOR3xp33_ASAP7_75t_L g2840 ( 
.A(n_2744),
.B(n_458),
.C(n_460),
.Y(n_2840)
);

AOI21xp5_ASAP7_75t_L g2841 ( 
.A1(n_2785),
.A2(n_461),
.B(n_462),
.Y(n_2841)
);

AOI221xp5_ASAP7_75t_L g2842 ( 
.A1(n_2783),
.A2(n_464),
.B1(n_461),
.B2(n_463),
.C(n_465),
.Y(n_2842)
);

AOI21xp5_ASAP7_75t_L g2843 ( 
.A1(n_2741),
.A2(n_464),
.B(n_466),
.Y(n_2843)
);

NOR4xp25_ASAP7_75t_L g2844 ( 
.A(n_2743),
.B(n_468),
.C(n_466),
.D(n_467),
.Y(n_2844)
);

OAI221xp5_ASAP7_75t_L g2845 ( 
.A1(n_2844),
.A2(n_2753),
.B1(n_2756),
.B2(n_2752),
.C(n_2750),
.Y(n_2845)
);

NOR2x1_ASAP7_75t_L g2846 ( 
.A(n_2814),
.B(n_2758),
.Y(n_2846)
);

CKINVDCx5p33_ASAP7_75t_R g2847 ( 
.A(n_2838),
.Y(n_2847)
);

AND2x4_ASAP7_75t_SL g2848 ( 
.A(n_2811),
.B(n_2760),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2829),
.Y(n_2849)
);

NOR3xp33_ASAP7_75t_L g2850 ( 
.A(n_2805),
.B(n_2762),
.C(n_2761),
.Y(n_2850)
);

OAI22xp5_ASAP7_75t_L g2851 ( 
.A1(n_2807),
.A2(n_2764),
.B1(n_2766),
.B2(n_2763),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2823),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_2809),
.B(n_2772),
.Y(n_2853)
);

AOI22xp5_ASAP7_75t_SL g2854 ( 
.A1(n_2834),
.A2(n_2773),
.B1(n_472),
.B2(n_469),
.Y(n_2854)
);

AND4x1_ASAP7_75t_L g2855 ( 
.A(n_2813),
.B(n_474),
.C(n_471),
.D(n_473),
.Y(n_2855)
);

OAI22xp5_ASAP7_75t_L g2856 ( 
.A1(n_2803),
.A2(n_477),
.B1(n_475),
.B2(n_476),
.Y(n_2856)
);

OAI322xp33_ASAP7_75t_L g2857 ( 
.A1(n_2839),
.A2(n_482),
.A3(n_481),
.B1(n_479),
.B2(n_475),
.C1(n_478),
.C2(n_480),
.Y(n_2857)
);

A2O1A1Ixp33_ASAP7_75t_SL g2858 ( 
.A1(n_2826),
.A2(n_483),
.B(n_479),
.C(n_481),
.Y(n_2858)
);

NOR3xp33_ASAP7_75t_L g2859 ( 
.A(n_2819),
.B(n_483),
.C(n_485),
.Y(n_2859)
);

OAI21xp33_ASAP7_75t_L g2860 ( 
.A1(n_2810),
.A2(n_2808),
.B(n_2812),
.Y(n_2860)
);

INVx1_ASAP7_75t_SL g2861 ( 
.A(n_2830),
.Y(n_2861)
);

OAI21xp5_ASAP7_75t_L g2862 ( 
.A1(n_2837),
.A2(n_491),
.B(n_492),
.Y(n_2862)
);

NAND4xp75_ASAP7_75t_L g2863 ( 
.A(n_2824),
.B(n_494),
.C(n_492),
.D(n_493),
.Y(n_2863)
);

AOI221xp5_ASAP7_75t_L g2864 ( 
.A1(n_2841),
.A2(n_2843),
.B1(n_2822),
.B2(n_2817),
.C(n_2815),
.Y(n_2864)
);

AOI22xp33_ASAP7_75t_L g2865 ( 
.A1(n_2833),
.A2(n_498),
.B1(n_496),
.B2(n_497),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2832),
.B(n_497),
.Y(n_2866)
);

OAI221xp5_ASAP7_75t_R g2867 ( 
.A1(n_2804),
.A2(n_501),
.B1(n_498),
.B2(n_499),
.C(n_502),
.Y(n_2867)
);

OAI221xp5_ASAP7_75t_L g2868 ( 
.A1(n_2818),
.A2(n_507),
.B1(n_504),
.B2(n_505),
.C(n_508),
.Y(n_2868)
);

AOI22xp33_ASAP7_75t_L g2869 ( 
.A1(n_2821),
.A2(n_508),
.B1(n_504),
.B2(n_505),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2835),
.Y(n_2870)
);

AOI22xp33_ASAP7_75t_L g2871 ( 
.A1(n_2820),
.A2(n_511),
.B1(n_509),
.B2(n_510),
.Y(n_2871)
);

AOI221xp5_ASAP7_75t_L g2872 ( 
.A1(n_2828),
.A2(n_513),
.B1(n_509),
.B2(n_512),
.C(n_514),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2836),
.Y(n_2873)
);

OAI21xp5_ASAP7_75t_L g2874 ( 
.A1(n_2806),
.A2(n_517),
.B(n_519),
.Y(n_2874)
);

NAND3xp33_ASAP7_75t_L g2875 ( 
.A(n_2840),
.B(n_520),
.C(n_521),
.Y(n_2875)
);

AOI221xp5_ASAP7_75t_L g2876 ( 
.A1(n_2827),
.A2(n_524),
.B1(n_521),
.B2(n_523),
.C(n_525),
.Y(n_2876)
);

OAI221xp5_ASAP7_75t_L g2877 ( 
.A1(n_2825),
.A2(n_526),
.B1(n_523),
.B2(n_524),
.C(n_527),
.Y(n_2877)
);

AND2x2_ASAP7_75t_L g2878 ( 
.A(n_2816),
.B(n_528),
.Y(n_2878)
);

A2O1A1Ixp33_ASAP7_75t_L g2879 ( 
.A1(n_2831),
.A2(n_531),
.B(n_529),
.C(n_530),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2842),
.Y(n_2880)
);

NOR3xp33_ASAP7_75t_SL g2881 ( 
.A(n_2814),
.B(n_534),
.C(n_535),
.Y(n_2881)
);

XOR2x2_ASAP7_75t_L g2882 ( 
.A(n_2863),
.B(n_535),
.Y(n_2882)
);

NOR2x1_ASAP7_75t_L g2883 ( 
.A(n_2846),
.B(n_536),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_2854),
.B(n_536),
.Y(n_2884)
);

AND2x2_ASAP7_75t_L g2885 ( 
.A(n_2847),
.B(n_537),
.Y(n_2885)
);

INVx2_ASAP7_75t_L g2886 ( 
.A(n_2878),
.Y(n_2886)
);

OR2x2_ASAP7_75t_L g2887 ( 
.A(n_2849),
.B(n_537),
.Y(n_2887)
);

AND2x2_ASAP7_75t_L g2888 ( 
.A(n_2848),
.B(n_538),
.Y(n_2888)
);

INVx3_ASAP7_75t_L g2889 ( 
.A(n_2855),
.Y(n_2889)
);

OR2x2_ASAP7_75t_L g2890 ( 
.A(n_2853),
.B(n_540),
.Y(n_2890)
);

NOR2xp33_ASAP7_75t_L g2891 ( 
.A(n_2861),
.B(n_541),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2866),
.Y(n_2892)
);

NOR2x1_ASAP7_75t_L g2893 ( 
.A(n_2856),
.B(n_542),
.Y(n_2893)
);

AND2x2_ASAP7_75t_L g2894 ( 
.A(n_2881),
.B(n_543),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2857),
.Y(n_2895)
);

NAND2x1p5_ASAP7_75t_L g2896 ( 
.A(n_2852),
.B(n_545),
.Y(n_2896)
);

INVx2_ASAP7_75t_SL g2897 ( 
.A(n_2851),
.Y(n_2897)
);

OR2x2_ASAP7_75t_L g2898 ( 
.A(n_2845),
.B(n_546),
.Y(n_2898)
);

XNOR2xp5_ASAP7_75t_L g2899 ( 
.A(n_2877),
.B(n_546),
.Y(n_2899)
);

AO22x2_ASAP7_75t_L g2900 ( 
.A1(n_2880),
.A2(n_2850),
.B1(n_2874),
.B2(n_2873),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2870),
.Y(n_2901)
);

NAND2xp5_ASAP7_75t_L g2902 ( 
.A(n_2858),
.B(n_2860),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_SL g2903 ( 
.A(n_2883),
.B(n_2864),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_SL g2904 ( 
.A(n_2889),
.B(n_2862),
.Y(n_2904)
);

NAND2xp33_ASAP7_75t_SL g2905 ( 
.A(n_2897),
.B(n_2888),
.Y(n_2905)
);

NOR2xp33_ASAP7_75t_R g2906 ( 
.A(n_2885),
.B(n_2865),
.Y(n_2906)
);

NAND2xp33_ASAP7_75t_SL g2907 ( 
.A(n_2890),
.B(n_2867),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_L g2908 ( 
.A(n_2886),
.B(n_2894),
.Y(n_2908)
);

NOR2xp33_ASAP7_75t_R g2909 ( 
.A(n_2902),
.B(n_2869),
.Y(n_2909)
);

NAND2xp33_ASAP7_75t_SL g2910 ( 
.A(n_2898),
.B(n_2871),
.Y(n_2910)
);

XNOR2x1_ASAP7_75t_L g2911 ( 
.A(n_2900),
.B(n_2875),
.Y(n_2911)
);

NOR2xp33_ASAP7_75t_R g2912 ( 
.A(n_2901),
.B(n_548),
.Y(n_2912)
);

NOR2xp33_ASAP7_75t_R g2913 ( 
.A(n_2899),
.B(n_549),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2896),
.B(n_2879),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2911),
.Y(n_2915)
);

AOI22xp5_ASAP7_75t_L g2916 ( 
.A1(n_2907),
.A2(n_2892),
.B1(n_2893),
.B2(n_2891),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2914),
.Y(n_2917)
);

INVx2_ASAP7_75t_L g2918 ( 
.A(n_2904),
.Y(n_2918)
);

AOI221x1_ASAP7_75t_L g2919 ( 
.A1(n_2905),
.A2(n_2900),
.B1(n_2895),
.B2(n_2884),
.C(n_2859),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2918),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2915),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2920),
.Y(n_2922)
);

INVx1_ASAP7_75t_SL g2923 ( 
.A(n_2921),
.Y(n_2923)
);

AOI22xp33_ASAP7_75t_L g2924 ( 
.A1(n_2923),
.A2(n_2910),
.B1(n_2917),
.B2(n_2903),
.Y(n_2924)
);

AOI31xp33_ASAP7_75t_L g2925 ( 
.A1(n_2922),
.A2(n_2916),
.A3(n_2908),
.B(n_2887),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_SL g2926 ( 
.A(n_2924),
.B(n_2912),
.Y(n_2926)
);

XNOR2xp5_ASAP7_75t_L g2927 ( 
.A(n_2925),
.B(n_2882),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2927),
.Y(n_2928)
);

XNOR2xp5_ASAP7_75t_L g2929 ( 
.A(n_2926),
.B(n_2919),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2929),
.Y(n_2930)
);

OAI221xp5_ASAP7_75t_R g2931 ( 
.A1(n_2930),
.A2(n_2928),
.B1(n_2909),
.B2(n_2913),
.C(n_2906),
.Y(n_2931)
);

AOI211xp5_ASAP7_75t_L g2932 ( 
.A1(n_2931),
.A2(n_2868),
.B(n_2876),
.C(n_2872),
.Y(n_2932)
);


endmodule