module fake_jpeg_10607_n_278 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_278);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_278;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_41),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

CKINVDCx6p67_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_19),
.Y(n_60)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_8),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_44),
.B(n_24),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_34),
.B1(n_19),
.B2(n_42),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_45),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_48),
.Y(n_85)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_51),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_39),
.B(n_17),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_54),
.Y(n_71)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_66),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_20),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_34),
.B1(n_23),
.B2(n_20),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_68),
.A2(n_17),
.B1(n_24),
.B2(n_29),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_69),
.B(n_73),
.Y(n_105)
);

AO22x1_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_72),
.A2(n_86),
.B(n_30),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_51),
.A2(n_26),
.B1(n_32),
.B2(n_25),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_79),
.A2(n_52),
.B1(n_58),
.B2(n_67),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_0),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_83),
.A2(n_87),
.B(n_62),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_0),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_23),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_89),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_33),
.Y(n_89)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_92),
.Y(n_101)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_94),
.A2(n_109),
.B1(n_113),
.B2(n_115),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

OA21x2_ASAP7_75t_L g118 ( 
.A1(n_96),
.A2(n_72),
.B(n_73),
.Y(n_118)
);

AOI32xp33_ASAP7_75t_L g97 ( 
.A1(n_89),
.A2(n_57),
.A3(n_67),
.B1(n_63),
.B2(n_52),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_100),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_98),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_31),
.B(n_68),
.C(n_27),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_99),
.B(n_103),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_59),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_104),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_47),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_107),
.Y(n_131)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_108),
.B(n_93),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_46),
.B1(n_53),
.B2(n_49),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_110),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_59),
.C(n_64),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_116),
.Y(n_120)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_79),
.A2(n_48),
.B1(n_65),
.B2(n_25),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_47),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_114),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_79),
.A2(n_28),
.B1(n_46),
.B2(n_27),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_59),
.C(n_47),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_46),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_83),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_118),
.A2(n_140),
.B1(n_30),
.B2(n_2),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_124),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_87),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_87),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_129),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_127),
.B(n_135),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_84),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_141),
.Y(n_165)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_99),
.A2(n_69),
.B(n_76),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_139),
.Y(n_163)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g140 ( 
.A1(n_94),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_98),
.B(n_71),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_105),
.B(n_78),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_28),
.Y(n_167)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_30),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_130),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_145),
.C(n_146),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_116),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_96),
.C(n_115),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_137),
.B(n_141),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_147),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_143),
.A2(n_112),
.B1(n_110),
.B2(n_107),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_148),
.A2(n_170),
.B1(n_125),
.B2(n_132),
.Y(n_181)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_149),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_123),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_152),
.Y(n_171)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

O2A1O1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_95),
.B(n_74),
.C(n_102),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_154),
.A2(n_155),
.B(n_157),
.Y(n_175)
);

AND2x6_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_1),
.Y(n_155)
);

NOR2x1_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_75),
.Y(n_156)
);

AO21x1_ASAP7_75t_L g180 ( 
.A1(n_156),
.A2(n_166),
.B(n_167),
.Y(n_180)
);

AND2x6_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_128),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_119),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_159),
.A2(n_162),
.B(n_169),
.Y(n_192)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_164),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_128),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_138),
.A2(n_30),
.B1(n_2),
.B2(n_4),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_168),
.A2(n_123),
.B1(n_125),
.B2(n_137),
.Y(n_183)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_163),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_178),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_120),
.C(n_126),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_179),
.C(n_189),
.Y(n_195)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_165),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_122),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_181),
.A2(n_183),
.B1(n_169),
.B2(n_159),
.Y(n_204)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_184),
.Y(n_197)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

NAND2xp33_ASAP7_75t_SL g185 ( 
.A(n_156),
.B(n_140),
.Y(n_185)
);

AOI21xp33_ASAP7_75t_L g209 ( 
.A1(n_185),
.A2(n_190),
.B(n_164),
.Y(n_209)
);

AO21x1_ASAP7_75t_L g186 ( 
.A1(n_151),
.A2(n_118),
.B(n_124),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_188),
.Y(n_205)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_167),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_151),
.B(n_134),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_L g190 ( 
.A1(n_158),
.A2(n_140),
.B(n_118),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_170),
.A2(n_118),
.B1(n_140),
.B2(n_135),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_191),
.A2(n_154),
.B1(n_162),
.B2(n_158),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_150),
.Y(n_193)
);

INVxp33_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_121),
.C(n_139),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_146),
.C(n_160),
.Y(n_206)
);

NOR2xp67_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_155),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_198),
.B(n_199),
.Y(n_218)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_192),
.B(n_157),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_200),
.B(n_175),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_201),
.A2(n_183),
.B1(n_187),
.B2(n_180),
.Y(n_229)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_207),
.C(n_208),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_168),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_161),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_209),
.A2(n_187),
.B(n_174),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_152),
.C(n_121),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_182),
.C(n_178),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_192),
.Y(n_212)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_212),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_189),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_175),
.A2(n_149),
.B1(n_4),
.B2(n_5),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_214),
.A2(n_177),
.B1(n_7),
.B2(n_9),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_1),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_6),
.Y(n_232)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_230),
.C(n_206),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_222),
.A2(n_203),
.B(n_207),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_213),
.A2(n_172),
.B1(n_184),
.B2(n_191),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_225),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_188),
.Y(n_226)
);

O2A1O1Ixp33_ASAP7_75t_L g239 ( 
.A1(n_226),
.A2(n_229),
.B(n_200),
.C(n_203),
.Y(n_239)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_215),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_232),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_177),
.C(n_180),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_231),
.A2(n_205),
.B1(n_201),
.B2(n_214),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_237),
.C(n_240),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_195),
.C(n_211),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_233),
.C(n_220),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_208),
.Y(n_237)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_238),
.Y(n_245)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_239),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_230),
.C(n_221),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_224),
.C(n_226),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_223),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_244),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_250),
.C(n_254),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_225),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_251),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_218),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_239),
.A2(n_217),
.B1(n_229),
.B2(n_216),
.Y(n_253)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_253),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_222),
.C(n_232),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_236),
.Y(n_255)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_255),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_245),
.A2(n_252),
.B1(n_234),
.B2(n_248),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_256),
.B(n_258),
.Y(n_267)
);

OAI21x1_ASAP7_75t_L g257 ( 
.A1(n_247),
.A2(n_234),
.B(n_210),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_257),
.B(n_6),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_231),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_6),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_7),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_263),
.A2(n_264),
.B1(n_10),
.B2(n_11),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_260),
.A2(n_16),
.B1(n_10),
.B2(n_11),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_265),
.B(n_13),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_255),
.Y(n_268)
);

A2O1A1Ixp33_ASAP7_75t_SL g272 ( 
.A1(n_268),
.A2(n_262),
.B(n_14),
.C(n_15),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_270),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_267),
.A2(n_259),
.B(n_261),
.Y(n_271)
);

INVxp33_ASAP7_75t_L g273 ( 
.A(n_271),
.Y(n_273)
);

INVxp33_ASAP7_75t_L g275 ( 
.A(n_273),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_275),
.A2(n_266),
.B(n_274),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_272),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_13),
.Y(n_278)
);


endmodule