module fake_aes_7068_n_857 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_857);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_857;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_227;
wire n_384;
wire n_163;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_455;
wire n_529;
wire n_312;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_490;
wire n_247;
wire n_393;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_482;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_466;
wire n_302;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g111 ( .A(n_58), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_53), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_41), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_103), .Y(n_114) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_39), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_6), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_14), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_15), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_9), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_104), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_96), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_65), .Y(n_122) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_79), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_19), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_107), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_33), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_106), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_56), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_12), .Y(n_129) );
INVx1_ASAP7_75t_SL g130 ( .A(n_98), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_51), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_7), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_91), .Y(n_133) );
BUFx2_ASAP7_75t_L g134 ( .A(n_5), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_7), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_59), .Y(n_136) );
CKINVDCx16_ASAP7_75t_R g137 ( .A(n_38), .Y(n_137) );
BUFx10_ASAP7_75t_L g138 ( .A(n_74), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_44), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_55), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_31), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_88), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_87), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_14), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g145 ( .A(n_47), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_67), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_105), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_42), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_75), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_27), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_84), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_25), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_100), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_95), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_85), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_117), .B(n_0), .Y(n_156) );
INVx2_ASAP7_75t_SL g157 ( .A(n_138), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_134), .B(n_0), .Y(n_158) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_134), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_117), .B(n_1), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_115), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_123), .B(n_118), .Y(n_162) );
INVx5_ASAP7_75t_L g163 ( .A(n_115), .Y(n_163) );
BUFx3_ASAP7_75t_L g164 ( .A(n_114), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_111), .B(n_1), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_111), .B(n_2), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_115), .Y(n_167) );
INVx4_ASAP7_75t_L g168 ( .A(n_150), .Y(n_168) );
BUFx12f_ASAP7_75t_L g169 ( .A(n_138), .Y(n_169) );
BUFx8_ASAP7_75t_SL g170 ( .A(n_116), .Y(n_170) );
INVx2_ASAP7_75t_SL g171 ( .A(n_138), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_115), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_115), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_114), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_150), .Y(n_175) );
BUFx3_ASAP7_75t_L g176 ( .A(n_138), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_113), .B(n_2), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_113), .B(n_3), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_118), .B(n_3), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_156), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_156), .Y(n_181) );
AOI22xp5_ASAP7_75t_L g182 ( .A1(n_159), .A2(n_137), .B1(n_119), .B2(n_141), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_168), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_159), .A2(n_126), .B1(n_132), .B2(n_135), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_156), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_158), .A2(n_124), .B1(n_152), .B2(n_129), .Y(n_186) );
OAI22xp33_ASAP7_75t_SL g187 ( .A1(n_162), .A2(n_129), .B1(n_152), .B2(n_155), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_168), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_156), .Y(n_189) );
OAI22xp33_ASAP7_75t_SL g190 ( .A1(n_162), .A2(n_155), .B1(n_154), .B2(n_125), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_168), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_176), .B(n_150), .Y(n_192) );
INVx2_ASAP7_75t_SL g193 ( .A(n_176), .Y(n_193) );
XNOR2xp5_ASAP7_75t_L g194 ( .A(n_158), .B(n_144), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_176), .B(n_150), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_170), .Y(n_196) );
AO22x2_ASAP7_75t_L g197 ( .A1(n_177), .A2(n_143), .B1(n_128), .B2(n_151), .Y(n_197) );
OAI22xp33_ASAP7_75t_L g198 ( .A1(n_179), .A2(n_150), .B1(n_145), .B2(n_153), .Y(n_198) );
OAI22xp33_ASAP7_75t_L g199 ( .A1(n_179), .A2(n_154), .B1(n_151), .B2(n_125), .Y(n_199) );
NAND3x1_ASAP7_75t_L g200 ( .A(n_158), .B(n_128), .C(n_131), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_158), .A2(n_131), .B1(n_143), .B2(n_147), .Y(n_201) );
AO22x2_ASAP7_75t_L g202 ( .A1(n_177), .A2(n_130), .B1(n_5), .B2(n_6), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_156), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_156), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_176), .B(n_112), .Y(n_205) );
OAI22xp5_ASAP7_75t_SL g206 ( .A1(n_170), .A2(n_149), .B1(n_148), .B2(n_146), .Y(n_206) );
OAI22xp33_ASAP7_75t_SL g207 ( .A1(n_162), .A2(n_142), .B1(n_140), .B2(n_139), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_156), .Y(n_208) );
OAI22xp5_ASAP7_75t_L g209 ( .A1(n_176), .A2(n_133), .B1(n_127), .B2(n_122), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_161), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_169), .A2(n_136), .B1(n_121), .B2(n_120), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g212 ( .A1(n_169), .A2(n_4), .B1(n_8), .B2(n_9), .Y(n_212) );
AO22x2_ASAP7_75t_L g213 ( .A1(n_177), .A2(n_4), .B1(n_8), .B2(n_10), .Y(n_213) );
OAI22xp33_ASAP7_75t_L g214 ( .A1(n_179), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_157), .B(n_34), .Y(n_215) );
OR2x2_ASAP7_75t_L g216 ( .A(n_157), .B(n_11), .Y(n_216) );
AO22x2_ASAP7_75t_L g217 ( .A1(n_177), .A2(n_13), .B1(n_15), .B2(n_16), .Y(n_217) );
HB1xp67_ASAP7_75t_L g218 ( .A(n_169), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_169), .B(n_13), .Y(n_219) );
OAI22xp33_ASAP7_75t_L g220 ( .A1(n_157), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_160), .Y(n_221) );
AND2x2_ASAP7_75t_L g222 ( .A(n_157), .B(n_17), .Y(n_222) );
BUFx3_ASAP7_75t_L g223 ( .A(n_164), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_171), .B(n_18), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_171), .B(n_19), .Y(n_225) );
INVxp67_ASAP7_75t_L g226 ( .A(n_171), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_171), .B(n_20), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_168), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_180), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_223), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_193), .A2(n_177), .B(n_164), .Y(n_231) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_223), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_192), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_195), .Y(n_234) );
INVx1_ASAP7_75t_SL g235 ( .A(n_219), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_181), .Y(n_236) );
INVx3_ASAP7_75t_L g237 ( .A(n_185), .Y(n_237) );
AND2x4_ASAP7_75t_L g238 ( .A(n_218), .B(n_189), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_203), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_204), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_208), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_218), .B(n_177), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_183), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_221), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_196), .Y(n_245) );
BUFx6f_ASAP7_75t_SL g246 ( .A(n_213), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_222), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_226), .B(n_177), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_196), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_206), .Y(n_250) );
INVxp33_ASAP7_75t_L g251 ( .A(n_182), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_222), .Y(n_252) );
CKINVDCx14_ASAP7_75t_R g253 ( .A(n_209), .Y(n_253) );
CKINVDCx14_ASAP7_75t_R g254 ( .A(n_211), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_216), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_201), .B(n_165), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_197), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_193), .A2(n_164), .B(n_160), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_197), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_197), .Y(n_260) );
CKINVDCx16_ASAP7_75t_R g261 ( .A(n_194), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_224), .Y(n_262) );
INVxp33_ASAP7_75t_L g263 ( .A(n_184), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_227), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_225), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_199), .B(n_160), .Y(n_266) );
XOR2xp5_ASAP7_75t_L g267 ( .A(n_198), .B(n_160), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_200), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_183), .Y(n_269) );
BUFx3_ASAP7_75t_L g270 ( .A(n_215), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_188), .Y(n_271) );
XOR2xp5_ASAP7_75t_L g272 ( .A(n_198), .B(n_160), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_200), .Y(n_273) );
AND2x6_ASAP7_75t_L g274 ( .A(n_215), .B(n_160), .Y(n_274) );
BUFx5_ASAP7_75t_L g275 ( .A(n_213), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_213), .Y(n_276) );
AND2x6_ASAP7_75t_L g277 ( .A(n_212), .B(n_160), .Y(n_277) );
NOR2xp33_ASAP7_75t_SL g278 ( .A(n_220), .B(n_165), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_217), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_217), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_217), .Y(n_281) );
XOR2xp5_ASAP7_75t_L g282 ( .A(n_207), .B(n_20), .Y(n_282) );
OAI21xp5_ASAP7_75t_L g283 ( .A1(n_188), .A2(n_164), .B(n_178), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_191), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_199), .B(n_164), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_187), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_190), .Y(n_287) );
INVxp33_ASAP7_75t_SL g288 ( .A(n_186), .Y(n_288) );
INVxp33_ASAP7_75t_SL g289 ( .A(n_202), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_202), .B(n_166), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_202), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_205), .B(n_166), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_220), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_191), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_243), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_255), .B(n_247), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_243), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_269), .Y(n_298) );
BUFx5_ASAP7_75t_L g299 ( .A(n_257), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_252), .B(n_214), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_269), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_237), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_287), .B(n_214), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_238), .B(n_178), .Y(n_304) );
AND2x6_ASAP7_75t_L g305 ( .A(n_259), .B(n_174), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_286), .B(n_228), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_271), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_256), .B(n_228), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_267), .B(n_168), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_267), .B(n_168), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_272), .B(n_168), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_271), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_275), .B(n_174), .Y(n_313) );
INVxp67_ASAP7_75t_L g314 ( .A(n_238), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_284), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_237), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_263), .B(n_21), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_237), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_244), .B(n_174), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_272), .B(n_21), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_284), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_232), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_238), .B(n_260), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_263), .B(n_22), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_276), .B(n_22), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_294), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_244), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_275), .B(n_23), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_275), .B(n_23), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_262), .B(n_174), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_294), .Y(n_331) );
AND2x4_ASAP7_75t_L g332 ( .A(n_279), .B(n_24), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_275), .B(n_24), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_275), .B(n_25), .Y(n_334) );
BUFx3_ASAP7_75t_L g335 ( .A(n_232), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_232), .Y(n_336) );
INVx2_ASAP7_75t_SL g337 ( .A(n_232), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_275), .B(n_26), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_232), .Y(n_339) );
BUFx3_ASAP7_75t_L g340 ( .A(n_275), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_230), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_290), .B(n_26), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_230), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_229), .Y(n_344) );
INVx2_ASAP7_75t_SL g345 ( .A(n_270), .Y(n_345) );
INVx4_ASAP7_75t_L g346 ( .A(n_246), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_290), .B(n_27), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_235), .B(n_28), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_280), .B(n_28), .Y(n_349) );
BUFx8_ASAP7_75t_L g350 ( .A(n_320), .Y(n_350) );
NOR2xp33_ASAP7_75t_SL g351 ( .A(n_346), .B(n_246), .Y(n_351) );
NOR2xp33_ASAP7_75t_SL g352 ( .A(n_346), .B(n_246), .Y(n_352) );
INVx1_ASAP7_75t_SL g353 ( .A(n_328), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_346), .B(n_323), .Y(n_354) );
BUFx4f_ASAP7_75t_L g355 ( .A(n_323), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_327), .B(n_293), .Y(n_356) );
CKINVDCx8_ASAP7_75t_R g357 ( .A(n_305), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_320), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_327), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_327), .B(n_277), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_314), .B(n_288), .Y(n_361) );
BUFx3_ASAP7_75t_L g362 ( .A(n_322), .Y(n_362) );
BUFx12f_ASAP7_75t_L g363 ( .A(n_346), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_320), .B(n_265), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_326), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_326), .Y(n_366) );
AND2x6_ASAP7_75t_L g367 ( .A(n_340), .B(n_281), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_314), .B(n_288), .Y(n_368) );
INVx2_ASAP7_75t_SL g369 ( .A(n_326), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_320), .B(n_264), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_296), .B(n_251), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_344), .B(n_277), .Y(n_372) );
OR2x6_ASAP7_75t_L g373 ( .A(n_346), .B(n_268), .Y(n_373) );
NAND2x1p5_ASAP7_75t_L g374 ( .A(n_346), .B(n_236), .Y(n_374) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_322), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_323), .B(n_273), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_326), .B(n_266), .Y(n_377) );
INVx5_ASAP7_75t_L g378 ( .A(n_305), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_331), .Y(n_379) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_322), .Y(n_380) );
CKINVDCx6p67_ASAP7_75t_R g381 ( .A(n_325), .Y(n_381) );
BUFx12f_ASAP7_75t_L g382 ( .A(n_325), .Y(n_382) );
AND2x2_ASAP7_75t_SL g383 ( .A(n_328), .B(n_291), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_379), .Y(n_384) );
BUFx2_ASAP7_75t_L g385 ( .A(n_382), .Y(n_385) );
BUFx4_ASAP7_75t_SL g386 ( .A(n_379), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_365), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_359), .B(n_344), .Y(n_388) );
INVx3_ASAP7_75t_L g389 ( .A(n_365), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_365), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_350), .Y(n_391) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_375), .Y(n_392) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_375), .Y(n_393) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_375), .Y(n_394) );
BUFx3_ASAP7_75t_L g395 ( .A(n_363), .Y(n_395) );
INVxp67_ASAP7_75t_L g396 ( .A(n_366), .Y(n_396) );
INVx1_ASAP7_75t_SL g397 ( .A(n_366), .Y(n_397) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_375), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_366), .Y(n_399) );
BUFx3_ASAP7_75t_L g400 ( .A(n_363), .Y(n_400) );
BUFx12f_ASAP7_75t_L g401 ( .A(n_350), .Y(n_401) );
INVx1_ASAP7_75t_SL g402 ( .A(n_381), .Y(n_402) );
BUFx3_ASAP7_75t_L g403 ( .A(n_363), .Y(n_403) );
NAND2x1p5_ASAP7_75t_L g404 ( .A(n_369), .B(n_340), .Y(n_404) );
BUFx12f_ASAP7_75t_L g405 ( .A(n_350), .Y(n_405) );
BUFx10_ASAP7_75t_L g406 ( .A(n_354), .Y(n_406) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_375), .Y(n_407) );
BUFx2_ASAP7_75t_L g408 ( .A(n_382), .Y(n_408) );
INVx5_ASAP7_75t_L g409 ( .A(n_382), .Y(n_409) );
INVx2_ASAP7_75t_SL g410 ( .A(n_355), .Y(n_410) );
CKINVDCx16_ASAP7_75t_R g411 ( .A(n_351), .Y(n_411) );
BUFx5_ASAP7_75t_L g412 ( .A(n_367), .Y(n_412) );
INVx3_ASAP7_75t_L g413 ( .A(n_375), .Y(n_413) );
BUFx2_ASAP7_75t_SL g414 ( .A(n_386), .Y(n_414) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_392), .Y(n_415) );
OAI22xp33_ASAP7_75t_L g416 ( .A1(n_409), .A2(n_289), .B1(n_381), .B2(n_353), .Y(n_416) );
BUFx12f_ASAP7_75t_L g417 ( .A(n_401), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_401), .A2(n_289), .B1(n_350), .B2(n_371), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_384), .Y(n_419) );
BUFx2_ASAP7_75t_SL g420 ( .A(n_386), .Y(n_420) );
BUFx2_ASAP7_75t_L g421 ( .A(n_397), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_411), .A2(n_353), .B1(n_383), .B2(n_358), .Y(n_422) );
NAND2x1p5_ASAP7_75t_L g423 ( .A(n_397), .B(n_369), .Y(n_423) );
CKINVDCx11_ASAP7_75t_R g424 ( .A(n_401), .Y(n_424) );
CKINVDCx11_ASAP7_75t_R g425 ( .A(n_405), .Y(n_425) );
BUFx3_ASAP7_75t_L g426 ( .A(n_395), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_399), .Y(n_427) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_405), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_384), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_399), .Y(n_430) );
BUFx12f_ASAP7_75t_L g431 ( .A(n_405), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_399), .Y(n_432) );
INVx6_ASAP7_75t_L g433 ( .A(n_406), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_409), .A2(n_277), .B1(n_317), .B2(n_324), .Y(n_434) );
BUFx2_ASAP7_75t_L g435 ( .A(n_396), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_388), .B(n_377), .Y(n_436) );
INVx1_ASAP7_75t_SL g437 ( .A(n_402), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_387), .Y(n_438) );
INVx6_ASAP7_75t_L g439 ( .A(n_406), .Y(n_439) );
BUFx3_ASAP7_75t_L g440 ( .A(n_395), .Y(n_440) );
BUFx4f_ASAP7_75t_SL g441 ( .A(n_395), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_411), .A2(n_383), .B1(n_357), .B2(n_347), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_409), .A2(n_383), .B1(n_357), .B2(n_347), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_391), .Y(n_444) );
INVx3_ASAP7_75t_L g445 ( .A(n_404), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_387), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_390), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_390), .B(n_359), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_396), .B(n_370), .Y(n_449) );
BUFx8_ASAP7_75t_SL g450 ( .A(n_400), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_388), .Y(n_451) );
BUFx4_ASAP7_75t_R g452 ( .A(n_412), .Y(n_452) );
OAI22xp33_ASAP7_75t_L g453 ( .A1(n_409), .A2(n_352), .B1(n_351), .B2(n_385), .Y(n_453) );
INVx2_ASAP7_75t_SL g454 ( .A(n_406), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_389), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_409), .A2(n_277), .B1(n_317), .B2(n_324), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_409), .A2(n_277), .B1(n_370), .B2(n_364), .Y(n_457) );
BUFx2_ASAP7_75t_L g458 ( .A(n_412), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_389), .Y(n_459) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_415), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_422), .A2(n_277), .B1(n_364), .B2(n_282), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_424), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_422), .A2(n_420), .B1(n_414), .B2(n_457), .Y(n_463) );
OAI22xp33_ASAP7_75t_L g464 ( .A1(n_441), .A2(n_409), .B1(n_352), .B2(n_385), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_419), .Y(n_465) );
NOR2x1_ASAP7_75t_SL g466 ( .A(n_414), .B(n_409), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_420), .A2(n_282), .B1(n_347), .B2(n_342), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_417), .B(n_261), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_457), .A2(n_342), .B1(n_347), .B2(n_408), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_419), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_438), .B(n_389), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_443), .A2(n_408), .B1(n_385), .B2(n_402), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_442), .A2(n_342), .B1(n_408), .B2(n_361), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_417), .B(n_250), .Y(n_474) );
BUFx12f_ASAP7_75t_L g475 ( .A(n_424), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_448), .B(n_342), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_429), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_427), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_429), .Y(n_479) );
INVx5_ASAP7_75t_SL g480 ( .A(n_425), .Y(n_480) );
BUFx4f_ASAP7_75t_SL g481 ( .A(n_417), .Y(n_481) );
BUFx10_ASAP7_75t_L g482 ( .A(n_433), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_443), .A2(n_410), .B1(n_400), .B2(n_403), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_442), .A2(n_410), .B1(n_400), .B2(n_403), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_434), .A2(n_368), .B1(n_310), .B2(n_309), .Y(n_485) );
AOI22xp33_ASAP7_75t_SL g486 ( .A1(n_433), .A2(n_403), .B1(n_410), .B2(n_412), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_416), .A2(n_278), .B1(n_311), .B2(n_309), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_438), .B(n_389), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_448), .B(n_349), .Y(n_489) );
BUFx3_ASAP7_75t_L g490 ( .A(n_441), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_438), .B(n_389), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_434), .A2(n_309), .B1(n_311), .B2(n_310), .Y(n_492) );
OAI22xp33_ASAP7_75t_L g493 ( .A1(n_431), .A2(n_355), .B1(n_374), .B2(n_372), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_427), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_456), .A2(n_309), .B1(n_311), .B2(n_310), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_446), .Y(n_496) );
OAI222xp33_ASAP7_75t_L g497 ( .A1(n_418), .A2(n_245), .B1(n_249), .B2(n_373), .C1(n_333), .C2(n_329), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_456), .A2(n_310), .B1(n_311), .B2(n_355), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_418), .A2(n_355), .B1(n_376), .B2(n_348), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_448), .B(n_349), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_416), .A2(n_376), .B1(n_348), .B2(n_372), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_446), .Y(n_502) );
BUFx3_ASAP7_75t_L g503 ( .A(n_450), .Y(n_503) );
BUFx4f_ASAP7_75t_SL g504 ( .A(n_431), .Y(n_504) );
BUFx12f_ASAP7_75t_L g505 ( .A(n_425), .Y(n_505) );
AOI22xp33_ASAP7_75t_SL g506 ( .A1(n_433), .A2(n_412), .B1(n_406), .B2(n_253), .Y(n_506) );
INVx1_ASAP7_75t_SL g507 ( .A(n_437), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_451), .A2(n_376), .B1(n_348), .B2(n_354), .Y(n_508) );
BUFx12f_ASAP7_75t_L g509 ( .A(n_444), .Y(n_509) );
AOI22xp33_ASAP7_75t_SL g510 ( .A1(n_433), .A2(n_412), .B1(n_406), .B2(n_253), .Y(n_510) );
OAI21xp5_ASAP7_75t_SL g511 ( .A1(n_453), .A2(n_374), .B(n_329), .Y(n_511) );
BUFx2_ASAP7_75t_L g512 ( .A(n_421), .Y(n_512) );
BUFx2_ASAP7_75t_L g513 ( .A(n_421), .Y(n_513) );
AOI22xp33_ASAP7_75t_SL g514 ( .A1(n_433), .A2(n_412), .B1(n_329), .B2(n_338), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_449), .A2(n_332), .B1(n_325), .B2(n_360), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_446), .B(n_413), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_449), .B(n_349), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_437), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_427), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_449), .B(n_349), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_447), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_447), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_447), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_450), .A2(n_325), .B1(n_332), .B2(n_333), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_430), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_436), .A2(n_325), .B1(n_332), .B2(n_333), .Y(n_526) );
OAI22xp33_ASAP7_75t_L g527 ( .A1(n_428), .A2(n_373), .B1(n_378), .B2(n_245), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_430), .B(n_413), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_439), .A2(n_334), .B1(n_329), .B2(n_338), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_436), .A2(n_332), .B1(n_325), .B2(n_334), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_461), .A2(n_473), .B1(n_463), .B2(n_467), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_487), .A2(n_440), .B1(n_426), .B2(n_458), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_487), .A2(n_440), .B1(n_426), .B2(n_458), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_498), .A2(n_440), .B1(n_426), .B2(n_458), .Y(n_534) );
AOI21xp5_ASAP7_75t_SL g535 ( .A1(n_466), .A2(n_453), .B(n_454), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_511), .A2(n_428), .B1(n_439), .B2(n_454), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_499), .A2(n_439), .B1(n_454), .B2(n_332), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_465), .B(n_435), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_511), .A2(n_439), .B1(n_435), .B2(n_445), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_469), .A2(n_439), .B1(n_334), .B2(n_338), .Y(n_540) );
AOI22xp33_ASAP7_75t_SL g541 ( .A1(n_466), .A2(n_445), .B1(n_435), .B2(n_412), .Y(n_541) );
OAI222xp33_ASAP7_75t_L g542 ( .A1(n_472), .A2(n_445), .B1(n_249), .B2(n_423), .C1(n_421), .C2(n_373), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_506), .A2(n_445), .B1(n_423), .B2(n_373), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_485), .A2(n_334), .B1(n_328), .B2(n_445), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_510), .A2(n_423), .B1(n_373), .B2(n_432), .Y(n_545) );
AOI22xp33_ASAP7_75t_SL g546 ( .A1(n_484), .A2(n_412), .B1(n_254), .B2(n_423), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_492), .A2(n_377), .B1(n_412), .B2(n_367), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_524), .A2(n_432), .B1(n_254), .B2(n_459), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_470), .B(n_432), .Y(n_549) );
AOI22xp33_ASAP7_75t_SL g550 ( .A1(n_483), .A2(n_504), .B1(n_481), .B2(n_480), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_495), .A2(n_412), .B1(n_367), .B2(n_303), .Y(n_551) );
NAND3xp33_ASAP7_75t_L g552 ( .A(n_514), .B(n_303), .C(n_173), .Y(n_552) );
AOI22xp33_ASAP7_75t_SL g553 ( .A1(n_480), .A2(n_412), .B1(n_452), .B2(n_250), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_501), .A2(n_412), .B1(n_367), .B2(n_303), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_527), .A2(n_367), .B1(n_455), .B2(n_459), .Y(n_555) );
NAND3xp33_ASAP7_75t_L g556 ( .A(n_477), .B(n_175), .C(n_173), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_496), .Y(n_557) );
AOI22xp33_ASAP7_75t_SL g558 ( .A1(n_480), .A2(n_452), .B1(n_413), .B2(n_378), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_529), .A2(n_367), .B1(n_356), .B2(n_362), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_503), .A2(n_367), .B1(n_362), .B2(n_300), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_503), .A2(n_367), .B1(n_362), .B2(n_300), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_508), .A2(n_344), .B1(n_251), .B2(n_296), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_476), .A2(n_304), .B1(n_274), .B2(n_305), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_517), .A2(n_304), .B1(n_274), .B2(n_305), .Y(n_564) );
BUFx3_ASAP7_75t_L g565 ( .A(n_490), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_526), .A2(n_404), .B1(n_378), .B2(n_296), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_530), .A2(n_378), .B1(n_413), .B2(n_340), .Y(n_567) );
AOI22xp33_ASAP7_75t_SL g568 ( .A1(n_480), .A2(n_413), .B1(n_378), .B2(n_415), .Y(n_568) );
OAI21xp5_ASAP7_75t_SL g569 ( .A1(n_497), .A2(n_304), .B(n_330), .Y(n_569) );
OAI222xp33_ASAP7_75t_L g570 ( .A1(n_486), .A2(n_378), .B1(n_330), .B2(n_304), .C1(n_313), .C2(n_340), .Y(n_570) );
NAND3xp33_ASAP7_75t_L g571 ( .A(n_479), .B(n_175), .C(n_167), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_520), .A2(n_304), .B1(n_274), .B2(n_305), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_496), .Y(n_573) );
OAI221xp5_ASAP7_75t_L g574 ( .A1(n_468), .A2(n_308), .B1(n_306), .B2(n_330), .C(n_292), .Y(n_574) );
NOR3xp33_ASAP7_75t_L g575 ( .A(n_474), .B(n_308), .C(n_167), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_490), .A2(n_304), .B1(n_274), .B2(n_305), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_502), .B(n_415), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_493), .A2(n_304), .B1(n_274), .B2(n_305), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_489), .A2(n_274), .B1(n_305), .B2(n_345), .Y(n_579) );
AOI22xp33_ASAP7_75t_SL g580 ( .A1(n_482), .A2(n_415), .B1(n_407), .B2(n_398), .Y(n_580) );
OA21x2_ASAP7_75t_L g581 ( .A1(n_502), .A2(n_319), .B(n_313), .Y(n_581) );
OAI22xp33_ASAP7_75t_L g582 ( .A1(n_475), .A2(n_415), .B1(n_407), .B2(n_398), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_464), .A2(n_331), .B1(n_345), .B2(n_394), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_500), .A2(n_305), .B1(n_345), .B2(n_380), .Y(n_584) );
AOI22xp33_ASAP7_75t_SL g585 ( .A1(n_482), .A2(n_407), .B1(n_398), .B2(n_394), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_515), .A2(n_331), .B1(n_398), .B2(n_394), .Y(n_586) );
NAND3xp33_ASAP7_75t_L g587 ( .A(n_462), .B(n_175), .C(n_167), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_475), .A2(n_305), .B1(n_380), .B2(n_299), .Y(n_588) );
OAI222xp33_ASAP7_75t_L g589 ( .A1(n_462), .A2(n_308), .B1(n_306), .B2(n_319), .C1(n_285), .C2(n_32), .Y(n_589) );
NOR2xp67_ASAP7_75t_L g590 ( .A(n_521), .B(n_392), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_505), .A2(n_407), .B1(n_398), .B2(n_394), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_505), .A2(n_305), .B1(n_380), .B2(n_299), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_507), .A2(n_305), .B1(n_380), .B2(n_299), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_507), .A2(n_380), .B1(n_299), .B2(n_323), .Y(n_594) );
AOI22xp33_ASAP7_75t_SL g595 ( .A1(n_482), .A2(n_407), .B1(n_398), .B2(n_394), .Y(n_595) );
INVxp67_ASAP7_75t_L g596 ( .A(n_518), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_518), .A2(n_299), .B1(n_323), .B2(n_394), .Y(n_597) );
OAI221xp5_ASAP7_75t_L g598 ( .A1(n_512), .A2(n_306), .B1(n_283), .B2(n_167), .C(n_173), .Y(n_598) );
OAI22xp33_ASAP7_75t_L g599 ( .A1(n_512), .A2(n_407), .B1(n_398), .B2(n_394), .Y(n_599) );
NAND3xp33_ASAP7_75t_L g600 ( .A(n_522), .B(n_175), .C(n_173), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_513), .A2(n_299), .B1(n_323), .B2(n_394), .Y(n_601) );
OAI221xp5_ASAP7_75t_SL g602 ( .A1(n_513), .A2(n_319), .B1(n_242), .B2(n_234), .C(n_233), .Y(n_602) );
OAI221xp5_ASAP7_75t_L g603 ( .A1(n_522), .A2(n_234), .B1(n_233), .B2(n_175), .C(n_241), .Y(n_603) );
OAI21xp5_ASAP7_75t_SL g604 ( .A1(n_523), .A2(n_174), .B(n_323), .Y(n_604) );
OAI22xp33_ASAP7_75t_L g605 ( .A1(n_509), .A2(n_407), .B1(n_398), .B2(n_393), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_516), .A2(n_299), .B1(n_393), .B2(n_392), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_516), .A2(n_299), .B1(n_393), .B2(n_392), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_523), .A2(n_407), .B1(n_393), .B2(n_392), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_471), .A2(n_299), .B1(n_321), .B2(n_298), .Y(n_609) );
AOI222xp33_ASAP7_75t_L g610 ( .A1(n_509), .A2(n_174), .B1(n_175), .B2(n_239), .C1(n_240), .C2(n_172), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_478), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_478), .A2(n_393), .B1(n_392), .B2(n_307), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_471), .A2(n_299), .B1(n_392), .B2(n_393), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_488), .A2(n_299), .B1(n_393), .B2(n_322), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_488), .A2(n_299), .B1(n_298), .B2(n_301), .Y(n_615) );
AOI22xp33_ASAP7_75t_SL g616 ( .A1(n_491), .A2(n_393), .B1(n_335), .B2(n_174), .Y(n_616) );
AOI22xp33_ASAP7_75t_SL g617 ( .A1(n_491), .A2(n_528), .B1(n_525), .B2(n_519), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_494), .A2(n_301), .B1(n_297), .B2(n_307), .Y(n_618) );
OAI221xp5_ASAP7_75t_SL g619 ( .A1(n_494), .A2(n_258), .B1(n_248), .B2(n_312), .C(n_295), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_519), .A2(n_299), .B1(n_335), .B2(n_337), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_460), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_460), .A2(n_337), .B1(n_270), .B2(n_339), .Y(n_622) );
AOI22xp33_ASAP7_75t_SL g623 ( .A1(n_460), .A2(n_174), .B1(n_297), .B2(n_312), .Y(n_623) );
AND2x6_ASAP7_75t_L g624 ( .A(n_536), .B(n_460), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_538), .B(n_460), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_596), .B(n_29), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_538), .B(n_29), .Y(n_627) );
NAND3xp33_ASAP7_75t_L g628 ( .A(n_550), .B(n_175), .C(n_172), .Y(n_628) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_531), .A2(n_175), .B1(n_174), .B2(n_172), .C(n_161), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_536), .A2(n_307), .B1(n_295), .B2(n_301), .Y(n_630) );
OAI21xp5_ASAP7_75t_SL g631 ( .A1(n_542), .A2(n_174), .B(n_175), .Y(n_631) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_589), .A2(n_175), .B1(n_172), .B2(n_161), .C(n_163), .Y(n_632) );
OAI21xp5_ASAP7_75t_SL g633 ( .A1(n_569), .A2(n_161), .B(n_172), .Y(n_633) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_574), .A2(n_161), .B1(n_172), .B2(n_163), .C(n_231), .Y(n_634) );
OAI21xp5_ASAP7_75t_SL g635 ( .A1(n_553), .A2(n_161), .B(n_172), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_573), .B(n_30), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_549), .B(n_30), .Y(n_637) );
OAI211xp5_ASAP7_75t_L g638 ( .A1(n_535), .A2(n_161), .B(n_172), .C(n_163), .Y(n_638) );
AOI221xp5_ASAP7_75t_L g639 ( .A1(n_575), .A2(n_161), .B1(n_172), .B2(n_163), .C(n_302), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_549), .B(n_31), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_617), .B(n_32), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_557), .B(n_33), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_577), .B(n_163), .Y(n_643) );
NAND3xp33_ASAP7_75t_L g644 ( .A(n_610), .B(n_163), .C(n_336), .Y(n_644) );
OAI21xp33_ASAP7_75t_L g645 ( .A1(n_535), .A2(n_339), .B(n_336), .Y(n_645) );
OAI221xp5_ASAP7_75t_L g646 ( .A1(n_604), .A2(n_163), .B1(n_302), .B2(n_316), .C(n_318), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_565), .B(n_163), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_611), .B(n_163), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_565), .B(n_163), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_539), .B(n_35), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_611), .B(n_312), .Y(n_651) );
AND2x2_ASAP7_75t_SL g652 ( .A(n_532), .B(n_315), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_548), .A2(n_339), .B1(n_336), .B2(n_343), .Y(n_653) );
NAND3xp33_ASAP7_75t_L g654 ( .A(n_587), .B(n_343), .C(n_341), .Y(n_654) );
NAND3xp33_ASAP7_75t_L g655 ( .A(n_546), .B(n_343), .C(n_341), .Y(n_655) );
NAND3xp33_ASAP7_75t_L g656 ( .A(n_533), .B(n_343), .C(n_341), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_562), .B(n_301), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_590), .B(n_36), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_562), .B(n_321), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_534), .B(n_37), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_552), .A2(n_341), .B1(n_321), .B2(n_295), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_543), .B(n_321), .Y(n_662) );
INVxp67_ASAP7_75t_SL g663 ( .A(n_605), .Y(n_663) );
NAND3xp33_ASAP7_75t_L g664 ( .A(n_602), .B(n_295), .C(n_315), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_541), .B(n_40), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_545), .B(n_315), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_580), .B(n_43), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_585), .B(n_45), .Y(n_668) );
NAND2xp5_ASAP7_75t_SL g669 ( .A(n_582), .B(n_307), .Y(n_669) );
NAND3xp33_ASAP7_75t_L g670 ( .A(n_619), .B(n_298), .C(n_297), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_595), .B(n_46), .Y(n_671) );
AOI221xp5_ASAP7_75t_L g672 ( .A1(n_603), .A2(n_318), .B1(n_316), .B2(n_302), .C(n_298), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_591), .B(n_609), .Y(n_673) );
NOR3xp33_ASAP7_75t_L g674 ( .A(n_552), .B(n_318), .C(n_316), .Y(n_674) );
OA21x2_ASAP7_75t_L g675 ( .A1(n_608), .A2(n_297), .B(n_49), .Y(n_675) );
NAND3xp33_ASAP7_75t_L g676 ( .A(n_616), .B(n_210), .C(n_50), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_615), .B(n_48), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_615), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_601), .B(n_52), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_606), .B(n_54), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_559), .A2(n_57), .B1(n_60), .B2(n_61), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_607), .B(n_62), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_618), .Y(n_683) );
NOR3xp33_ASAP7_75t_SL g684 ( .A(n_570), .B(n_63), .C(n_64), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_544), .A2(n_210), .B1(n_68), .B2(n_69), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_613), .B(n_66), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_598), .B(n_70), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_555), .A2(n_71), .B1(n_72), .B2(n_73), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_560), .B(n_76), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_540), .B(n_77), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_537), .A2(n_210), .B1(n_80), .B2(n_81), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_561), .A2(n_558), .B1(n_547), .B2(n_551), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_554), .A2(n_210), .B1(n_82), .B2(n_83), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_597), .B(n_78), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_614), .B(n_86), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_586), .B(n_89), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_594), .B(n_90), .Y(n_697) );
NAND2xp5_ASAP7_75t_SL g698 ( .A(n_599), .B(n_92), .Y(n_698) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_612), .Y(n_699) );
OAI22xp33_ASAP7_75t_L g700 ( .A1(n_566), .A2(n_93), .B1(n_94), .B2(n_97), .Y(n_700) );
OAI21xp5_ASAP7_75t_SL g701 ( .A1(n_568), .A2(n_99), .B(n_101), .Y(n_701) );
NAND4xp25_ASAP7_75t_L g702 ( .A(n_578), .B(n_102), .C(n_108), .D(n_109), .Y(n_702) );
NAND3xp33_ASAP7_75t_L g703 ( .A(n_623), .B(n_110), .C(n_556), .Y(n_703) );
NAND3xp33_ASAP7_75t_L g704 ( .A(n_571), .B(n_588), .C(n_592), .Y(n_704) );
NOR3xp33_ASAP7_75t_L g705 ( .A(n_600), .B(n_583), .C(n_567), .Y(n_705) );
OAI221xp5_ASAP7_75t_SL g706 ( .A1(n_563), .A2(n_564), .B1(n_572), .B2(n_576), .C(n_579), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_620), .A2(n_581), .B1(n_593), .B2(n_584), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_622), .B(n_596), .Y(n_708) );
NAND3xp33_ASAP7_75t_L g709 ( .A(n_596), .B(n_550), .C(n_610), .Y(n_709) );
OA21x2_ASAP7_75t_L g710 ( .A1(n_621), .A2(n_511), .B(n_536), .Y(n_710) );
OA21x2_ASAP7_75t_L g711 ( .A1(n_621), .A2(n_511), .B(n_536), .Y(n_711) );
OAI221xp5_ASAP7_75t_SL g712 ( .A1(n_633), .A2(n_631), .B1(n_701), .B2(n_635), .C(n_709), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_699), .B(n_663), .Y(n_713) );
OR2x6_ASAP7_75t_L g714 ( .A(n_645), .B(n_698), .Y(n_714) );
INVx2_ASAP7_75t_SL g715 ( .A(n_647), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_692), .A2(n_652), .B1(n_678), .B2(n_624), .Y(n_716) );
NOR3xp33_ASAP7_75t_L g717 ( .A(n_641), .B(n_626), .C(n_702), .Y(n_717) );
NAND4xp75_ASAP7_75t_L g718 ( .A(n_652), .B(n_684), .C(n_710), .D(n_711), .Y(n_718) );
AND2x2_ASAP7_75t_L g719 ( .A(n_711), .B(n_673), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_642), .Y(n_720) );
AO21x2_ASAP7_75t_L g721 ( .A1(n_636), .A2(n_627), .B(n_643), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_704), .A2(n_644), .B1(n_683), .B2(n_705), .Y(n_722) );
AOI22xp5_ASAP7_75t_L g723 ( .A1(n_624), .A2(n_650), .B1(n_708), .B2(n_674), .Y(n_723) );
OR2x2_ASAP7_75t_L g724 ( .A(n_625), .B(n_651), .Y(n_724) );
NAND3xp33_ASAP7_75t_L g725 ( .A(n_629), .B(n_684), .C(n_705), .Y(n_725) );
NAND4xp75_ASAP7_75t_L g726 ( .A(n_698), .B(n_665), .C(n_660), .D(n_667), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_637), .B(n_640), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_624), .B(n_666), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_706), .B(n_649), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_624), .B(n_658), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_674), .A2(n_632), .B1(n_662), .B2(n_707), .Y(n_731) );
NAND3xp33_ASAP7_75t_L g732 ( .A(n_628), .B(n_707), .C(n_669), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_679), .B(n_648), .Y(n_733) );
NAND3xp33_ASAP7_75t_L g734 ( .A(n_669), .B(n_656), .C(n_639), .Y(n_734) );
NAND3xp33_ASAP7_75t_L g735 ( .A(n_693), .B(n_675), .C(n_691), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_668), .B(n_671), .Y(n_736) );
NAND3xp33_ASAP7_75t_L g737 ( .A(n_693), .B(n_675), .C(n_691), .Y(n_737) );
AO21x2_ASAP7_75t_L g738 ( .A1(n_700), .A2(n_696), .B(n_677), .Y(n_738) );
AOI22xp33_ASAP7_75t_SL g739 ( .A1(n_675), .A2(n_646), .B1(n_655), .B2(n_638), .Y(n_739) );
NAND3xp33_ASAP7_75t_L g740 ( .A(n_687), .B(n_654), .C(n_685), .Y(n_740) );
NAND3xp33_ASAP7_75t_L g741 ( .A(n_687), .B(n_685), .C(n_634), .Y(n_741) );
OR2x2_ASAP7_75t_SL g742 ( .A(n_676), .B(n_664), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_690), .B(n_694), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_695), .A2(n_697), .B1(n_689), .B2(n_630), .Y(n_744) );
NAND3xp33_ASAP7_75t_L g745 ( .A(n_670), .B(n_703), .C(n_680), .Y(n_745) );
AND2x4_ASAP7_75t_L g746 ( .A(n_657), .B(n_659), .Y(n_746) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_682), .B(n_686), .Y(n_747) );
NOR3xp33_ASAP7_75t_SL g748 ( .A(n_700), .B(n_681), .C(n_688), .Y(n_748) );
BUFx3_ASAP7_75t_L g749 ( .A(n_661), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_653), .B(n_672), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_709), .A2(n_692), .B1(n_633), .B2(n_536), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_709), .A2(n_531), .B1(n_461), .B2(n_575), .Y(n_752) );
NAND3xp33_ASAP7_75t_L g753 ( .A(n_709), .B(n_631), .C(n_633), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_709), .A2(n_531), .B1(n_461), .B2(n_575), .Y(n_754) );
NAND3xp33_ASAP7_75t_L g755 ( .A(n_709), .B(n_631), .C(n_633), .Y(n_755) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_626), .B(n_475), .Y(n_756) );
NAND3xp33_ASAP7_75t_L g757 ( .A(n_709), .B(n_631), .C(n_633), .Y(n_757) );
NAND3xp33_ASAP7_75t_L g758 ( .A(n_709), .B(n_631), .C(n_633), .Y(n_758) );
INVxp67_ASAP7_75t_L g759 ( .A(n_663), .Y(n_759) );
NOR3xp33_ASAP7_75t_L g760 ( .A(n_633), .B(n_631), .C(n_709), .Y(n_760) );
OA211x2_ASAP7_75t_L g761 ( .A1(n_645), .A2(n_698), .B(n_709), .C(n_463), .Y(n_761) );
NAND3xp33_ASAP7_75t_L g762 ( .A(n_709), .B(n_631), .C(n_633), .Y(n_762) );
INVx2_ASAP7_75t_SL g763 ( .A(n_647), .Y(n_763) );
NAND4xp75_ASAP7_75t_L g764 ( .A(n_652), .B(n_536), .C(n_684), .D(n_641), .Y(n_764) );
NAND3xp33_ASAP7_75t_L g765 ( .A(n_709), .B(n_631), .C(n_633), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_626), .B(n_475), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_626), .B(n_475), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_759), .B(n_719), .Y(n_768) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_759), .Y(n_769) );
NAND4xp75_ASAP7_75t_L g770 ( .A(n_761), .B(n_751), .C(n_716), .D(n_748), .Y(n_770) );
NAND4xp75_ASAP7_75t_L g771 ( .A(n_748), .B(n_723), .C(n_766), .D(n_756), .Y(n_771) );
INVx2_ASAP7_75t_SL g772 ( .A(n_715), .Y(n_772) );
INVx1_ASAP7_75t_SL g773 ( .A(n_713), .Y(n_773) );
BUFx2_ASAP7_75t_L g774 ( .A(n_714), .Y(n_774) );
XNOR2xp5_ASAP7_75t_L g775 ( .A(n_726), .B(n_736), .Y(n_775) );
NOR2xp33_ASAP7_75t_L g776 ( .A(n_729), .B(n_767), .Y(n_776) );
NAND4xp75_ASAP7_75t_L g777 ( .A(n_747), .B(n_743), .C(n_750), .D(n_720), .Y(n_777) );
NAND4xp75_ASAP7_75t_SL g778 ( .A(n_730), .B(n_718), .C(n_764), .D(n_712), .Y(n_778) );
NAND3xp33_ASAP7_75t_SL g779 ( .A(n_760), .B(n_755), .C(n_765), .Y(n_779) );
NAND4xp75_ASAP7_75t_SL g780 ( .A(n_753), .B(n_757), .C(n_762), .D(n_758), .Y(n_780) );
INVx2_ASAP7_75t_SL g781 ( .A(n_763), .Y(n_781) );
AND2x2_ASAP7_75t_L g782 ( .A(n_746), .B(n_728), .Y(n_782) );
INVx4_ASAP7_75t_L g783 ( .A(n_714), .Y(n_783) );
OAI31xp33_ASAP7_75t_L g784 ( .A1(n_735), .A2(n_737), .A3(n_732), .B(n_740), .Y(n_784) );
NOR2x1_ASAP7_75t_L g785 ( .A(n_714), .B(n_734), .Y(n_785) );
INVx1_ASAP7_75t_SL g786 ( .A(n_724), .Y(n_786) );
XOR2xp5_ASAP7_75t_L g787 ( .A(n_752), .B(n_754), .Y(n_787) );
XNOR2x2_ASAP7_75t_L g788 ( .A(n_725), .B(n_741), .Y(n_788) );
BUFx2_ASAP7_75t_L g789 ( .A(n_721), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_749), .Y(n_790) );
INVx1_ASAP7_75t_SL g791 ( .A(n_742), .Y(n_791) );
AOI22xp5_ASAP7_75t_L g792 ( .A1(n_752), .A2(n_754), .B1(n_722), .B2(n_717), .Y(n_792) );
NAND4xp75_ASAP7_75t_L g793 ( .A(n_733), .B(n_727), .C(n_722), .D(n_739), .Y(n_793) );
NAND4xp75_ASAP7_75t_L g794 ( .A(n_739), .B(n_717), .C(n_731), .D(n_738), .Y(n_794) );
AND2x2_ASAP7_75t_L g795 ( .A(n_738), .B(n_744), .Y(n_795) );
HB1xp67_ASAP7_75t_L g796 ( .A(n_769), .Y(n_796) );
OAI22x1_ASAP7_75t_L g797 ( .A1(n_774), .A2(n_731), .B1(n_745), .B2(n_783), .Y(n_797) );
XNOR2xp5_ASAP7_75t_L g798 ( .A(n_787), .B(n_775), .Y(n_798) );
AND2x2_ASAP7_75t_L g799 ( .A(n_774), .B(n_782), .Y(n_799) );
XOR2x2_ASAP7_75t_L g800 ( .A(n_780), .B(n_787), .Y(n_800) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_783), .A2(n_785), .B1(n_793), .B2(n_771), .Y(n_801) );
INVxp67_ASAP7_75t_L g802 ( .A(n_785), .Y(n_802) );
BUFx3_ASAP7_75t_L g803 ( .A(n_772), .Y(n_803) );
INVx3_ASAP7_75t_L g804 ( .A(n_783), .Y(n_804) );
HB1xp67_ASAP7_75t_SL g805 ( .A(n_783), .Y(n_805) );
XNOR2x1_ASAP7_75t_L g806 ( .A(n_794), .B(n_793), .Y(n_806) );
XNOR2xp5_ASAP7_75t_L g807 ( .A(n_775), .B(n_778), .Y(n_807) );
INVxp67_ASAP7_75t_L g808 ( .A(n_776), .Y(n_808) );
XNOR2xp5_ASAP7_75t_L g809 ( .A(n_792), .B(n_770), .Y(n_809) );
INVx1_ASAP7_75t_SL g810 ( .A(n_786), .Y(n_810) );
BUFx3_ASAP7_75t_L g811 ( .A(n_781), .Y(n_811) );
CKINVDCx16_ASAP7_75t_R g812 ( .A(n_779), .Y(n_812) );
HB1xp67_ASAP7_75t_L g813 ( .A(n_796), .Y(n_813) );
INVxp67_ASAP7_75t_L g814 ( .A(n_809), .Y(n_814) );
AOI22x1_ASAP7_75t_L g815 ( .A1(n_797), .A2(n_791), .B1(n_788), .B2(n_795), .Y(n_815) );
HB1xp67_ASAP7_75t_L g816 ( .A(n_810), .Y(n_816) );
XNOR2x1_ASAP7_75t_L g817 ( .A(n_806), .B(n_794), .Y(n_817) );
OA22x2_ASAP7_75t_L g818 ( .A1(n_809), .A2(n_791), .B1(n_792), .B2(n_795), .Y(n_818) );
HB1xp67_ASAP7_75t_L g819 ( .A(n_803), .Y(n_819) );
XOR2x2_ASAP7_75t_L g820 ( .A(n_800), .B(n_788), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_799), .Y(n_821) );
INVx4_ASAP7_75t_L g822 ( .A(n_804), .Y(n_822) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_805), .A2(n_777), .B1(n_790), .B2(n_768), .Y(n_823) );
AOI22x1_ASAP7_75t_L g824 ( .A1(n_797), .A2(n_784), .B1(n_789), .B2(n_773), .Y(n_824) );
OAI322xp33_ASAP7_75t_L g825 ( .A1(n_818), .A2(n_812), .A3(n_806), .B1(n_801), .B2(n_798), .C1(n_802), .C2(n_807), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_813), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_816), .Y(n_827) );
BUFx2_ASAP7_75t_L g828 ( .A(n_819), .Y(n_828) );
AO22x1_ASAP7_75t_L g829 ( .A1(n_822), .A2(n_804), .B1(n_811), .B2(n_803), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_821), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_822), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_822), .Y(n_832) );
BUFx3_ASAP7_75t_L g833 ( .A(n_820), .Y(n_833) );
OAI22xp5_ASAP7_75t_L g834 ( .A1(n_833), .A2(n_817), .B1(n_818), .B2(n_807), .Y(n_834) );
OAI322xp33_ASAP7_75t_L g835 ( .A1(n_827), .A2(n_818), .A3(n_814), .B1(n_817), .B2(n_815), .C1(n_824), .C2(n_798), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_828), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_833), .A2(n_823), .B1(n_815), .B2(n_824), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_828), .Y(n_838) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_834), .A2(n_837), .B1(n_827), .B2(n_832), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_836), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_838), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_840), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_839), .B(n_820), .Y(n_843) );
NAND3xp33_ASAP7_75t_SL g844 ( .A(n_843), .B(n_841), .C(n_831), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_842), .Y(n_845) );
INVx2_ASAP7_75t_L g846 ( .A(n_845), .Y(n_846) );
INVx2_ASAP7_75t_L g847 ( .A(n_844), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_847), .Y(n_848) );
BUFx2_ASAP7_75t_L g849 ( .A(n_846), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_849), .Y(n_850) );
INVxp67_ASAP7_75t_L g851 ( .A(n_850), .Y(n_851) );
AOI22xp5_ASAP7_75t_L g852 ( .A1(n_851), .A2(n_848), .B1(n_849), .B2(n_800), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_852), .Y(n_853) );
AOI22xp5_ASAP7_75t_L g854 ( .A1(n_853), .A2(n_826), .B1(n_808), .B2(n_830), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_854), .Y(n_855) );
AOI221x1_ASAP7_75t_L g856 ( .A1(n_855), .A2(n_826), .B1(n_835), .B2(n_825), .C(n_829), .Y(n_856) );
AOI211xp5_ASAP7_75t_L g857 ( .A1(n_856), .A2(n_829), .B(n_799), .C(n_811), .Y(n_857) );
endmodule