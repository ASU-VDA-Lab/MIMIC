module fake_ibex_1026_n_957 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_181, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_957);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_957;

wire n_599;
wire n_822;
wire n_778;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_926;
wire n_328;
wire n_293;
wire n_372;
wire n_341;
wire n_418;
wire n_256;
wire n_510;
wire n_193;
wire n_845;
wire n_947;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_375;
wire n_317;
wire n_340;
wire n_708;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_259;
wire n_339;
wire n_276;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_798;
wire n_732;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_953;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_949;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_837;
wire n_797;
wire n_796;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_402;
wire n_725;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_444;
wire n_200;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_927;
wire n_684;
wire n_775;
wire n_934;
wire n_784;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_285;
wire n_247;
wire n_320;
wire n_379;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_820;
wire n_728;
wire n_670;
wire n_805;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_683;
wire n_631;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_897;
wire n_889;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_912;
wire n_921;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_175),
.Y(n_182)
);

INVxp67_ASAP7_75t_SL g183 ( 
.A(n_144),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_53),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_16),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_3),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_32),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_126),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_56),
.Y(n_189)
);

INVxp33_ASAP7_75t_SL g190 ( 
.A(n_47),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_64),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_48),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_96),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_12),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_157),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_121),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_5),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_12),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_43),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_92),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_91),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_42),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_94),
.Y(n_206)
);

NOR2xp67_ASAP7_75t_L g207 ( 
.A(n_117),
.B(n_78),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_90),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_141),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_127),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_33),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_14),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_4),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_61),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_97),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_37),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_28),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_54),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_95),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_11),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_137),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_132),
.Y(n_223)
);

INVxp33_ASAP7_75t_L g224 ( 
.A(n_21),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_116),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_123),
.Y(n_226)
);

BUFx10_ASAP7_75t_L g227 ( 
.A(n_75),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_178),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_149),
.B(n_32),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_156),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_136),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_30),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_151),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_179),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_49),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_41),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_150),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_155),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_0),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_128),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_146),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_17),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_77),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_118),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_69),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_122),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_27),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_27),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_100),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_60),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_36),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_14),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_41),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_120),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_11),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_43),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_135),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_88),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_21),
.Y(n_259)
);

INVxp67_ASAP7_75t_SL g260 ( 
.A(n_36),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_5),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_28),
.Y(n_262)
);

NOR2xp67_ASAP7_75t_L g263 ( 
.A(n_71),
.B(n_163),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_152),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_142),
.B(n_25),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_30),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_170),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_161),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_158),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_74),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_153),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_37),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_70),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_81),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_134),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_171),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_160),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_85),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_139),
.Y(n_279)
);

BUFx8_ASAP7_75t_SL g280 ( 
.A(n_65),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_80),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_62),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_87),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_76),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_148),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_50),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_166),
.B(n_79),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_44),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_59),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_143),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_168),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_68),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_44),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_51),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_106),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_119),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_177),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_173),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_52),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_89),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_165),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_147),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_103),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_154),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_236),
.B(n_0),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_224),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_217),
.B(n_1),
.Y(n_307)
);

OAI22x1_ASAP7_75t_SL g308 ( 
.A1(n_186),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_182),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_189),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_224),
.B(n_6),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_198),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_288),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_280),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_225),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_230),
.B(n_7),
.Y(n_316)
);

OA21x2_ASAP7_75t_L g317 ( 
.A1(n_219),
.A2(n_86),
.B(n_176),
.Y(n_317)
);

AND2x4_ASAP7_75t_L g318 ( 
.A(n_214),
.B(n_261),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_219),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_182),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_221),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_214),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_261),
.Y(n_323)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_271),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_182),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_227),
.B(n_8),
.Y(n_326)
);

AND2x6_ASAP7_75t_L g327 ( 
.A(n_267),
.B(n_46),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_237),
.Y(n_328)
);

BUFx12f_ASAP7_75t_L g329 ( 
.A(n_227),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_293),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_182),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_210),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_184),
.B(n_188),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_210),
.Y(n_334)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_227),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_267),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_187),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_191),
.Y(n_338)
);

AND2x4_ASAP7_75t_L g339 ( 
.A(n_299),
.B(n_8),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_210),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_192),
.B(n_9),
.Y(n_341)
);

AND2x4_ASAP7_75t_L g342 ( 
.A(n_299),
.B(n_9),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_210),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_237),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_193),
.Y(n_345)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_185),
.Y(n_346)
);

AND2x4_ASAP7_75t_L g347 ( 
.A(n_268),
.B(n_10),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_281),
.B(n_55),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_185),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_200),
.Y(n_350)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_268),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_233),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_185),
.Y(n_353)
);

INVx5_ASAP7_75t_L g354 ( 
.A(n_220),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_195),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_277),
.Y(n_356)
);

AND2x4_ASAP7_75t_L g357 ( 
.A(n_277),
.B(n_10),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_197),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_213),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_185),
.Y(n_360)
);

AND2x4_ASAP7_75t_L g361 ( 
.A(n_218),
.B(n_13),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_199),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_190),
.A2(n_242),
.B1(n_195),
.B2(n_231),
.Y(n_363)
);

AND2x4_ASAP7_75t_L g364 ( 
.A(n_232),
.B(n_13),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_233),
.B(n_15),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_206),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_204),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_220),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_220),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_220),
.Y(n_370)
);

OA21x2_ASAP7_75t_L g371 ( 
.A1(n_208),
.A2(n_93),
.B(n_174),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_209),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_239),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_242),
.Y(n_374)
);

INVx5_ASAP7_75t_L g375 ( 
.A(n_190),
.Y(n_375)
);

AOI22x1_ASAP7_75t_SL g376 ( 
.A1(n_186),
.A2(n_272),
.B1(n_231),
.B2(n_274),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_248),
.B(n_16),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_252),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_338),
.B(n_211),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_L g380 ( 
.A1(n_347),
.A2(n_256),
.B1(n_255),
.B2(n_302),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_347),
.Y(n_381)
);

AND2x6_ASAP7_75t_L g382 ( 
.A(n_339),
.B(n_215),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_355),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_L g384 ( 
.A1(n_347),
.A2(n_235),
.B1(n_264),
.B2(n_301),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_339),
.B(n_216),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_339),
.B(n_222),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_338),
.B(n_223),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_324),
.B(n_238),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_L g389 ( 
.A1(n_357),
.A2(n_258),
.B1(n_226),
.B2(n_228),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_336),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_335),
.B(n_194),
.Y(n_391)
);

AND2x6_ASAP7_75t_L g392 ( 
.A(n_342),
.B(n_234),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_318),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_345),
.B(n_243),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_318),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_318),
.Y(n_396)
);

XNOR2x2_ASAP7_75t_SL g397 ( 
.A(n_363),
.B(n_272),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_357),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_357),
.Y(n_399)
);

OR2x2_ASAP7_75t_L g400 ( 
.A(n_313),
.B(n_260),
.Y(n_400)
);

OR2x6_ASAP7_75t_L g401 ( 
.A(n_329),
.B(n_265),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_361),
.Y(n_402)
);

AND2x6_ASAP7_75t_L g403 ( 
.A(n_342),
.B(n_245),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_314),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_355),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_324),
.B(n_269),
.Y(n_406)
);

OR2x6_ASAP7_75t_L g407 ( 
.A(n_329),
.B(n_229),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_372),
.Y(n_408)
);

AND2x6_ASAP7_75t_L g409 ( 
.A(n_342),
.B(n_246),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_374),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_361),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_324),
.B(n_284),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_335),
.B(n_292),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_309),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g415 ( 
.A(n_312),
.B(n_201),
.Y(n_415)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_327),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_311),
.A2(n_274),
.B1(n_257),
.B2(n_206),
.Y(n_417)
);

AND2x6_ASAP7_75t_L g418 ( 
.A(n_365),
.B(n_249),
.Y(n_418)
);

BUFx10_ASAP7_75t_L g419 ( 
.A(n_352),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_315),
.B(n_254),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_364),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_309),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_310),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_378),
.Y(n_424)
);

OAI22xp33_ASAP7_75t_L g425 ( 
.A1(n_306),
.A2(n_253),
.B1(n_205),
.B2(n_247),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_375),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_378),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_310),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_321),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_311),
.B(n_194),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_309),
.Y(n_431)
);

NOR2x1p5_ASAP7_75t_L g432 ( 
.A(n_366),
.B(n_202),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_378),
.Y(n_433)
);

INVx5_ASAP7_75t_L g434 ( 
.A(n_327),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_345),
.B(n_273),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_375),
.B(n_304),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_351),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_319),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_375),
.B(n_275),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_365),
.B(n_337),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_375),
.B(n_276),
.Y(n_441)
);

AND2x6_ASAP7_75t_L g442 ( 
.A(n_358),
.B(n_282),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_319),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_351),
.Y(n_444)
);

INVxp33_ASAP7_75t_L g445 ( 
.A(n_305),
.Y(n_445)
);

AND2x2_ASAP7_75t_SL g446 ( 
.A(n_348),
.B(n_287),
.Y(n_446)
);

AND3x1_ASAP7_75t_L g447 ( 
.A(n_307),
.B(n_316),
.C(n_377),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_328),
.Y(n_448)
);

OAI22xp33_ASAP7_75t_L g449 ( 
.A1(n_366),
.A2(n_259),
.B1(n_262),
.B2(n_266),
.Y(n_449)
);

NOR2x1_ASAP7_75t_L g450 ( 
.A(n_350),
.B(n_359),
.Y(n_450)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_327),
.Y(n_451)
);

NAND2xp33_ASAP7_75t_L g452 ( 
.A(n_327),
.B(n_303),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_344),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_356),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_356),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_358),
.B(n_283),
.Y(n_456)
);

AO22x2_ASAP7_75t_L g457 ( 
.A1(n_376),
.A2(n_326),
.B1(n_367),
.B2(n_362),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_SL g458 ( 
.A1(n_376),
.A2(n_257),
.B1(n_298),
.B2(n_295),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_373),
.Y(n_459)
);

INVx5_ASAP7_75t_L g460 ( 
.A(n_354),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_330),
.Y(n_461)
);

INVxp33_ASAP7_75t_L g462 ( 
.A(n_333),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_362),
.B(n_290),
.Y(n_463)
);

AND2x6_ASAP7_75t_L g464 ( 
.A(n_367),
.B(n_296),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_322),
.B(n_297),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_322),
.B(n_196),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_323),
.B(n_196),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_466),
.B(n_341),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_405),
.B(n_321),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_418),
.A2(n_323),
.B1(n_298),
.B2(n_295),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_447),
.A2(n_418),
.B1(n_425),
.B2(n_420),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_424),
.B(n_285),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_416),
.B(n_286),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_427),
.B(n_289),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_433),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_430),
.B(n_183),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_437),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_444),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_418),
.A2(n_212),
.B1(n_251),
.B2(n_308),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_440),
.B(n_203),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_451),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_462),
.B(n_270),
.Y(n_482)
);

AO22x1_ASAP7_75t_L g483 ( 
.A1(n_404),
.A2(n_279),
.B1(n_240),
.B2(n_241),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_388),
.B(n_244),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_402),
.B(n_317),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_411),
.B(n_317),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_410),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_445),
.B(n_250),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_451),
.B(n_434),
.Y(n_489)
);

AOI22xp33_ASAP7_75t_L g490 ( 
.A1(n_418),
.A2(n_317),
.B1(n_349),
.B2(n_346),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_L g491 ( 
.A1(n_382),
.A2(n_353),
.B1(n_349),
.B2(n_360),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_401),
.B(n_207),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g493 ( 
.A(n_405),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_383),
.Y(n_494)
);

INVx8_ASAP7_75t_L g495 ( 
.A(n_401),
.Y(n_495)
);

AND2x6_ASAP7_75t_L g496 ( 
.A(n_421),
.B(n_360),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_406),
.B(n_278),
.Y(n_497)
);

NOR3xp33_ASAP7_75t_SL g498 ( 
.A(n_449),
.B(n_291),
.C(n_294),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_393),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_395),
.Y(n_500)
);

BUFx12f_ASAP7_75t_L g501 ( 
.A(n_401),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_425),
.A2(n_300),
.B1(n_263),
.B2(n_371),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_420),
.B(n_407),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_396),
.Y(n_504)
);

INVx8_ASAP7_75t_L g505 ( 
.A(n_392),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_429),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_392),
.A2(n_371),
.B1(n_354),
.B2(n_369),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_406),
.B(n_371),
.Y(n_508)
);

NAND2x1p5_ASAP7_75t_L g509 ( 
.A(n_446),
.B(n_354),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_385),
.A2(n_354),
.B(n_369),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_412),
.B(n_309),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_390),
.Y(n_512)
);

NAND2x1_ASAP7_75t_L g513 ( 
.A(n_392),
.B(n_309),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_412),
.B(n_320),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_467),
.B(n_320),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_446),
.A2(n_370),
.B1(n_369),
.B2(n_368),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_400),
.B(n_18),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_461),
.Y(n_518)
);

NOR3xp33_ASAP7_75t_L g519 ( 
.A(n_449),
.B(n_458),
.C(n_391),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_415),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_413),
.B(n_57),
.Y(n_521)
);

NOR3xp33_ASAP7_75t_L g522 ( 
.A(n_458),
.B(n_18),
.C(n_19),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_392),
.A2(n_370),
.B1(n_369),
.B2(n_368),
.Y(n_523)
);

BUFx6f_ASAP7_75t_SL g524 ( 
.A(n_407),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_428),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_442),
.B(n_320),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_380),
.A2(n_370),
.B1(n_369),
.B2(n_368),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_419),
.Y(n_528)
);

AND2x6_ASAP7_75t_L g529 ( 
.A(n_381),
.B(n_325),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_419),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_423),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_380),
.B(n_325),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_413),
.B(n_58),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_384),
.B(n_325),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_384),
.B(n_389),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_459),
.B(n_325),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_389),
.B(n_331),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_407),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_467),
.B(n_450),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_432),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_392),
.A2(n_343),
.B1(n_340),
.B2(n_334),
.Y(n_541)
);

OR2x2_ASAP7_75t_L g542 ( 
.A(n_379),
.B(n_20),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_442),
.B(n_343),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_485),
.A2(n_452),
.B(n_386),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_476),
.B(n_398),
.Y(n_545)
);

O2A1O1Ixp33_ASAP7_75t_SL g546 ( 
.A1(n_513),
.A2(n_386),
.B(n_379),
.C(n_387),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_493),
.A2(n_403),
.B1(n_409),
.B2(n_457),
.Y(n_547)
);

O2A1O1Ixp5_ASAP7_75t_L g548 ( 
.A1(n_508),
.A2(n_439),
.B(n_441),
.C(n_463),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_476),
.B(n_399),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_539),
.B(n_403),
.Y(n_550)
);

A2O1A1Ixp33_ASAP7_75t_L g551 ( 
.A1(n_502),
.A2(n_463),
.B(n_441),
.C(n_439),
.Y(n_551)
);

AOI33xp33_ASAP7_75t_L g552 ( 
.A1(n_520),
.A2(n_453),
.A3(n_455),
.B1(n_438),
.B2(n_448),
.B3(n_443),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_473),
.B(n_426),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_477),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_487),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_486),
.A2(n_436),
.B(n_435),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_478),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_486),
.A2(n_436),
.B(n_435),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_503),
.B(n_394),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_468),
.B(n_472),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_471),
.A2(n_394),
.B1(n_456),
.B2(n_457),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_489),
.A2(n_465),
.B(n_408),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_494),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_481),
.B(n_465),
.Y(n_564)
);

NAND2x1p5_ASAP7_75t_L g565 ( 
.A(n_530),
.B(n_454),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_470),
.A2(n_457),
.B1(n_403),
.B2(n_409),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_468),
.B(n_403),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_535),
.A2(n_403),
.B1(n_409),
.B2(n_442),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_475),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_472),
.B(n_409),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_503),
.B(n_442),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_SL g572 ( 
.A1(n_495),
.A2(n_397),
.B1(n_442),
.B2(n_464),
.Y(n_572)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_469),
.Y(n_573)
);

OR2x6_ASAP7_75t_L g574 ( 
.A(n_495),
.B(n_501),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_509),
.A2(n_397),
.B1(n_460),
.B2(n_340),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_474),
.B(n_542),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_499),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_474),
.B(n_464),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_488),
.B(n_464),
.Y(n_579)
);

O2A1O1Ixp5_ASAP7_75t_L g580 ( 
.A1(n_534),
.A2(n_464),
.B(n_431),
.C(n_422),
.Y(n_580)
);

O2A1O1Ixp33_ASAP7_75t_L g581 ( 
.A1(n_532),
.A2(n_20),
.B(n_22),
.C(n_23),
.Y(n_581)
);

OAI22x1_ASAP7_75t_L g582 ( 
.A1(n_479),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_517),
.B(n_24),
.Y(n_583)
);

O2A1O1Ixp33_ASAP7_75t_L g584 ( 
.A1(n_537),
.A2(n_25),
.B(n_26),
.C(n_29),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_538),
.B(n_482),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_480),
.B(n_26),
.Y(n_586)
);

NAND2xp33_ASAP7_75t_L g587 ( 
.A(n_505),
.B(n_460),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_528),
.B(n_29),
.Y(n_588)
);

INVxp67_ASAP7_75t_L g589 ( 
.A(n_524),
.Y(n_589)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_511),
.A2(n_514),
.B(n_490),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_L g591 ( 
.A1(n_507),
.A2(n_460),
.B(n_431),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_495),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_500),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_506),
.Y(n_594)
);

NAND3xp33_ASAP7_75t_SL g595 ( 
.A(n_522),
.B(n_519),
.C(n_498),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_515),
.A2(n_422),
.B(n_414),
.Y(n_596)
);

NAND3xp33_ASAP7_75t_SL g597 ( 
.A(n_516),
.B(n_31),
.C(n_33),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_505),
.A2(n_334),
.B1(n_332),
.B2(n_331),
.Y(n_598)
);

O2A1O1Ixp33_ASAP7_75t_SL g599 ( 
.A1(n_543),
.A2(n_108),
.B(n_181),
.C(n_169),
.Y(n_599)
);

NAND2xp33_ASAP7_75t_L g600 ( 
.A(n_481),
.B(n_331),
.Y(n_600)
);

NAND2xp33_ASAP7_75t_SL g601 ( 
.A(n_524),
.B(n_331),
.Y(n_601)
);

A2O1A1Ixp33_ASAP7_75t_L g602 ( 
.A1(n_521),
.A2(n_334),
.B(n_332),
.C(n_331),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_481),
.B(n_332),
.Y(n_603)
);

O2A1O1Ixp33_ASAP7_75t_L g604 ( 
.A1(n_527),
.A2(n_34),
.B(n_35),
.C(n_38),
.Y(n_604)
);

AOI21x1_ASAP7_75t_L g605 ( 
.A1(n_543),
.A2(n_334),
.B(n_332),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_483),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_492),
.B(n_35),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_526),
.B(n_39),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_L g609 ( 
.A1(n_504),
.A2(n_39),
.B1(n_40),
.B2(n_45),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_531),
.B(n_40),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_492),
.B(n_45),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_518),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_484),
.B(n_63),
.Y(n_613)
);

A2O1A1Ixp33_ASAP7_75t_L g614 ( 
.A1(n_533),
.A2(n_66),
.B(n_67),
.C(n_72),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_497),
.B(n_73),
.Y(n_615)
);

AO21x1_ASAP7_75t_L g616 ( 
.A1(n_527),
.A2(n_82),
.B(n_83),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_526),
.B(n_84),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_540),
.B(n_98),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_525),
.A2(n_99),
.B1(n_101),
.B2(n_102),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_554),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_563),
.Y(n_621)
);

OAI21x1_ASAP7_75t_L g622 ( 
.A1(n_580),
.A2(n_510),
.B(n_536),
.Y(n_622)
);

AO21x2_ASAP7_75t_L g623 ( 
.A1(n_591),
.A2(n_510),
.B(n_523),
.Y(n_623)
);

INVx5_ASAP7_75t_L g624 ( 
.A(n_592),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_592),
.B(n_491),
.Y(n_625)
);

INVxp67_ASAP7_75t_L g626 ( 
.A(n_555),
.Y(n_626)
);

OAI21x1_ASAP7_75t_L g627 ( 
.A1(n_605),
.A2(n_541),
.B(n_512),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_L g628 ( 
.A1(n_548),
.A2(n_544),
.B(n_590),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_557),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_569),
.Y(n_630)
);

AOI21xp33_ASAP7_75t_L g631 ( 
.A1(n_585),
.A2(n_496),
.B(n_105),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_574),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_556),
.A2(n_496),
.B(n_529),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_577),
.Y(n_634)
);

BUFx12f_ASAP7_75t_L g635 ( 
.A(n_574),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_L g636 ( 
.A1(n_548),
.A2(n_529),
.B(n_107),
.Y(n_636)
);

AO31x2_ASAP7_75t_L g637 ( 
.A1(n_561),
.A2(n_602),
.A3(n_551),
.B(n_614),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_593),
.Y(n_638)
);

CKINVDCx11_ASAP7_75t_R g639 ( 
.A(n_574),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_558),
.A2(n_104),
.B(n_109),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_570),
.A2(n_110),
.B(n_111),
.Y(n_641)
);

BUFx4_ASAP7_75t_SL g642 ( 
.A(n_594),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_567),
.A2(n_112),
.B(n_113),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_568),
.A2(n_114),
.B(n_115),
.Y(n_644)
);

AOI221xp5_ASAP7_75t_L g645 ( 
.A1(n_573),
.A2(n_124),
.B1(n_125),
.B2(n_129),
.C(n_130),
.Y(n_645)
);

NOR2xp67_ASAP7_75t_SL g646 ( 
.A(n_606),
.B(n_131),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_595),
.A2(n_133),
.B1(n_138),
.B2(n_140),
.Y(n_647)
);

OR2x2_ASAP7_75t_L g648 ( 
.A(n_575),
.B(n_145),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_578),
.A2(n_159),
.B(n_162),
.Y(n_649)
);

INVx3_ASAP7_75t_SL g650 ( 
.A(n_571),
.Y(n_650)
);

O2A1O1Ixp5_ASAP7_75t_L g651 ( 
.A1(n_553),
.A2(n_579),
.B(n_615),
.C(n_613),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_546),
.A2(n_550),
.B(n_562),
.Y(n_652)
);

OR2x6_ASAP7_75t_L g653 ( 
.A(n_565),
.B(n_589),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_564),
.A2(n_545),
.B(n_549),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_583),
.B(n_547),
.Y(n_655)
);

NOR2x1_ASAP7_75t_R g656 ( 
.A(n_572),
.B(n_588),
.Y(n_656)
);

A2O1A1Ixp33_ASAP7_75t_L g657 ( 
.A1(n_552),
.A2(n_604),
.B(n_581),
.C(n_584),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_582),
.Y(n_658)
);

O2A1O1Ixp33_ASAP7_75t_L g659 ( 
.A1(n_604),
.A2(n_610),
.B(n_609),
.C(n_584),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_565),
.B(n_607),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_612),
.Y(n_661)
);

AO32x2_ASAP7_75t_L g662 ( 
.A1(n_598),
.A2(n_619),
.A3(n_597),
.B1(n_581),
.B2(n_599),
.Y(n_662)
);

OAI21x1_ASAP7_75t_L g663 ( 
.A1(n_603),
.A2(n_617),
.B(n_608),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_597),
.Y(n_664)
);

NAND3xp33_ASAP7_75t_SL g665 ( 
.A(n_611),
.B(n_618),
.C(n_601),
.Y(n_665)
);

AO31x2_ASAP7_75t_L g666 ( 
.A1(n_600),
.A2(n_616),
.A3(n_508),
.B(n_561),
.Y(n_666)
);

OAI22x1_ASAP7_75t_L g667 ( 
.A1(n_587),
.A2(n_417),
.B1(n_366),
.B2(n_471),
.Y(n_667)
);

NAND2x1p5_ASAP7_75t_L g668 ( 
.A(n_592),
.B(n_487),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_SL g669 ( 
.A1(n_575),
.A2(n_376),
.B1(n_366),
.B2(n_487),
.Y(n_669)
);

BUFx12f_ASAP7_75t_L g670 ( 
.A(n_574),
.Y(n_670)
);

INVx3_ASAP7_75t_SL g671 ( 
.A(n_574),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_573),
.B(n_487),
.Y(n_672)
);

OAI21x1_ASAP7_75t_L g673 ( 
.A1(n_580),
.A2(n_605),
.B(n_596),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_559),
.B(n_560),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_559),
.B(n_560),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_569),
.Y(n_676)
);

OAI22x1_ASAP7_75t_L g677 ( 
.A1(n_547),
.A2(n_417),
.B1(n_366),
.B2(n_471),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_573),
.A2(n_487),
.B1(n_366),
.B2(n_417),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_559),
.B(n_560),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_554),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_559),
.B(n_560),
.Y(n_681)
);

AO32x2_ASAP7_75t_L g682 ( 
.A1(n_561),
.A2(n_566),
.A3(n_527),
.B1(n_609),
.B2(n_575),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_592),
.B(n_571),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_573),
.B(n_487),
.Y(n_684)
);

AO31x2_ASAP7_75t_L g685 ( 
.A1(n_616),
.A2(n_508),
.A3(n_561),
.B(n_602),
.Y(n_685)
);

OAI22xp5_ASAP7_75t_L g686 ( 
.A1(n_576),
.A2(n_471),
.B1(n_470),
.B2(n_566),
.Y(n_686)
);

A2O1A1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_560),
.A2(n_586),
.B(n_548),
.C(n_576),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_573),
.B(n_487),
.Y(n_688)
);

OAI21x1_ASAP7_75t_L g689 ( 
.A1(n_580),
.A2(n_605),
.B(n_596),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_559),
.B(n_560),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_573),
.B(n_487),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_559),
.B(n_560),
.Y(n_692)
);

OAI21x1_ASAP7_75t_L g693 ( 
.A1(n_580),
.A2(n_605),
.B(n_596),
.Y(n_693)
);

OAI22xp5_ASAP7_75t_L g694 ( 
.A1(n_576),
.A2(n_471),
.B1(n_470),
.B2(n_566),
.Y(n_694)
);

A2O1A1Ixp33_ASAP7_75t_L g695 ( 
.A1(n_560),
.A2(n_586),
.B(n_548),
.C(n_576),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_554),
.Y(n_696)
);

AO31x2_ASAP7_75t_L g697 ( 
.A1(n_616),
.A2(n_508),
.A3(n_561),
.B(n_602),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_554),
.Y(n_698)
);

AO31x2_ASAP7_75t_L g699 ( 
.A1(n_616),
.A2(n_508),
.A3(n_561),
.B(n_602),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_574),
.Y(n_700)
);

OAI21xp5_ASAP7_75t_L g701 ( 
.A1(n_548),
.A2(n_544),
.B(n_590),
.Y(n_701)
);

OAI21xp5_ASAP7_75t_L g702 ( 
.A1(n_548),
.A2(n_544),
.B(n_590),
.Y(n_702)
);

INVx8_ASAP7_75t_L g703 ( 
.A(n_574),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_573),
.B(n_487),
.Y(n_704)
);

OAI22x1_ASAP7_75t_L g705 ( 
.A1(n_547),
.A2(n_417),
.B1(n_366),
.B2(n_471),
.Y(n_705)
);

OR2x6_ASAP7_75t_L g706 ( 
.A(n_703),
.B(n_635),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_674),
.B(n_675),
.Y(n_707)
);

INVxp67_ASAP7_75t_L g708 ( 
.A(n_684),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_676),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_686),
.A2(n_694),
.B1(n_655),
.B2(n_648),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_672),
.B(n_688),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_620),
.Y(n_712)
);

NOR2x1_ASAP7_75t_SL g713 ( 
.A(n_624),
.B(n_653),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_679),
.B(n_681),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_680),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_624),
.B(n_683),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_624),
.Y(n_717)
);

A2O1A1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_687),
.A2(n_695),
.B(n_659),
.C(n_654),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_683),
.Y(n_719)
);

AND2x4_ASAP7_75t_SL g720 ( 
.A(n_621),
.B(n_653),
.Y(n_720)
);

INVxp67_ASAP7_75t_L g721 ( 
.A(n_691),
.Y(n_721)
);

BUFx12f_ASAP7_75t_L g722 ( 
.A(n_639),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_703),
.Y(n_723)
);

AO21x2_ASAP7_75t_L g724 ( 
.A1(n_636),
.A2(n_657),
.B(n_652),
.Y(n_724)
);

OA21x2_ASAP7_75t_L g725 ( 
.A1(n_673),
.A2(n_689),
.B(n_693),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_629),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_690),
.B(n_692),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_669),
.A2(n_705),
.B1(n_677),
.B2(n_667),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_630),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_634),
.B(n_638),
.Y(n_730)
);

OAI21xp5_ASAP7_75t_L g731 ( 
.A1(n_633),
.A2(n_644),
.B(n_651),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_671),
.Y(n_732)
);

HB1xp67_ASAP7_75t_L g733 ( 
.A(n_642),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_678),
.B(n_704),
.Y(n_734)
);

NAND2x1p5_ASAP7_75t_L g735 ( 
.A(n_632),
.B(n_700),
.Y(n_735)
);

OAI22xp33_ASAP7_75t_L g736 ( 
.A1(n_658),
.A2(n_670),
.B1(n_668),
.B2(n_626),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_650),
.Y(n_737)
);

OAI21x1_ASAP7_75t_L g738 ( 
.A1(n_622),
.A2(n_663),
.B(n_627),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_696),
.Y(n_739)
);

AO31x2_ASAP7_75t_L g740 ( 
.A1(n_640),
.A2(n_649),
.A3(n_641),
.B(n_643),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_698),
.Y(n_741)
);

AOI221xp5_ASAP7_75t_L g742 ( 
.A1(n_638),
.A2(n_661),
.B1(n_660),
.B2(n_664),
.C(n_665),
.Y(n_742)
);

BUFx2_ASAP7_75t_L g743 ( 
.A(n_656),
.Y(n_743)
);

HB1xp67_ASAP7_75t_L g744 ( 
.A(n_625),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_631),
.A2(n_623),
.B(n_664),
.Y(n_745)
);

AOI21xp33_ASAP7_75t_L g746 ( 
.A1(n_646),
.A2(n_647),
.B(n_645),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_682),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_682),
.B(n_637),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_682),
.B(n_662),
.Y(n_749)
);

HB1xp67_ASAP7_75t_L g750 ( 
.A(n_637),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_662),
.B(n_666),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_685),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_685),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_662),
.B(n_666),
.Y(n_754)
);

CKINVDCx11_ASAP7_75t_R g755 ( 
.A(n_685),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_699),
.B(n_697),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_697),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_699),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_684),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_621),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_686),
.A2(n_694),
.B1(n_655),
.B2(n_648),
.Y(n_761)
);

A2O1A1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_687),
.A2(n_695),
.B(n_659),
.C(n_654),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_624),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_674),
.B(n_675),
.Y(n_764)
);

AND2x4_ASAP7_75t_SL g765 ( 
.A(n_621),
.B(n_592),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_620),
.Y(n_766)
);

XNOR2xp5_ASAP7_75t_L g767 ( 
.A(n_621),
.B(n_397),
.Y(n_767)
);

CKINVDCx11_ASAP7_75t_R g768 ( 
.A(n_639),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_678),
.B(n_366),
.Y(n_769)
);

OA21x2_ASAP7_75t_L g770 ( 
.A1(n_628),
.A2(n_702),
.B(n_701),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_624),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_674),
.B(n_675),
.Y(n_772)
);

INVx1_ASAP7_75t_SL g773 ( 
.A(n_672),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_620),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_674),
.B(n_675),
.Y(n_775)
);

HB1xp67_ASAP7_75t_L g776 ( 
.A(n_711),
.Y(n_776)
);

NAND2x1p5_ASAP7_75t_L g777 ( 
.A(n_717),
.B(n_771),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_717),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_730),
.Y(n_779)
);

INVxp33_ASAP7_75t_L g780 ( 
.A(n_733),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_709),
.Y(n_781)
);

OR2x6_ASAP7_75t_L g782 ( 
.A(n_710),
.B(n_761),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_717),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_716),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_727),
.B(n_707),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_716),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_773),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_773),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_771),
.Y(n_789)
);

BUFx3_ASAP7_75t_L g790 ( 
.A(n_763),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_765),
.Y(n_791)
);

INVxp67_ASAP7_75t_L g792 ( 
.A(n_760),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_R g793 ( 
.A(n_706),
.B(n_743),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_726),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_720),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_729),
.Y(n_796)
);

AO31x2_ASAP7_75t_L g797 ( 
.A1(n_751),
.A2(n_754),
.A3(n_718),
.B(n_762),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_712),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_706),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_706),
.Y(n_800)
);

BUFx2_ASAP7_75t_L g801 ( 
.A(n_770),
.Y(n_801)
);

INVxp67_ASAP7_75t_L g802 ( 
.A(n_714),
.Y(n_802)
);

OAI21x1_ASAP7_75t_L g803 ( 
.A1(n_738),
.A2(n_731),
.B(n_745),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_725),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_739),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_741),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_714),
.B(n_775),
.Y(n_807)
);

HB1xp67_ASAP7_75t_L g808 ( 
.A(n_715),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_750),
.Y(n_809)
);

CKINVDCx20_ASAP7_75t_R g810 ( 
.A(n_768),
.Y(n_810)
);

AO21x2_ASAP7_75t_L g811 ( 
.A1(n_756),
.A2(n_731),
.B(n_724),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_764),
.B(n_775),
.Y(n_812)
);

INVxp67_ASAP7_75t_L g813 ( 
.A(n_764),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_766),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_772),
.B(n_774),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_772),
.B(n_734),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_747),
.B(n_758),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_769),
.B(n_708),
.Y(n_818)
);

INVx1_ASAP7_75t_SL g819 ( 
.A(n_737),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_752),
.Y(n_820)
);

AO21x2_ASAP7_75t_L g821 ( 
.A1(n_724),
.A2(n_757),
.B(n_749),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_744),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_748),
.B(n_753),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_713),
.Y(n_824)
);

OA21x2_ASAP7_75t_L g825 ( 
.A1(n_742),
.A2(n_710),
.B(n_761),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_721),
.B(n_759),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_820),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_824),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_782),
.B(n_823),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_782),
.B(n_755),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_787),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_782),
.B(n_728),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_793),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_807),
.B(n_767),
.Y(n_834)
);

HB1xp67_ASAP7_75t_L g835 ( 
.A(n_788),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_782),
.B(n_719),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_823),
.B(n_737),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_812),
.B(n_719),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_812),
.B(n_736),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_817),
.Y(n_840)
);

INVxp67_ASAP7_75t_SL g841 ( 
.A(n_798),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_776),
.Y(n_842)
);

AOI21xp33_ASAP7_75t_L g843 ( 
.A1(n_816),
.A2(n_746),
.B(n_723),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_815),
.B(n_797),
.Y(n_844)
);

HB1xp67_ASAP7_75t_L g845 ( 
.A(n_808),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_783),
.Y(n_846)
);

NOR2x1_ASAP7_75t_R g847 ( 
.A(n_791),
.B(n_722),
.Y(n_847)
);

INVxp67_ASAP7_75t_SL g848 ( 
.A(n_814),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_815),
.B(n_735),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_SL g850 ( 
.A(n_810),
.B(n_732),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_797),
.B(n_740),
.Y(n_851)
);

OR2x2_ASAP7_75t_L g852 ( 
.A(n_785),
.B(n_740),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_802),
.B(n_740),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_790),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_813),
.B(n_779),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_797),
.B(n_781),
.Y(n_856)
);

OR2x2_ASAP7_75t_L g857 ( 
.A(n_822),
.B(n_809),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_804),
.Y(n_858)
);

INVxp33_ASAP7_75t_L g859 ( 
.A(n_795),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_790),
.Y(n_860)
);

BUFx2_ASAP7_75t_SL g861 ( 
.A(n_790),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_844),
.B(n_856),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_844),
.B(n_801),
.Y(n_863)
);

NAND2x1p5_ASAP7_75t_L g864 ( 
.A(n_828),
.B(n_846),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_856),
.B(n_801),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_827),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_858),
.Y(n_867)
);

OR2x6_ASAP7_75t_L g868 ( 
.A(n_861),
.B(n_803),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_828),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_829),
.B(n_821),
.Y(n_870)
);

AND2x6_ASAP7_75t_SL g871 ( 
.A(n_847),
.B(n_818),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_829),
.B(n_821),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_SL g873 ( 
.A(n_861),
.B(n_799),
.Y(n_873)
);

OR2x2_ASAP7_75t_L g874 ( 
.A(n_857),
.B(n_852),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_839),
.B(n_800),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_857),
.B(n_811),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_845),
.Y(n_877)
);

NOR2x1_ASAP7_75t_L g878 ( 
.A(n_869),
.B(n_837),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_866),
.Y(n_879)
);

OR2x2_ASAP7_75t_L g880 ( 
.A(n_874),
.B(n_852),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_862),
.B(n_870),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_862),
.B(n_851),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_870),
.B(n_872),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_872),
.B(n_851),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_874),
.B(n_853),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_867),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_877),
.B(n_842),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_863),
.B(n_851),
.Y(n_888)
);

OR2x2_ASAP7_75t_L g889 ( 
.A(n_876),
.B(n_840),
.Y(n_889)
);

OR2x2_ASAP7_75t_L g890 ( 
.A(n_876),
.B(n_831),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_871),
.B(n_780),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_877),
.B(n_841),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_868),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_880),
.B(n_865),
.Y(n_894)
);

AOI221xp5_ASAP7_75t_L g895 ( 
.A1(n_887),
.A2(n_843),
.B1(n_832),
.B2(n_875),
.C(n_835),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_891),
.B(n_871),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_890),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_892),
.B(n_819),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_880),
.B(n_865),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_890),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_879),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_881),
.B(n_832),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_886),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_885),
.B(n_837),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_878),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_881),
.B(n_882),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_878),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_906),
.B(n_883),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_897),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_896),
.A2(n_875),
.B1(n_884),
.B2(n_882),
.Y(n_910)
);

INVx1_ASAP7_75t_SL g911 ( 
.A(n_894),
.Y(n_911)
);

BUFx2_ASAP7_75t_SL g912 ( 
.A(n_905),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_896),
.A2(n_884),
.B1(n_833),
.B2(n_888),
.Y(n_913)
);

XOR2x2_ASAP7_75t_L g914 ( 
.A(n_904),
.B(n_850),
.Y(n_914)
);

NOR3xp33_ASAP7_75t_L g915 ( 
.A(n_895),
.B(n_847),
.C(n_826),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_900),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_904),
.B(n_883),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_903),
.Y(n_918)
);

OAI21xp33_ASAP7_75t_SL g919 ( 
.A1(n_907),
.A2(n_893),
.B(n_888),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_898),
.A2(n_830),
.B1(n_836),
.B2(n_838),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_919),
.A2(n_873),
.B(n_833),
.Y(n_921)
);

AOI21xp33_ASAP7_75t_SL g922 ( 
.A1(n_915),
.A2(n_864),
.B(n_898),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_912),
.B(n_792),
.Y(n_923)
);

AOI211xp5_ASAP7_75t_L g924 ( 
.A1(n_915),
.A2(n_859),
.B(n_830),
.C(n_893),
.Y(n_924)
);

O2A1O1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_909),
.A2(n_834),
.B(n_800),
.C(n_799),
.Y(n_925)
);

OAI31xp33_ASAP7_75t_L g926 ( 
.A1(n_911),
.A2(n_869),
.A3(n_893),
.B(n_864),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_918),
.Y(n_927)
);

AOI221xp5_ASAP7_75t_L g928 ( 
.A1(n_922),
.A2(n_916),
.B1(n_920),
.B2(n_917),
.C(n_910),
.Y(n_928)
);

NAND4xp25_ASAP7_75t_L g929 ( 
.A(n_924),
.B(n_913),
.C(n_920),
.D(n_873),
.Y(n_929)
);

AOI221xp5_ASAP7_75t_L g930 ( 
.A1(n_925),
.A2(n_902),
.B1(n_908),
.B2(n_901),
.C(n_918),
.Y(n_930)
);

NAND4xp75_ASAP7_75t_L g931 ( 
.A(n_928),
.B(n_921),
.C(n_926),
.D(n_923),
.Y(n_931)
);

AOI221x1_ASAP7_75t_L g932 ( 
.A1(n_929),
.A2(n_927),
.B1(n_914),
.B2(n_789),
.C(n_778),
.Y(n_932)
);

NOR4xp25_ASAP7_75t_L g933 ( 
.A(n_931),
.B(n_930),
.C(n_791),
.D(n_806),
.Y(n_933)
);

NAND3xp33_ASAP7_75t_L g934 ( 
.A(n_932),
.B(n_860),
.C(n_854),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_934),
.Y(n_935)
);

NAND4xp75_ASAP7_75t_L g936 ( 
.A(n_933),
.B(n_825),
.C(n_786),
.D(n_784),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_935),
.B(n_893),
.Y(n_937)
);

NOR2x1_ASAP7_75t_L g938 ( 
.A(n_936),
.B(n_869),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_937),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_938),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_937),
.Y(n_941)
);

OA21x2_ASAP7_75t_L g942 ( 
.A1(n_939),
.A2(n_848),
.B(n_855),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_SL g943 ( 
.A1(n_940),
.A2(n_864),
.B1(n_777),
.B2(n_784),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_940),
.A2(n_899),
.B1(n_885),
.B2(n_889),
.Y(n_944)
);

AOI22x1_ASAP7_75t_L g945 ( 
.A1(n_941),
.A2(n_777),
.B1(n_778),
.B2(n_789),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_939),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_946),
.A2(n_786),
.B1(n_849),
.B2(n_789),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_942),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_945),
.A2(n_777),
.B(n_796),
.Y(n_949)
);

INVxp67_ASAP7_75t_L g950 ( 
.A(n_943),
.Y(n_950)
);

INVxp67_ASAP7_75t_L g951 ( 
.A(n_944),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_946),
.B(n_794),
.Y(n_952)
);

NAND3xp33_ASAP7_75t_L g953 ( 
.A(n_950),
.B(n_951),
.C(n_948),
.Y(n_953)
);

NOR2x1_ASAP7_75t_R g954 ( 
.A(n_952),
.B(n_846),
.Y(n_954)
);

AOI21xp33_ASAP7_75t_L g955 ( 
.A1(n_949),
.A2(n_806),
.B(n_805),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_954),
.Y(n_956)
);

AOI22xp33_ASAP7_75t_L g957 ( 
.A1(n_956),
.A2(n_953),
.B1(n_955),
.B2(n_947),
.Y(n_957)
);


endmodule