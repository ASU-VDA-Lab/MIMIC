module fake_jpeg_19136_n_174 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_174);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx6f_ASAP7_75t_SL g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_SL g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g30 ( 
.A(n_15),
.B(n_0),
.CON(n_30),
.SN(n_30)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_18),
.B(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_34),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_35),
.A2(n_22),
.B1(n_20),
.B2(n_24),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_40),
.A2(n_50),
.B1(n_19),
.B2(n_25),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_48),
.B1(n_26),
.B2(n_15),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_21),
.B1(n_24),
.B2(n_14),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_14),
.B1(n_18),
.B2(n_28),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_45),
.B(n_31),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_52),
.B(n_54),
.Y(n_80)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_57),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_32),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_38),
.B1(n_28),
.B2(n_16),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_55),
.A2(n_58),
.B1(n_60),
.B2(n_43),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_59),
.Y(n_90)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_37),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_16),
.B1(n_19),
.B2(n_27),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_63),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_37),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_62),
.B(n_66),
.Y(n_92)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_72),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_33),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_27),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_67),
.B(n_68),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_27),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_23),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_73),
.B(n_76),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_23),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_23),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_29),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_2),
.Y(n_94)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_82),
.A2(n_89),
.B1(n_55),
.B2(n_70),
.Y(n_110)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_65),
.A2(n_43),
.B1(n_29),
.B2(n_39),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_84),
.A2(n_88),
.B1(n_6),
.B2(n_7),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_2),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_70),
.B(n_73),
.Y(n_108)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_65),
.A2(n_39),
.B1(n_25),
.B2(n_4),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_62),
.A2(n_25),
.B1(n_3),
.B2(n_4),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_9),
.Y(n_98)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_98),
.B(n_100),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_53),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_61),
.Y(n_101)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_51),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_104),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_51),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_58),
.Y(n_105)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

AND2x4_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_73),
.Y(n_107)
);

AND2x4_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_81),
.Y(n_120)
);

NOR3xp33_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_89),
.C(n_81),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_111),
.B1(n_116),
.B2(n_87),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_82),
.A2(n_97),
.B1(n_92),
.B2(n_83),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_77),
.A2(n_75),
.B(n_5),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_112),
.A2(n_114),
.B(n_7),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_78),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_79),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_77),
.A2(n_4),
.B(n_5),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_6),
.Y(n_115)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_95),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_107),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_80),
.C(n_78),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_130),
.C(n_114),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_119),
.A2(n_120),
.B(n_126),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_110),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_129),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_112),
.A2(n_107),
.B(n_111),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_128),
.A2(n_115),
.B(n_108),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_103),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_79),
.C(n_8),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_137),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_142),
.B(n_143),
.Y(n_147)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_124),
.B1(n_121),
.B2(n_105),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_106),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_139),
.B(n_140),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_107),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_117),
.B(n_106),
.Y(n_141)
);

OA21x2_ASAP7_75t_SL g145 ( 
.A1(n_141),
.A2(n_120),
.B(n_127),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_99),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_107),
.B(n_109),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_145),
.B(n_133),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_120),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_148),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_128),
.B(n_122),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_131),
.Y(n_155)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_150),
.A2(n_136),
.B(n_143),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_157),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_158),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_152),
.A2(n_140),
.B(n_123),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_113),
.B(n_109),
.Y(n_158)
);

OAI22x1_ASAP7_75t_L g161 ( 
.A1(n_156),
.A2(n_147),
.B1(n_151),
.B2(n_146),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_161),
.A2(n_144),
.B1(n_103),
.B2(n_11),
.Y(n_167)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_165),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_144),
.C(n_132),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_160),
.B(n_131),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_167),
.Y(n_171)
);

AOI31xp33_ASAP7_75t_L g169 ( 
.A1(n_163),
.A2(n_8),
.A3(n_11),
.B(n_79),
.Y(n_169)
);

NAND2xp33_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_161),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_170),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_162),
.B1(n_167),
.B2(n_168),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_171),
.Y(n_174)
);


endmodule