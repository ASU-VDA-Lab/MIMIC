module fake_jpeg_20387_n_274 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_274);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g26 ( 
.A(n_17),
.Y(n_26)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_25),
.Y(n_34)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

HAxp5_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_28),
.CON(n_42),
.SN(n_42)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_30),
.A2(n_23),
.B1(n_14),
.B2(n_15),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_26),
.B1(n_29),
.B2(n_25),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_32),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_24),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_55),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_30),
.B1(n_26),
.B2(n_23),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_47),
.A2(n_38),
.B1(n_29),
.B2(n_25),
.Y(n_69)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_57),
.B1(n_38),
.B2(n_37),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_53),
.B(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_11),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_32),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_34),
.A2(n_26),
.B1(n_29),
.B2(n_31),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_23),
.B1(n_33),
.B2(n_26),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_60),
.A2(n_34),
.B1(n_38),
.B2(n_25),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_27),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_69),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_62),
.A2(n_44),
.B1(n_57),
.B2(n_60),
.Y(n_84)
);

AO21x2_ASAP7_75t_L g63 ( 
.A1(n_56),
.A2(n_38),
.B(n_39),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_77),
.B1(n_46),
.B2(n_40),
.Y(n_90)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_70),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_72),
.A2(n_73),
.B1(n_46),
.B2(n_41),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_31),
.B1(n_33),
.B2(n_27),
.Y(n_73)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_31),
.B1(n_41),
.B2(n_33),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_74),
.A2(n_55),
.B(n_35),
.Y(n_86)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_43),
.A2(n_41),
.B1(n_27),
.B2(n_16),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_56),
.B(n_44),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_67),
.B(n_62),
.Y(n_99)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_74),
.B1(n_73),
.B2(n_70),
.Y(n_105)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g120 ( 
.A1(n_86),
.A2(n_89),
.B1(n_90),
.B2(n_94),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_58),
.C(n_52),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_84),
.C(n_97),
.Y(n_104)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_88),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_72),
.B1(n_65),
.B2(n_63),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_98),
.B1(n_75),
.B2(n_66),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_65),
.A2(n_53),
.B1(n_40),
.B2(n_51),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_96),
.Y(n_107)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_93),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_63),
.A2(n_51),
.B1(n_40),
.B2(n_50),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_63),
.A2(n_40),
.B1(n_24),
.B2(n_32),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_63),
.A2(n_39),
.B1(n_24),
.B2(n_32),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_99),
.A2(n_81),
.B(n_12),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_82),
.B(n_64),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_101),
.B(n_116),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_102),
.B(n_114),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_119),
.C(n_96),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_121),
.B1(n_28),
.B2(n_39),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_112),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_74),
.B1(n_68),
.B2(n_71),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_109),
.A2(n_110),
.B1(n_59),
.B2(n_39),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_83),
.A2(n_68),
.B1(n_71),
.B2(n_80),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_64),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_87),
.B(n_78),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_113),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_85),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_78),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_59),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_35),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_90),
.B(n_20),
.Y(n_117)
);

XOR2x1_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_94),
.Y(n_126)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_80),
.C(n_24),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_103),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_124),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_123),
.B(n_120),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_103),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_106),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_130),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_126),
.A2(n_133),
.B1(n_147),
.B2(n_100),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_95),
.C(n_98),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_132),
.C(n_150),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_129),
.A2(n_144),
.B(n_148),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_106),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_81),
.C(n_66),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_134),
.A2(n_141),
.B1(n_149),
.B2(n_100),
.Y(n_158)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

BUFx4f_ASAP7_75t_SL g139 ( 
.A(n_118),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_145),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_108),
.A2(n_22),
.B1(n_12),
.B2(n_13),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_142),
.Y(n_160)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_143),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_10),
.B(n_9),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_28),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_15),
.B1(n_22),
.B2(n_12),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_111),
.A2(n_22),
.B1(n_15),
.B2(n_13),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_99),
.B(n_59),
.C(n_21),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_135),
.B(n_132),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_153),
.Y(n_183)
);

XNOR2x1_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_112),
.Y(n_153)
);

XNOR2x2_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_120),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_154),
.A2(n_131),
.B(n_6),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_105),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_159),
.C(n_169),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_157),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_158),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_119),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_162),
.A2(n_6),
.B1(n_9),
.B2(n_3),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_120),
.B1(n_13),
.B2(n_0),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_163),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_189)
);

INVxp33_ASAP7_75t_SL g166 ( 
.A(n_139),
.Y(n_166)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_6),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_133),
.A2(n_127),
.B1(n_146),
.B2(n_143),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_150),
.B1(n_145),
.B2(n_137),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_129),
.A2(n_120),
.B(n_21),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_173),
.B(n_149),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_18),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_175),
.C(n_172),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_18),
.C(n_11),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_177),
.B(n_181),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_142),
.Y(n_178)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_179),
.A2(n_189),
.B1(n_174),
.B2(n_156),
.Y(n_207)
);

AOI21x1_ASAP7_75t_L g180 ( 
.A1(n_154),
.A2(n_148),
.B(n_122),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_180),
.A2(n_188),
.B(n_153),
.Y(n_204)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_158),
.A2(n_136),
.B1(n_131),
.B2(n_141),
.Y(n_186)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_186),
.Y(n_200)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_190),
.A2(n_163),
.B1(n_168),
.B2(n_175),
.Y(n_202)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_176),
.Y(n_191)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_191),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_164),
.Y(n_192)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_193),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_0),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_194),
.Y(n_206)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_196),
.A2(n_155),
.B(n_7),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_197),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_152),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_203),
.Y(n_227)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_159),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_204),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_207),
.A2(n_188),
.B1(n_184),
.B2(n_191),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_169),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_182),
.C(n_197),
.Y(n_217)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_209),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_185),
.A2(n_155),
.B1(n_7),
.B2(n_3),
.Y(n_214)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_7),
.B1(n_9),
.B2(n_4),
.Y(n_215)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_218),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_192),
.Y(n_219)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_219),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_200),
.A2(n_184),
.B1(n_196),
.B2(n_195),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_220),
.A2(n_189),
.B1(n_211),
.B2(n_199),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_195),
.C(n_181),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_203),
.C(n_207),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_198),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_226),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_190),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_213),
.A2(n_178),
.B1(n_194),
.B2(n_180),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_222),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_231),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_204),
.B(n_206),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_212),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_235),
.Y(n_248)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_224),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_221),
.A2(n_206),
.B(n_202),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_237),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_4),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_239),
.B(n_240),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_4),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_223),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_242),
.B(n_250),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_233),
.B(n_224),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_249),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_238),
.A2(n_220),
.B(n_217),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_246),
.A2(n_247),
.B(n_236),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_238),
.A2(n_227),
.B(n_5),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_231),
.B(n_227),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_5),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_253),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_230),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_5),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_259),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_5),
.C(n_8),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_258),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_248),
.B(n_8),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_10),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_248),
.B(n_0),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_260),
.B(n_0),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_263),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_1),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_265),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_264),
.B(n_257),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_268),
.A2(n_262),
.B(n_260),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_261),
.C(n_254),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_269),
.A2(n_270),
.B(n_266),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_271),
.B(n_1),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_1),
.Y(n_273)
);

BUFx24_ASAP7_75t_SL g274 ( 
.A(n_273),
.Y(n_274)
);


endmodule