module fake_jpeg_30214_n_543 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_543);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_543;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_441;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_18;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_13),
.B(n_4),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_5),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_59),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_28),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_60),
.B(n_73),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_62),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_63),
.Y(n_125)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_65),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_67),
.Y(n_172)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_68),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_69),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_70),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_71),
.Y(n_170)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_28),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_74),
.Y(n_129)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_76),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_78),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_79),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_80),
.Y(n_156)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx4_ASAP7_75t_SL g84 ( 
.A(n_38),
.Y(n_84)
);

BUFx2_ASAP7_75t_R g139 ( 
.A(n_84),
.Y(n_139)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_88),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_92),
.Y(n_165)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_93),
.Y(n_166)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_94),
.Y(n_174)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_95),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_98),
.Y(n_136)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_101),
.Y(n_119)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_99),
.B(n_103),
.Y(n_146)
);

BUFx24_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_42),
.Y(n_118)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_27),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_105),
.Y(n_130)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_104),
.B(n_107),
.Y(n_149)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_16),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_106),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_48),
.B(n_9),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_43),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_108),
.A2(n_109),
.B1(n_49),
.B2(n_47),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_43),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_118),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_107),
.B(n_48),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_123),
.B(n_132),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_106),
.B(n_53),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_126),
.B(n_140),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_71),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_56),
.B(n_53),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_137),
.B(n_145),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_55),
.A2(n_109),
.B1(n_108),
.B2(n_104),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_138),
.A2(n_150),
.B1(n_159),
.B2(n_164),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_84),
.B(n_36),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_SL g141 ( 
.A1(n_100),
.A2(n_44),
.B(n_42),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_141),
.B(n_160),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_79),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_56),
.B(n_36),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_147),
.B(n_148),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_87),
.B(n_45),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_82),
.A2(n_51),
.B1(n_49),
.B2(n_47),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_154),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_63),
.A2(n_77),
.B1(n_99),
.B2(n_96),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_87),
.B(n_45),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_61),
.A2(n_50),
.B1(n_46),
.B2(n_19),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_163),
.B(n_167),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_66),
.A2(n_50),
.B1(n_46),
.B2(n_47),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_62),
.B(n_18),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_102),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_168),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_70),
.A2(n_49),
.B1(n_47),
.B2(n_43),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_176),
.A2(n_177),
.B1(n_42),
.B2(n_34),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_76),
.A2(n_49),
.B1(n_43),
.B2(n_27),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_166),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_179),
.Y(n_245)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_112),
.Y(n_180)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_180),
.Y(n_238)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_134),
.Y(n_181)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_181),
.Y(n_241)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_121),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_182),
.Y(n_250)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_116),
.Y(n_183)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_183),
.Y(n_235)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_116),
.Y(n_184)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_185),
.Y(n_273)
);

AO22x2_ASAP7_75t_L g186 ( 
.A1(n_141),
.A2(n_91),
.B1(n_89),
.B2(n_88),
.Y(n_186)
);

O2A1O1Ixp33_ASAP7_75t_SL g264 ( 
.A1(n_186),
.A2(n_159),
.B(n_119),
.C(n_128),
.Y(n_264)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_187),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_153),
.A2(n_83),
.B1(n_33),
.B2(n_29),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_188),
.A2(n_192),
.B1(n_197),
.B2(n_202),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_122),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_189),
.B(n_190),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_122),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_L g192 ( 
.A1(n_136),
.A2(n_33),
.B1(n_26),
.B2(n_29),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_193),
.Y(n_242)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_127),
.Y(n_195)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_195),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_139),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_196),
.B(n_199),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_120),
.A2(n_33),
.B1(n_26),
.B2(n_16),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_115),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_198),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_139),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_120),
.A2(n_33),
.B1(n_17),
.B2(n_20),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_127),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_203),
.Y(n_243)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_135),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_204),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_122),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_205),
.B(n_220),
.Y(n_252)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_124),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_206),
.Y(n_257)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_170),
.Y(n_209)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_209),
.Y(n_269)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_121),
.Y(n_210)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_210),
.Y(n_265)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_170),
.Y(n_211)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_124),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_212),
.Y(n_262)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_130),
.Y(n_213)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

BUFx2_ASAP7_75t_SL g216 ( 
.A(n_171),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_216),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_125),
.Y(n_217)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_217),
.Y(n_254)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_171),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_218),
.Y(n_270)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_110),
.Y(n_219)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_219),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_148),
.Y(n_220)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_125),
.Y(n_221)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_221),
.Y(n_266)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_157),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_223),
.Y(n_256)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_157),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_114),
.A2(n_22),
.B1(n_18),
.B2(n_19),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_225),
.A2(n_154),
.B1(n_177),
.B2(n_22),
.Y(n_251)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_144),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_228),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_150),
.Y(n_237)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_151),
.Y(n_228)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_151),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_229),
.B(n_230),
.Y(n_271)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_174),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_158),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_231),
.Y(n_272)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_175),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_232),
.A2(n_172),
.B1(n_171),
.B2(n_115),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_149),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_233),
.B(n_249),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_237),
.A2(n_251),
.B1(n_263),
.B2(n_264),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_208),
.A2(n_163),
.B(n_118),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_248),
.A2(n_274),
.B(n_129),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_215),
.B(n_146),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_200),
.B(n_117),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_258),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_194),
.A2(n_128),
.B1(n_173),
.B2(n_162),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_267),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_215),
.A2(n_165),
.B(n_131),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_264),
.A2(n_186),
.B1(n_201),
.B2(n_191),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_276),
.A2(n_280),
.B1(n_289),
.B2(n_247),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_248),
.B(n_192),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_277),
.Y(n_321)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_244),
.Y(n_278)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_278),
.Y(n_311)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_259),
.Y(n_279)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_279),
.Y(n_316)
);

OAI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_264),
.A2(n_191),
.B1(n_186),
.B2(n_225),
.Y(n_280)
);

OAI22x1_ASAP7_75t_L g281 ( 
.A1(n_251),
.A2(n_186),
.B1(n_178),
.B2(n_188),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g332 ( 
.A1(n_281),
.A2(n_285),
.B1(n_229),
.B2(n_228),
.Y(n_332)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_259),
.Y(n_283)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_283),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_246),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_284),
.B(n_288),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_263),
.A2(n_193),
.B1(n_156),
.B2(n_219),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_233),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_286),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_249),
.A2(n_224),
.B(n_207),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_287),
.A2(n_296),
.B(n_297),
.Y(n_327)
);

OAI32xp33_ASAP7_75t_L g288 ( 
.A1(n_258),
.A2(n_214),
.A3(n_202),
.B1(n_197),
.B2(n_142),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_239),
.A2(n_133),
.B1(n_162),
.B2(n_173),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_290),
.B(n_292),
.Y(n_323)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_256),
.Y(n_291)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_291),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_262),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_252),
.B(n_184),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_293),
.B(n_294),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_236),
.B(n_185),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_250),
.Y(n_295)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_295),
.Y(n_325)
);

A2O1A1Ixp33_ASAP7_75t_SL g297 ( 
.A1(n_237),
.A2(n_218),
.B(n_198),
.C(n_172),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_244),
.Y(n_298)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_298),
.Y(n_328)
);

INVx13_ASAP7_75t_L g299 ( 
.A(n_269),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_299),
.B(n_304),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_237),
.A2(n_129),
.B(n_155),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_307),
.Y(n_310)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_235),
.Y(n_302)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_302),
.Y(n_333)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_262),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_261),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_305),
.B(n_306),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_260),
.Y(n_306)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_255),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_303),
.A2(n_239),
.B1(n_261),
.B2(n_133),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_308),
.A2(n_314),
.B1(n_334),
.B2(n_289),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_309),
.A2(n_332),
.B1(n_275),
.B2(n_290),
.Y(n_347)
);

NOR2x1_ASAP7_75t_L g312 ( 
.A(n_277),
.B(n_270),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_312),
.B(n_313),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_279),
.B(n_270),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_303),
.A2(n_266),
.B1(n_245),
.B2(n_243),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_282),
.B(n_236),
.Y(n_317)
);

AO21x1_ASAP7_75t_L g350 ( 
.A1(n_317),
.A2(n_288),
.B(n_297),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_286),
.B(n_245),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_319),
.B(n_326),
.C(n_330),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_283),
.B(n_272),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_320),
.B(n_335),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_301),
.B(n_234),
.C(n_235),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_286),
.B(n_111),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_281),
.A2(n_266),
.B1(n_254),
.B2(n_210),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_301),
.B(n_272),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_296),
.B(n_257),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_337),
.B(n_277),
.Y(n_342)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_325),
.Y(n_338)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_338),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_325),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_340),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_341),
.A2(n_349),
.B1(n_366),
.B2(n_332),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_342),
.B(n_355),
.Y(n_390)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_320),
.Y(n_343)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_343),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_337),
.B(n_287),
.C(n_276),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_346),
.B(n_351),
.C(n_353),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_347),
.A2(n_362),
.B1(n_334),
.B2(n_322),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_313),
.B(n_335),
.Y(n_348)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_348),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_308),
.A2(n_275),
.B1(n_300),
.B2(n_291),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_350),
.B(n_352),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_337),
.B(n_306),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_309),
.A2(n_284),
.B1(n_297),
.B2(n_305),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_319),
.B(n_234),
.C(n_292),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_336),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_354),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_330),
.B(n_297),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_312),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_356),
.B(n_361),
.Y(n_384)
);

NAND2x1_ASAP7_75t_L g357 ( 
.A(n_312),
.B(n_321),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_357),
.A2(n_310),
.B(n_321),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_336),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_358),
.Y(n_379)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_316),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_359),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_317),
.B(n_253),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_360),
.B(n_363),
.Y(n_374)
);

AND2x2_ASAP7_75t_SL g361 ( 
.A(n_327),
.B(n_297),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_318),
.A2(n_295),
.B1(n_254),
.B2(n_250),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_323),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_316),
.B(n_302),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_364),
.B(n_322),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_315),
.B(n_307),
.C(n_240),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_365),
.B(n_323),
.C(n_331),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_314),
.A2(n_295),
.B1(n_250),
.B2(n_265),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_339),
.B(n_327),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_367),
.B(n_377),
.C(n_378),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_370),
.A2(n_396),
.B1(n_366),
.B2(n_364),
.Y(n_411)
);

OA21x2_ASAP7_75t_L g372 ( 
.A1(n_344),
.A2(n_318),
.B(n_310),
.Y(n_372)
);

OA22x2_ASAP7_75t_L g409 ( 
.A1(n_372),
.A2(n_357),
.B1(n_350),
.B2(n_352),
.Y(n_409)
);

CKINVDCx14_ASAP7_75t_R g418 ( 
.A(n_375),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_339),
.B(n_326),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_346),
.B(n_351),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_354),
.B(n_324),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_382),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_342),
.B(n_329),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_383),
.B(n_386),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_385),
.B(n_340),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_355),
.B(n_329),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_387),
.A2(n_389),
.B1(n_391),
.B2(n_394),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_388),
.B(n_392),
.C(n_365),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_341),
.A2(n_321),
.B1(n_324),
.B2(n_331),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_343),
.A2(n_333),
.B1(n_328),
.B2(n_311),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_353),
.B(n_333),
.C(n_328),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_338),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_393),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_349),
.A2(n_311),
.B1(n_265),
.B2(n_304),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_347),
.A2(n_268),
.B1(n_253),
.B2(n_242),
.Y(n_396)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_395),
.Y(n_399)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_399),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_419),
.C(n_423),
.Y(n_426)
);

INVx5_ASAP7_75t_L g402 ( 
.A(n_393),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_402),
.B(n_404),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_L g403 ( 
.A1(n_376),
.A2(n_358),
.B1(n_363),
.B2(n_359),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_403),
.A2(n_413),
.B1(n_424),
.B2(n_269),
.Y(n_447)
);

NOR3xp33_ASAP7_75t_L g404 ( 
.A(n_379),
.B(n_361),
.C(n_344),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_377),
.B(n_361),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_405),
.B(n_421),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_384),
.A2(n_356),
.B(n_357),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_407),
.B(n_410),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_372),
.B(n_348),
.Y(n_408)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_408),
.Y(n_428)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_409),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_374),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_411),
.A2(n_425),
.B1(n_373),
.B2(n_396),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_372),
.B(n_345),
.Y(n_412)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_412),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_387),
.A2(n_345),
.B1(n_268),
.B2(n_340),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_380),
.Y(n_414)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_414),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_388),
.B(n_298),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_415),
.B(n_420),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_417),
.B(n_422),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_392),
.B(n_369),
.C(n_367),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_380),
.B(n_240),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_391),
.B(n_278),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_384),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_369),
.B(n_273),
.C(n_269),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_368),
.Y(n_424)
);

OAI22xp33_ASAP7_75t_SL g425 ( 
.A1(n_381),
.A2(n_255),
.B1(n_242),
.B2(n_221),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_401),
.A2(n_371),
.B1(n_370),
.B2(n_385),
.Y(n_431)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_431),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_419),
.B(n_378),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_432),
.B(n_433),
.C(n_434),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_400),
.B(n_386),
.C(n_383),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_423),
.B(n_389),
.C(n_371),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_397),
.B(n_390),
.C(n_394),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_436),
.B(n_445),
.C(n_449),
.Y(n_461)
);

INVx13_ASAP7_75t_L g437 ( 
.A(n_402),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_437),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_401),
.A2(n_413),
.B1(n_422),
.B2(n_414),
.Y(n_441)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_441),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_443),
.A2(n_438),
.B1(n_421),
.B2(n_435),
.Y(n_454)
);

NOR2xp67_ASAP7_75t_SL g444 ( 
.A(n_406),
.B(n_390),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_444),
.B(n_398),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_397),
.B(n_368),
.C(n_273),
.Y(n_445)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_447),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_417),
.A2(n_217),
.B1(n_182),
.B2(n_238),
.Y(n_448)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_448),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_405),
.B(n_241),
.C(n_238),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_440),
.B(n_418),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_450),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_430),
.B(n_399),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_451),
.B(n_457),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_454),
.B(n_20),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_455),
.B(n_468),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_428),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_442),
.A2(n_407),
.B(n_431),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_458),
.A2(n_169),
.B(n_17),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_441),
.A2(n_409),
.B1(n_424),
.B2(n_416),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_463),
.A2(n_465),
.B1(n_466),
.B2(n_452),
.Y(n_477)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_427),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_464),
.B(n_467),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_439),
.A2(n_442),
.B1(n_448),
.B2(n_429),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_442),
.A2(n_409),
.B1(n_416),
.B2(n_398),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_446),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_437),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_426),
.B(n_445),
.C(n_432),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_469),
.B(n_241),
.C(n_211),
.Y(n_476)
);

OAI321xp33_ASAP7_75t_L g470 ( 
.A1(n_451),
.A2(n_409),
.A3(n_443),
.B1(n_434),
.B2(n_429),
.C(n_449),
.Y(n_470)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_470),
.Y(n_490)
);

FAx1_ASAP7_75t_SL g471 ( 
.A(n_466),
.B(n_433),
.CI(n_436),
.CON(n_471),
.SN(n_471)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_471),
.B(n_476),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_458),
.A2(n_426),
.B(n_299),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_472),
.A2(n_481),
.B(n_8),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_461),
.B(n_299),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_475),
.B(n_477),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_479),
.A2(n_10),
.B(n_15),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_469),
.A2(n_209),
.B(n_143),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_453),
.B(n_143),
.C(n_113),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_482),
.B(n_486),
.C(n_487),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_450),
.B(n_34),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_483),
.B(n_484),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_461),
.B(n_155),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_485),
.B(n_456),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_465),
.B(n_113),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_454),
.B(n_161),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_474),
.A2(n_452),
.B1(n_459),
.B2(n_463),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_491),
.B(n_496),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_480),
.Y(n_493)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_493),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_478),
.A2(n_456),
.B1(n_460),
.B2(n_462),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_494),
.A2(n_498),
.B1(n_489),
.B2(n_14),
.Y(n_514)
);

OAI21x1_ASAP7_75t_L g495 ( 
.A1(n_473),
.A2(n_453),
.B(n_462),
.Y(n_495)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_495),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_475),
.B(n_460),
.C(n_161),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_497),
.B(n_503),
.Y(n_511)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_499),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_476),
.B(n_10),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_500),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_SL g501 ( 
.A(n_471),
.B(n_11),
.Y(n_501)
);

XNOR2x1_ASAP7_75t_L g513 ( 
.A(n_501),
.B(n_5),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_502),
.B(n_8),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_484),
.B(n_482),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_490),
.A2(n_485),
.B(n_479),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_504),
.B(n_507),
.Y(n_521)
);

OAI221xp5_ASAP7_75t_L g505 ( 
.A1(n_501),
.A2(n_471),
.B1(n_488),
.B2(n_492),
.C(n_499),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_505),
.B(n_514),
.Y(n_520)
);

AOI21x1_ASAP7_75t_SL g506 ( 
.A1(n_497),
.A2(n_487),
.B(n_486),
.Y(n_506)
);

AOI21x1_ASAP7_75t_SL g523 ( 
.A1(n_506),
.A2(n_509),
.B(n_513),
.Y(n_523)
);

AO22x1_ASAP7_75t_L g509 ( 
.A1(n_498),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_489),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_512),
.A2(n_3),
.B1(n_12),
.B2(n_2),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_SL g524 ( 
.A(n_513),
.B(n_12),
.Y(n_524)
);

NOR2xp67_ASAP7_75t_SL g518 ( 
.A(n_516),
.B(n_3),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_518),
.A2(n_517),
.B(n_508),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_515),
.B(n_35),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_519),
.B(n_522),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_523),
.B(n_524),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_511),
.B(n_44),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_525),
.B(n_526),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_511),
.B(n_44),
.C(n_35),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_527),
.B(n_528),
.C(n_530),
.Y(n_534)
);

FAx1_ASAP7_75t_SL g528 ( 
.A(n_521),
.B(n_510),
.CI(n_509),
.CON(n_528),
.SN(n_528)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_520),
.A2(n_506),
.B(n_44),
.Y(n_530)
);

INVxp33_ASAP7_75t_L g533 ( 
.A(n_532),
.Y(n_533)
);

NAND4xp25_ASAP7_75t_L g538 ( 
.A(n_533),
.B(n_535),
.C(n_35),
.D(n_1),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_529),
.A2(n_520),
.B(n_35),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_531),
.B(n_44),
.C(n_35),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_536),
.B(n_531),
.C(n_44),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_537),
.B(n_538),
.C(n_534),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_539),
.B(n_0),
.C(n_1),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_540),
.A2(n_2),
.B(n_0),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_541),
.B(n_0),
.C(n_1),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_542),
.B(n_1),
.Y(n_543)
);


endmodule