module fake_jpeg_26056_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_288;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_5),
.B(n_14),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_14),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g33 ( 
.A(n_16),
.Y(n_33)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_39),
.Y(n_44)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_41),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_42),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_43),
.B(n_48),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_49),
.Y(n_72)
);

CKINVDCx12_ASAP7_75t_R g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_57),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_33),
.A2(n_15),
.B1(n_21),
.B2(n_30),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_51),
.A2(n_55),
.B1(n_26),
.B2(n_30),
.Y(n_75)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_15),
.B1(n_21),
.B2(n_22),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_54),
.A2(n_22),
.B1(n_24),
.B2(n_41),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_33),
.A2(n_38),
.B1(n_37),
.B2(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_39),
.B(n_19),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_18),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_63),
.A2(n_11),
.B(n_14),
.Y(n_88)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_44),
.A2(n_38),
.B1(n_33),
.B2(n_34),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_70),
.B1(n_52),
.B2(n_53),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_38),
.B1(n_33),
.B2(n_34),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_36),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_71),
.A2(n_74),
.B(n_79),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_36),
.C(n_32),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_56),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_36),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_75),
.A2(n_76),
.B1(n_61),
.B2(n_43),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_52),
.A2(n_26),
.B1(n_23),
.B2(n_28),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_32),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_86),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_66),
.Y(n_102)
);

AOI22x1_ASAP7_75t_SL g83 ( 
.A1(n_50),
.A2(n_41),
.B1(n_40),
.B2(n_22),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_45),
.B(n_66),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_12),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_85),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_90),
.B(n_97),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_92),
.A2(n_108),
.B1(n_109),
.B2(n_68),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_59),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_102),
.Y(n_119)
);

OAI32xp33_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_60),
.A3(n_45),
.B1(n_48),
.B2(n_65),
.Y(n_95)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_96),
.A2(n_99),
.B(n_107),
.Y(n_121)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_98),
.B(n_104),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_73),
.A2(n_61),
.B1(n_58),
.B2(n_66),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_112),
.B1(n_74),
.B2(n_70),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_87),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_79),
.B(n_56),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_106),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_85),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_79),
.B(n_56),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_71),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_83),
.A2(n_41),
.B1(n_40),
.B2(n_61),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_0),
.B(n_1),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_110),
.A2(n_74),
.B(n_67),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_110),
.B(n_94),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_80),
.A2(n_56),
.B1(n_29),
.B2(n_31),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_114),
.B(n_132),
.Y(n_139)
);

OA21x2_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_88),
.B(n_80),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_99),
.B(n_106),
.Y(n_143)
);

BUFx8_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_107),
.A2(n_78),
.B1(n_74),
.B2(n_77),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_117),
.A2(n_122),
.B(n_125),
.Y(n_144)
);

BUFx24_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_69),
.B1(n_86),
.B2(n_81),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_123),
.A2(n_112),
.B1(n_109),
.B2(n_102),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_92),
.B1(n_107),
.B2(n_98),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_77),
.B(n_72),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_69),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_130),
.Y(n_146)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_134),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_31),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_92),
.Y(n_142)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_133),
.B(n_135),
.Y(n_153)
);

BUFx24_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_27),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_112),
.Y(n_152)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_102),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_140),
.A2(n_142),
.B1(n_159),
.B2(n_135),
.Y(n_166)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_141),
.B(n_145),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_143),
.A2(n_157),
.B(n_158),
.Y(n_182)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_97),
.C(n_104),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_136),
.C(n_125),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_113),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_148),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_126),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_149),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_118),
.A2(n_111),
.B(n_108),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_150),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_122),
.Y(n_176)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_155),
.Y(n_172)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_160),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_115),
.A2(n_68),
.B(n_89),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_115),
.A2(n_89),
.B(n_72),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_133),
.A2(n_24),
.B1(n_20),
.B2(n_27),
.Y(n_159)
);

AND2x6_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_9),
.Y(n_160)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_163),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_164),
.B(n_175),
.C(n_179),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_166),
.A2(n_151),
.B1(n_163),
.B2(n_154),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_139),
.B(n_119),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_167),
.B(n_169),
.Y(n_200)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_177),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_148),
.B(n_119),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_147),
.B(n_132),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_174),
.B(n_176),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_137),
.C(n_128),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_186),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_128),
.C(n_118),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_142),
.A2(n_134),
.B1(n_120),
.B2(n_117),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_181),
.A2(n_158),
.B1(n_157),
.B2(n_145),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_161),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_184),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_149),
.B(n_120),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_185),
.B(n_187),
.Y(n_209)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_138),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

XOR2x2_ASAP7_75t_L g188 ( 
.A(n_144),
.B(n_134),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_188),
.A2(n_171),
.B(n_144),
.Y(n_199)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_183),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_191),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_181),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_196),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_187),
.Y(n_196)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_20),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_28),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_175),
.Y(n_202)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_173),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_203),
.Y(n_219)
);

NAND2x1_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_162),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_197),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_186),
.A2(n_142),
.B1(n_134),
.B2(n_160),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_205),
.A2(n_210),
.B1(n_211),
.B2(n_171),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_152),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_165),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_170),
.A2(n_159),
.B1(n_162),
.B2(n_120),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_180),
.A2(n_161),
.B1(n_24),
.B2(n_116),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_179),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_174),
.Y(n_217)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_204),
.Y(n_214)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_214),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_215),
.A2(n_206),
.B(n_194),
.Y(n_245)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_216),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_220),
.C(n_221),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_164),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_224),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_182),
.C(n_168),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_182),
.C(n_177),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_178),
.C(n_165),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_227),
.C(n_221),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_205),
.A2(n_173),
.B1(n_189),
.B2(n_116),
.Y(n_226)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_84),
.C(n_62),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_200),
.B(n_9),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_230),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_191),
.Y(n_237)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_215),
.A2(n_198),
.B1(n_192),
.B2(n_204),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_238),
.A2(n_241),
.B1(n_249),
.B2(n_0),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_222),
.A2(n_196),
.B1(n_190),
.B2(n_199),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_209),
.Y(n_244)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_244),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_245),
.A2(n_6),
.B(n_13),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_84),
.C(n_46),
.Y(n_259)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_247),
.B(n_248),
.Y(n_253)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_222),
.A2(n_195),
.B1(n_194),
.B2(n_206),
.Y(n_249)
);

OAI21xp33_ASAP7_75t_L g250 ( 
.A1(n_234),
.A2(n_225),
.B(n_214),
.Y(n_250)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_240),
.B(n_229),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_251),
.Y(n_273)
);

A2O1A1O1Ixp25_ASAP7_75t_L g252 ( 
.A1(n_245),
.A2(n_224),
.B(n_220),
.C(n_223),
.D(n_227),
.Y(n_252)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_252),
.Y(n_270)
);

AOI322xp5_ASAP7_75t_SL g254 ( 
.A1(n_244),
.A2(n_7),
.A3(n_13),
.B1(n_12),
.B2(n_10),
.C1(n_8),
.C2(n_5),
.Y(n_254)
);

NOR2xp67_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_6),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_7),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_255),
.A2(n_10),
.B(n_8),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_235),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_257),
.B(n_259),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_84),
.C(n_62),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_233),
.C(n_62),
.Y(n_274)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_262),
.Y(n_272)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_237),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_263),
.A2(n_243),
.B(n_239),
.Y(n_267)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_264),
.Y(n_275)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_267),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_268),
.B(n_255),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_258),
.A2(n_242),
.B1(n_236),
.B2(n_238),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_274),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g271 ( 
.A(n_252),
.B(n_235),
.CI(n_242),
.CON(n_271),
.SN(n_271)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_260),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_276),
.B(n_254),
.Y(n_279)
);

OAI21x1_ASAP7_75t_L g277 ( 
.A1(n_265),
.A2(n_253),
.B(n_250),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_277),
.A2(n_266),
.B1(n_269),
.B2(n_274),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_279),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_280),
.A2(n_283),
.B(n_271),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_256),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_282),
.B(n_284),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_6),
.B(n_8),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_1),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_288),
.Y(n_292)
);

AOI21x1_ASAP7_75t_L g289 ( 
.A1(n_285),
.A2(n_271),
.B(n_267),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_289),
.A2(n_278),
.B1(n_272),
.B2(n_3),
.Y(n_294)
);

BUFx24_ASAP7_75t_SL g293 ( 
.A(n_290),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_281),
.B(n_275),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_1),
.C(n_2),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_295),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_292),
.A2(n_286),
.B(n_287),
.Y(n_297)
);

OAI321xp33_ASAP7_75t_L g298 ( 
.A1(n_297),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_293),
.C(n_296),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_2),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_4),
.Y(n_300)
);


endmodule