module fake_jpeg_904_n_121 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_121);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx5_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_46),
.Y(n_56)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_48),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_28),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_32),
.B1(n_41),
.B2(n_39),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_52),
.A2(n_56),
.B1(n_49),
.B2(n_54),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_1),
.Y(n_70)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

OAI21xp33_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_59),
.B(n_37),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_32),
.B1(n_38),
.B2(n_33),
.Y(n_57)
);

OAI22x1_ASAP7_75t_SL g62 ( 
.A1(n_57),
.A2(n_33),
.B1(n_36),
.B2(n_34),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_40),
.Y(n_59)
);

AOI32xp33_ASAP7_75t_L g60 ( 
.A1(n_50),
.A2(n_53),
.A3(n_59),
.B1(n_46),
.B2(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_69),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_57),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_61),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_63),
.B1(n_64),
.B2(n_58),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_50),
.B1(n_52),
.B2(n_49),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_56),
.B(n_36),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_66),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_56),
.B(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_68),
.Y(n_83)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_51),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_3),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_27),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_2),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_81),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_55),
.C(n_54),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_75),
.C(n_80),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_55),
.B(n_58),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_58),
.B(n_62),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_79),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_4),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_4),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_54),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_94),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_11),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_87),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_89),
.C(n_91),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_25),
.C(n_24),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_90),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_76),
.C(n_83),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_23),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_93),
.B(n_10),
.Y(n_98)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_9),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_95),
.B(n_17),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_15),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_99),
.A2(n_101),
.B(n_104),
.Y(n_107)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_102),
.A2(n_105),
.B1(n_92),
.B2(n_16),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_13),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_91),
.A2(n_15),
.B1(n_16),
.B2(n_19),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_93),
.C(n_89),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_108),
.A2(n_111),
.B(n_105),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_96),
.Y(n_115)
);

AOI322xp5_ASAP7_75t_L g113 ( 
.A1(n_107),
.A2(n_99),
.A3(n_103),
.B1(n_96),
.B2(n_102),
.C1(n_20),
.C2(n_22),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_113),
.B(n_109),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_115),
.A2(n_116),
.B(n_114),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_115),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_108),
.C(n_111),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_119),
.B(n_110),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_106),
.Y(n_121)
);


endmodule