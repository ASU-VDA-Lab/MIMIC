module fake_jpeg_628_n_216 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_216);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_10),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_2),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_8),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_35),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_24),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_30),
.B(n_29),
.Y(n_74)
);

BUFx24_ASAP7_75t_L g75 ( 
.A(n_8),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_0),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_L g88 ( 
.A1(n_77),
.A2(n_83),
.B(n_74),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_75),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_79),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_20),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_56),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_81),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_49),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_85),
.A2(n_60),
.B1(n_75),
.B2(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_88),
.Y(n_105)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_85),
.B1(n_79),
.B2(n_59),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_65),
.B1(n_53),
.B2(n_57),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_73),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_95),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_51),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_69),
.B1(n_72),
.B2(n_53),
.Y(n_96)
);

AO22x1_ASAP7_75t_SL g101 ( 
.A1(n_96),
.A2(n_83),
.B1(n_65),
.B2(n_72),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_84),
.B1(n_69),
.B2(n_61),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_61),
.Y(n_116)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_100),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_101),
.A2(n_117),
.B1(n_116),
.B2(n_92),
.Y(n_125)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_114),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_118),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_68),
.B(n_62),
.Y(n_129)
);

NOR2x1_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_52),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_101),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_122),
.A2(n_136),
.B1(n_4),
.B2(n_5),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_125),
.A2(n_25),
.B1(n_45),
.B2(n_44),
.Y(n_148)
);

BUFx12_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_126),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_105),
.C(n_55),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_134),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_129),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_71),
.B(n_70),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_3),
.B(n_4),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_66),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_135),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_67),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_133),
.B(n_32),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_57),
.C(n_50),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_0),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_112),
.A2(n_68),
.B1(n_62),
.B2(n_76),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_1),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_5),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_122),
.B(n_125),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_143),
.A2(n_146),
.B(n_27),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_126),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_149),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_68),
.B(n_76),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_138),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_148),
.B1(n_156),
.B2(n_167),
.Y(n_178)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_140),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_151),
.Y(n_172)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_126),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_153),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_127),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_158),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_6),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_160),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_134),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_128),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_165),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_123),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_36),
.C(n_43),
.Y(n_171)
);

AOI32xp33_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_7),
.A3(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_164),
.A2(n_13),
.B(n_14),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_7),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_166),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_125),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_47),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_173),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_177),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_175),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_33),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_181),
.B1(n_149),
.B2(n_147),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_39),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_157),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_179),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_143),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_188),
.Y(n_197)
);

OAI21xp33_ASAP7_75t_SL g188 ( 
.A1(n_168),
.A2(n_162),
.B(n_146),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_184),
.B(n_145),
.Y(n_189)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_189),
.Y(n_196)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_176),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_192),
.A2(n_180),
.B1(n_183),
.B2(n_181),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_156),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_171),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_193),
.B(n_173),
.C(n_169),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_200),
.C(n_201),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_188),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_198),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_175),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_202),
.C(n_185),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_191),
.C(n_187),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_205),
.B(n_196),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_197),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_207),
.A2(n_208),
.B1(n_198),
.B2(n_204),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_209),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_203),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_174),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_178),
.C(n_19),
.Y(n_213)
);

BUFx24_ASAP7_75t_SL g214 ( 
.A(n_213),
.Y(n_214)
);

BUFx24_ASAP7_75t_SL g215 ( 
.A(n_214),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_178),
.Y(n_216)
);


endmodule