module fake_jpeg_28456_n_320 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_42),
.Y(n_67)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_48),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

CKINVDCx6p67_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_26),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx5_ASAP7_75t_SL g53 ( 
.A(n_49),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_50),
.B(n_51),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_32),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_18),
.B1(n_23),
.B2(n_27),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_52),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_88)
);

INVx5_ASAP7_75t_SL g54 ( 
.A(n_46),
.Y(n_54)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_49),
.A2(n_17),
.B1(n_33),
.B2(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_34),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_57),
.B(n_35),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_17),
.B1(n_33),
.B2(n_30),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_46),
.A2(n_17),
.B1(n_33),
.B2(n_30),
.Y(n_59)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_17),
.B1(n_33),
.B2(n_30),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_63),
.A2(n_71),
.B1(n_80),
.B2(n_29),
.Y(n_92)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_47),
.A2(n_17),
.B1(n_23),
.B2(n_18),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_74),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_40),
.A2(n_27),
.B1(n_23),
.B2(n_18),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_67),
.B(n_38),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_82),
.Y(n_124)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_67),
.B(n_38),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_85),
.B(n_87),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_43),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_89),
.B(n_93),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_64),
.A2(n_43),
.B(n_44),
.C(n_42),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_90),
.B(n_66),
.Y(n_123)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_92),
.A2(n_27),
.B1(n_23),
.B2(n_75),
.Y(n_129)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

AND2x4_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_19),
.Y(n_94)
);

OR2x4_ASAP7_75t_L g145 ( 
.A(n_94),
.B(n_19),
.Y(n_145)
);

AOI21xp33_ASAP7_75t_L g95 ( 
.A1(n_64),
.A2(n_37),
.B(n_22),
.Y(n_95)
);

AOI21xp33_ASAP7_75t_L g127 ( 
.A1(n_95),
.A2(n_101),
.B(n_20),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_44),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_117),
.C(n_36),
.Y(n_134)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

OR2x2_ASAP7_75t_SL g101 ( 
.A(n_76),
.B(n_27),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_53),
.A2(n_42),
.B(n_34),
.C(n_28),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_70),
.Y(n_121)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_53),
.B(n_37),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_110),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g112 ( 
.A(n_55),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_112),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_61),
.B(n_28),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_22),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_60),
.B(n_35),
.C(n_24),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_137),
.Y(n_154)
);

NOR2xp67_ASAP7_75t_R g172 ( 
.A(n_121),
.B(n_123),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_105),
.B(n_24),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_122),
.B(n_151),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_127),
.A2(n_130),
.B(n_145),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_101),
.A2(n_65),
.B1(n_69),
.B2(n_72),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_88),
.B1(n_83),
.B2(n_84),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_129),
.A2(n_115),
.B1(n_99),
.B2(n_118),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_94),
.A2(n_55),
.B(n_19),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_132),
.B(n_134),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_68),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_138),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_102),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_68),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_68),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_143),
.Y(n_165)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_90),
.B(n_55),
.C(n_36),
.Y(n_143)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_86),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_148),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_20),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_114),
.B(n_8),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_98),
.B(n_19),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_99),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_156),
.A2(n_139),
.B1(n_143),
.B2(n_138),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_157),
.A2(n_160),
.B1(n_161),
.B2(n_169),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_112),
.B(n_98),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_158),
.A2(n_185),
.B(n_147),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_137),
.A2(n_111),
.B1(n_84),
.B2(n_103),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_121),
.A2(n_103),
.B1(n_97),
.B2(n_107),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_149),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_167),
.B(n_175),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_121),
.A2(n_107),
.B1(n_104),
.B2(n_113),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_171),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_86),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_129),
.A2(n_104),
.B1(n_118),
.B2(n_91),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_173),
.A2(n_140),
.B1(n_141),
.B2(n_125),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_126),
.B(n_124),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_122),
.B(n_7),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_176),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_11),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_180),
.Y(n_187)
);

AOI22x1_ASAP7_75t_SL g178 ( 
.A1(n_145),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_178),
.A2(n_125),
.B(n_135),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_0),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_181),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_11),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_124),
.B(n_0),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_12),
.Y(n_182)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_133),
.B(n_2),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_144),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_130),
.A2(n_2),
.B(n_3),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_149),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_186),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_188),
.A2(n_190),
.B1(n_196),
.B2(n_202),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_183),
.B(n_155),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_211),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_156),
.A2(n_126),
.B1(n_134),
.B2(n_130),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_191),
.A2(n_178),
.B(n_185),
.Y(n_229)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_193),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_195),
.B(n_201),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_156),
.A2(n_128),
.B1(n_153),
.B2(n_131),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_136),
.C(n_144),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_155),
.C(n_159),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_154),
.A2(n_119),
.B1(n_131),
.B2(n_136),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_154),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_207),
.Y(n_239)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_168),
.Y(n_206)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_206),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_172),
.A2(n_119),
.B(n_147),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_208),
.A2(n_181),
.B(n_160),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_170),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_210),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_158),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_165),
.B(n_152),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_173),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_172),
.Y(n_213)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_213),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_163),
.A2(n_146),
.B1(n_125),
.B2(n_135),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_214),
.A2(n_169),
.B1(n_157),
.B2(n_161),
.Y(n_223)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_160),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_215),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_216),
.A2(n_166),
.B(n_174),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_199),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_222),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_219),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_205),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_230),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_183),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_229),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_228),
.C(n_233),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_159),
.C(n_163),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_205),
.Y(n_230)
);

A2O1A1O1Ixp25_ASAP7_75t_L g231 ( 
.A1(n_208),
.A2(n_171),
.B(n_184),
.C(n_185),
.D(n_178),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_234),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_210),
.A2(n_162),
.B(n_175),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_194),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_186),
.C(n_167),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_190),
.B(n_166),
.C(n_177),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_188),
.C(n_191),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_214),
.B1(n_215),
.B2(n_213),
.Y(n_255)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_239),
.Y(n_241)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_242),
.A2(n_254),
.B(n_249),
.Y(n_273)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_250),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_226),
.C(n_235),
.Y(n_261)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_227),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_247),
.Y(n_260)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_240),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_251),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_187),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_253),
.B(n_232),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_225),
.A2(n_195),
.B1(n_207),
.B2(n_213),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_255),
.A2(n_256),
.B1(n_258),
.B2(n_259),
.Y(n_262)
);

INVx3_ASAP7_75t_SL g256 ( 
.A(n_219),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_225),
.A2(n_197),
.B1(n_198),
.B2(n_204),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_237),
.A2(n_197),
.B1(n_201),
.B2(n_206),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_272),
.C(n_277),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_243),
.A2(n_176),
.B(n_164),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_263),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_269),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_224),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_268),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_221),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_246),
.A2(n_164),
.B(n_220),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_245),
.B(n_179),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_192),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_221),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_259),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_228),
.C(n_217),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_273),
.A2(n_275),
.B1(n_212),
.B2(n_247),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_258),
.A2(n_217),
.B1(n_223),
.B2(n_219),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_236),
.C(n_234),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_271),
.C(n_272),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_268),
.C(n_266),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_192),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_284),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_276),
.A2(n_257),
.B(n_255),
.Y(n_283)
);

A2O1A1O1Ixp25_ASAP7_75t_L g293 ( 
.A1(n_283),
.A2(n_276),
.B(n_229),
.C(n_277),
.D(n_274),
.Y(n_293)
);

NOR3xp33_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_216),
.C(n_231),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_262),
.A2(n_256),
.B1(n_257),
.B2(n_220),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_193),
.C(n_260),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_267),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_286),
.B(n_274),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_288),
.A2(n_289),
.B1(n_146),
.B2(n_14),
.Y(n_298)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_260),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_294),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_293),
.A2(n_296),
.B1(n_298),
.B2(n_283),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_280),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_278),
.B(n_174),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_299),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_290),
.B(n_13),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_292),
.B(n_279),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_300),
.A2(n_306),
.B(n_307),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_302),
.A2(n_5),
.B1(n_14),
.B2(n_15),
.Y(n_312)
);

NOR3xp33_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_279),
.C(n_289),
.Y(n_304)
);

AOI21xp33_ASAP7_75t_L g309 ( 
.A1(n_304),
.A2(n_285),
.B(n_287),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_135),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_294),
.B(n_281),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_292),
.B(n_287),
.Y(n_307)
);

AOI322xp5_ASAP7_75t_L g314 ( 
.A1(n_309),
.A2(n_311),
.A3(n_312),
.B1(n_303),
.B2(n_14),
.C1(n_15),
.C2(n_16),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_310),
.A2(n_303),
.B(n_5),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_301),
.A2(n_5),
.B(n_11),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_313),
.B(n_314),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_308),
.A2(n_3),
.A3(n_4),
.B1(n_15),
.B2(n_16),
.C1(n_310),
.C2(n_274),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_315),
.B(n_16),
.C(n_3),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_317),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_316),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_3),
.Y(n_320)
);


endmodule