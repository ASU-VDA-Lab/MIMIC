module real_jpeg_11998_n_17 (n_5, n_4, n_8, n_0, n_12, n_324, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_324;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g98 ( 
.A(n_0),
.Y(n_98)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_3),
.A2(n_40),
.B1(n_41),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_3),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_3),
.A2(n_28),
.B1(n_30),
.B2(n_81),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_3),
.A2(n_58),
.B1(n_62),
.B2(n_81),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_81),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_4),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_4),
.A2(n_28),
.B1(n_30),
.B2(n_43),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_43),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_4),
.A2(n_43),
.B1(n_58),
.B2(n_62),
.Y(n_268)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_6),
.A2(n_28),
.B1(n_30),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_6),
.A2(n_36),
.B1(n_58),
.B2(n_62),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_7),
.A2(n_40),
.B1(n_41),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_7),
.A2(n_28),
.B1(n_30),
.B2(n_50),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_50),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_7),
.A2(n_50),
.B1(n_58),
.B2(n_62),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_8),
.A2(n_40),
.B1(n_41),
.B2(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_8),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_110),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_8),
.A2(n_58),
.B1(n_62),
.B2(n_110),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_8),
.A2(n_28),
.B1(n_30),
.B2(n_110),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_9),
.A2(n_40),
.B1(n_41),
.B2(n_73),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_9),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_9),
.A2(n_28),
.B1(n_30),
.B2(n_73),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_73),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_9),
.A2(n_58),
.B1(n_62),
.B2(n_73),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_10),
.A2(n_40),
.B1(n_41),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_10),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_10),
.A2(n_58),
.B1(n_62),
.B2(n_144),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_144),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_10),
.A2(n_28),
.B1(n_30),
.B2(n_144),
.Y(n_254)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_12),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_12),
.A2(n_58),
.B1(n_62),
.B2(n_176),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_12),
.A2(n_28),
.B1(n_30),
.B2(n_176),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_12),
.A2(n_40),
.B1(n_41),
.B2(n_176),
.Y(n_278)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_164),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_14),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_14),
.B(n_58),
.C(n_61),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_14),
.B(n_31),
.Y(n_172)
);

OAI21xp33_ASAP7_75t_L g196 ( 
.A1(n_14),
.A2(n_135),
.B(n_180),
.Y(n_196)
);

O2A1O1Ixp33_ASAP7_75t_L g206 ( 
.A1(n_14),
.A2(n_27),
.B(n_30),
.C(n_207),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_14),
.A2(n_28),
.B1(n_30),
.B2(n_164),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_14),
.B(n_51),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_14),
.B(n_40),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_15),
.A2(n_28),
.B1(n_30),
.B2(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_15),
.A2(n_40),
.B1(n_41),
.B2(n_47),
.Y(n_48)
);

NAND2xp33_ASAP7_75t_SL g264 ( 
.A(n_15),
.B(n_28),
.Y(n_264)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_88),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_87),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_74),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_21),
.B(n_74),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_54),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_37),
.B1(n_52),
.B2(n_53),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_23),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_31),
.B(n_34),
.Y(n_23)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_24),
.A2(n_31),
.B1(n_84),
.B2(n_86),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_24),
.B(n_214),
.Y(n_228)
);

NOR2x1_ASAP7_75t_R g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_25)
);

AO22x1_ASAP7_75t_SL g31 ( 
.A1(n_26),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_L g207 ( 
.A1(n_26),
.A2(n_32),
.B(n_164),
.Y(n_207)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI32xp33_ASAP7_75t_L g263 ( 
.A1(n_30),
.A2(n_41),
.A3(n_47),
.B1(n_251),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_31),
.B(n_214),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_32),
.A2(n_33),
.B1(n_60),
.B2(n_61),
.Y(n_64)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_33),
.B(n_168),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_35),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_67)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_44),
.B1(n_49),
.B2(n_51),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_39),
.A2(n_45),
.B1(n_46),
.B2(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

O2A1O1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_41),
.A2(n_45),
.B(n_164),
.C(n_250),
.Y(n_249)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_44),
.B(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_46),
.B1(n_72),
.B2(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_45),
.A2(n_143),
.B(n_145),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_45),
.A2(n_46),
.B1(n_143),
.B2(n_278),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_48),
.Y(n_45)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_46),
.A2(n_80),
.B(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_46),
.B(n_109),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_46),
.A2(n_107),
.B(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_67),
.C(n_71),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_67),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_55),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_SL g82 ( 
.A(n_55),
.B(n_79),
.C(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_55),
.A2(n_78),
.B1(n_83),
.B2(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_63),
.B(n_65),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_56),
.A2(n_63),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_56),
.A2(n_63),
.B1(n_103),
.B2(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_56),
.B(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_56),
.A2(n_63),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_56),
.A2(n_63),
.B1(n_139),
.B2(n_257),
.Y(n_283)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_57),
.A2(n_66),
.B1(n_105),
.B2(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_57),
.A2(n_175),
.B(n_177),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_57),
.B(n_164),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_57),
.A2(n_177),
.B(n_256),
.Y(n_255)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_58),
.Y(n_62)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_62),
.B(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_62),
.B(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_63),
.B(n_166),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_68),
.A2(n_70),
.B1(n_85),
.B2(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_68),
.A2(n_70),
.B1(n_114),
.B2(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_68),
.A2(n_212),
.B(n_213),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_68),
.A2(n_70),
.B1(n_227),
.B2(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_68),
.A2(n_213),
.B(n_254),
.Y(n_276)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_70),
.A2(n_227),
.B(n_228),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_70),
.A2(n_141),
.B(n_228),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.C(n_82),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_75),
.A2(n_79),
.B1(n_118),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_75),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_79),
.A2(n_118),
.B1(n_119),
.B2(n_121),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_79),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_82),
.B(n_149),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_83),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AO21x1_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_152),
.B(n_320),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_147),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_122),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_91),
.B(n_122),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_111),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_92),
.B(n_112),
.C(n_117),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_96),
.B(n_106),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_93),
.A2(n_94),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_101),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_95),
.A2(n_96),
.B1(n_106),
.B2(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_95),
.A2(n_96),
.B1(n_101),
.B2(n_102),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_98),
.B(n_99),
.Y(n_96)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_97),
.A2(n_98),
.B1(n_185),
.B2(n_187),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_97),
.B(n_181),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_97),
.A2(n_98),
.B1(n_134),
.B2(n_268),
.Y(n_282)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_98),
.B(n_181),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_100),
.A2(n_133),
.B1(n_135),
.B2(n_136),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_117),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_113),
.B(n_115),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_116),
.A2(n_163),
.B(n_165),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_116),
.A2(n_165),
.B(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_119),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_128),
.C(n_129),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_123),
.A2(n_124),
.B1(n_128),
.B2(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_128),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_129),
.B(n_317),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_140),
.C(n_142),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_130),
.A2(n_131),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_137),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_132),
.A2(n_137),
.B1(n_138),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_132),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_135),
.A2(n_179),
.B(n_180),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_135),
.A2(n_136),
.B1(n_209),
.B2(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_135),
.A2(n_136),
.B1(n_234),
.B2(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_136),
.A2(n_186),
.B(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_136),
.B(n_164),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_136),
.A2(n_194),
.B(n_209),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_140),
.B(n_142),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_146),
.B(n_249),
.Y(n_248)
);

OAI21xp33_ASAP7_75t_L g320 ( 
.A1(n_147),
.A2(n_321),
.B(n_322),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_148),
.B(n_151),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_314),
.B(n_319),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_302),
.B(n_313),
.Y(n_153)
);

OAI321xp33_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_270),
.A3(n_295),
.B1(n_300),
.B2(n_301),
.C(n_324),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_243),
.B(n_269),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_221),
.B(n_242),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_202),
.B(n_220),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_182),
.B(n_201),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_169),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_160),
.B(n_169),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_167),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_161),
.A2(n_162),
.B1(n_167),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_167),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_178),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_174),
.C(n_178),
.Y(n_203)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_179),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_190),
.B(n_200),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_188),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_184),
.B(n_188),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_195),
.B(n_199),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_192),
.B(n_193),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_203),
.B(n_204),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_210),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_215),
.C(n_219),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_208),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_208),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_215),
.B1(n_218),
.B2(n_219),
.Y(n_210)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_211),
.Y(n_219)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_217),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_222),
.B(n_223),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_235),
.B2(n_236),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_238),
.C(n_240),
.Y(n_244)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_229),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_230),
.C(n_233),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_240),
.B2(n_241),
.Y(n_236)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_237),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_238),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_244),
.B(n_245),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_259),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_246),
.B(n_260),
.C(n_261),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_252),
.B2(n_258),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_247),
.B(n_253),
.C(n_255),
.Y(n_284)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_252),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_265),
.B2(n_266),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_266),
.Y(n_280)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_285),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_271),
.B(n_285),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_281),
.C(n_284),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_272),
.A2(n_273),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_280),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_277),
.B2(n_279),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_279),
.C(n_280),
.Y(n_294)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_277),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_281),
.B(n_284),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_283),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_294),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_289),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_287),
.B(n_289),
.C(n_294),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_293),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_292),
.C(n_293),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_296),
.B(n_297),
.Y(n_300)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_312),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_312),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_307),
.C(n_308),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_316),
.Y(n_319)
);


endmodule