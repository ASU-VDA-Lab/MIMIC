module fake_jpeg_5863_n_324 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx11_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_13),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_12),
.B(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_16),
.Y(n_33)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_41),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_24),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_0),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_43),
.Y(n_49)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_37),
.B1(n_36),
.B2(n_43),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_44),
.A2(n_52),
.B1(n_54),
.B2(n_58),
.Y(n_75)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_32),
.B1(n_23),
.B2(n_19),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_34),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_53),
.A2(n_21),
.B1(n_25),
.B2(n_27),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_32),
.B1(n_20),
.B2(n_23),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_56),
.Y(n_69)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_61),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_32),
.B1(n_20),
.B2(n_23),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_29),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_60),
.B(n_29),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_21),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_35),
.A2(n_32),
.B1(n_31),
.B2(n_30),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_31),
.B1(n_22),
.B2(n_11),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_72),
.B(n_73),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_27),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_18),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_52),
.B1(n_66),
.B2(n_44),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_77),
.A2(n_83),
.B1(n_86),
.B2(n_88),
.Y(n_107)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_80),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_79),
.Y(n_95)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_49),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_81),
.B(n_84),
.Y(n_109)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_25),
.B1(n_30),
.B2(n_24),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_54),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_42),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_18),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_25),
.B1(n_30),
.B2(n_24),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_87),
.A2(n_46),
.B1(n_18),
.B2(n_64),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_63),
.A2(n_40),
.B1(n_27),
.B2(n_22),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_28),
.B(n_17),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_50),
.B1(n_51),
.B2(n_48),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_94),
.A2(n_106),
.B1(n_74),
.B2(n_90),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_96),
.B(n_101),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_56),
.C(n_42),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_99),
.C(n_114),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_69),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_102),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_71),
.A2(n_84),
.B(n_85),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_71),
.A2(n_28),
.B(n_47),
.C(n_35),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_111),
.Y(n_121)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_103),
.Y(n_132)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_77),
.A2(n_42),
.B1(n_62),
.B2(n_46),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_108),
.A2(n_113),
.B1(n_78),
.B2(n_82),
.Y(n_124)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_110),
.Y(n_131)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_42),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_18),
.B(n_79),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_75),
.A2(n_42),
.B1(n_62),
.B2(n_35),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_67),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_116),
.Y(n_135)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_67),
.Y(n_117)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_118),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_101),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_124),
.A2(n_126),
.B1(n_130),
.B2(n_133),
.Y(n_157)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_127),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_113),
.A2(n_72),
.B1(n_70),
.B2(n_93),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_129),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_70),
.B1(n_93),
.B2(n_90),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_92),
.C(n_79),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_137),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_92),
.C(n_79),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_142),
.B(n_100),
.Y(n_147)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_139),
.B(n_111),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_99),
.B(n_79),
.C(n_74),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_117),
.Y(n_167)
);

OR2x6_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_74),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_144),
.B(n_119),
.Y(n_169)
);

OA21x2_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_18),
.B(n_17),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g144 ( 
.A(n_112),
.B(n_17),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_94),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_146),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_147),
.A2(n_169),
.B(n_141),
.Y(n_189)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_149),
.Y(n_181)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_126),
.Y(n_151)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_152),
.B(n_159),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_145),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_154),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_98),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_160),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_136),
.C(n_123),
.Y(n_173)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_116),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_125),
.B(n_100),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_163),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_145),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_162),
.Y(n_187)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_165),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_135),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_140),
.Y(n_185)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_168),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_143),
.B(n_107),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_172),
.Y(n_192)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_194),
.C(n_198),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_166),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_175),
.B(n_184),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_156),
.B(n_143),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_182),
.B(n_191),
.Y(n_202)
);

OA22x2_ASAP7_75t_L g183 ( 
.A1(n_150),
.A2(n_141),
.B1(n_144),
.B2(n_142),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_183),
.A2(n_106),
.B1(n_120),
.B2(n_124),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_160),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_189),
.Y(n_200)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_190),
.Y(n_222)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_193),
.B(n_161),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_153),
.B(n_138),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_152),
.A2(n_141),
.B(n_144),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_196),
.A2(n_169),
.B1(n_164),
.B2(n_141),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_143),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_197),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_153),
.B(n_167),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_199),
.B(n_177),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_183),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_220),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_176),
.A2(n_157),
.B1(n_163),
.B2(n_150),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_204),
.A2(n_206),
.B1(n_213),
.B2(n_214),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_183),
.A2(n_176),
.B1(n_141),
.B2(n_151),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_205),
.A2(n_186),
.B1(n_193),
.B2(n_190),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_179),
.A2(n_157),
.B1(n_149),
.B2(n_147),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_208),
.Y(n_242)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_192),
.A2(n_170),
.B1(n_172),
.B2(n_133),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_209),
.A2(n_197),
.B1(n_182),
.B2(n_178),
.Y(n_229)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_211),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_148),
.Y(n_212)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_179),
.A2(n_120),
.B1(n_162),
.B2(n_154),
.Y(n_214)
);

AND2x2_ASAP7_75t_SL g215 ( 
.A(n_183),
.B(n_158),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_SL g241 ( 
.A(n_215),
.B(n_95),
.C(n_131),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_158),
.C(n_119),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_173),
.C(n_196),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_191),
.B(n_139),
.Y(n_218)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_192),
.A2(n_128),
.B1(n_107),
.B2(n_142),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_219),
.A2(n_221),
.B1(n_181),
.B2(n_187),
.Y(n_237)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_183),
.A2(n_110),
.B1(n_102),
.B2(n_103),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_180),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_223),
.B(n_180),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_227),
.A2(n_222),
.B(n_212),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_194),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_228),
.B(n_234),
.Y(n_262)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_230),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_209),
.A2(n_178),
.B1(n_177),
.B2(n_189),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_239),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_233),
.A2(n_237),
.B(n_241),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_185),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_223),
.B(n_195),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_235),
.B(n_244),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_240),
.C(n_215),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_205),
.A2(n_188),
.B1(n_187),
.B2(n_175),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_195),
.C(n_95),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_171),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_217),
.Y(n_248)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_208),
.Y(n_245)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

NAND4xp25_ASAP7_75t_SL g246 ( 
.A(n_242),
.B(n_132),
.C(n_105),
.D(n_131),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_2),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_250),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_253),
.C(n_236),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_225),
.A2(n_202),
.B(n_215),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_251),
.A2(n_256),
.B(n_1),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_203),
.C(n_220),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_207),
.Y(n_255)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_255),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_226),
.A2(n_203),
.B(n_199),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_238),
.B(n_219),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_257),
.B(n_234),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_237),
.A2(n_221),
.B1(n_213),
.B2(n_105),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_258),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_0),
.Y(n_261)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_261),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_0),
.Y(n_263)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_263),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_271),
.C(n_262),
.Y(n_287)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_246),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_269),
.A2(n_276),
.B(n_277),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g270 ( 
.A(n_247),
.B(n_233),
.CI(n_231),
.CON(n_270),
.SN(n_270)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_272),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_228),
.C(n_243),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_259),
.B(n_8),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_274),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_275),
.A2(n_261),
.B1(n_250),
.B2(n_260),
.Y(n_284)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_254),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_279),
.Y(n_282)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_245),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_265),
.A2(n_260),
.B1(n_252),
.B2(n_256),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_280),
.B(n_284),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_276),
.B(n_263),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_283),
.A2(n_267),
.B(n_10),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_247),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_286),
.A2(n_288),
.B(n_293),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_271),
.Y(n_295)
);

NAND2x1p5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_251),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_264),
.A2(n_249),
.B1(n_262),
.B2(n_248),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_273),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_9),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_292),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_9),
.Y(n_292)
);

NAND2xp33_ASAP7_75t_L g293 ( 
.A(n_270),
.B(n_8),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_303),
.Y(n_307)
);

AO21x1_ASAP7_75t_L g306 ( 
.A1(n_297),
.A2(n_291),
.B(n_290),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_285),
.B(n_266),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_298),
.B(n_302),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_301),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_3),
.Y(n_301)
);

INVx6_ASAP7_75t_L g302 ( 
.A(n_288),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_3),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_289),
.A2(n_15),
.B(n_14),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_292),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_311),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_302),
.Y(n_308)
);

AO221x1_ASAP7_75t_L g318 ( 
.A1(n_308),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.C(n_11),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_309),
.B(n_296),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_287),
.Y(n_310)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_310),
.Y(n_313)
);

BUFx24_ASAP7_75t_SL g311 ( 
.A(n_299),
.Y(n_311)
);

A2O1A1O1Ixp25_ASAP7_75t_L g319 ( 
.A1(n_315),
.A2(n_318),
.B(n_305),
.C(n_15),
.D(n_5),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_294),
.Y(n_316)
);

AOI321xp33_ASAP7_75t_L g320 ( 
.A1(n_316),
.A2(n_317),
.A3(n_3),
.B1(n_4),
.B2(n_6),
.C(n_7),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_307),
.A2(n_297),
.B(n_4),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_319),
.A2(n_320),
.B(n_313),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_321),
.A2(n_314),
.B(n_6),
.Y(n_322)
);

AOI221xp5_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.C(n_293),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_4),
.Y(n_324)
);


endmodule