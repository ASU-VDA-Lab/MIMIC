module fake_jpeg_7692_n_276 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_276);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_276;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx8_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_37),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_40),
.B(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_22),
.B(n_9),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_24),
.Y(n_54)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_46),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_26),
.C(n_22),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_47),
.Y(n_66)
);

OR2x4_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_29),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_63),
.Y(n_75)
);

INVx5_ASAP7_75t_SL g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_59),
.Y(n_69)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_54),
.B(n_34),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_28),
.B1(n_27),
.B2(n_32),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_57),
.B1(n_17),
.B2(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_27),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_23),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_28),
.B1(n_33),
.B2(n_32),
.Y(n_57)
);

INVx5_ASAP7_75t_SL g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_60),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_17),
.B1(n_33),
.B2(n_32),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_17),
.B1(n_33),
.B2(n_42),
.Y(n_67)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_39),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_34),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_65),
.B(n_79),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_67),
.A2(n_19),
.B1(n_39),
.B2(n_60),
.Y(n_111)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_72),
.A2(n_75),
.B1(n_92),
.B2(n_39),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_31),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_74),
.Y(n_119)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_78),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_31),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_54),
.B(n_20),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_80),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_87),
.Y(n_125)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_82),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_48),
.A2(n_26),
.B1(n_23),
.B2(n_20),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_44),
.Y(n_86)
);

NAND3xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_0),
.C(n_1),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_25),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_49),
.Y(n_88)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_93),
.Y(n_105)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_53),
.Y(n_91)
);

NOR3xp33_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_94),
.C(n_101),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_48),
.A2(n_25),
.B1(n_24),
.B2(n_40),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_35),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_53),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_53),
.A2(n_40),
.B1(n_37),
.B2(n_30),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_97),
.A2(n_59),
.B1(n_37),
.B2(n_29),
.Y(n_107)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_29),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_108),
.B1(n_82),
.B2(n_99),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_86),
.A2(n_59),
.B1(n_29),
.B2(n_19),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_29),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_114),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_111),
.A2(n_116),
.B1(n_126),
.B2(n_97),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_112),
.B(n_13),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_70),
.B(n_19),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_0),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_117),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_116),
.A2(n_14),
.B(n_1),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_70),
.B(n_0),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_86),
.B(n_93),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_39),
.Y(n_158)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_130),
.B(n_131),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_104),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_132),
.B(n_135),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_74),
.B1(n_76),
.B2(n_67),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_138),
.B1(n_141),
.B2(n_150),
.Y(n_163)
);

MAJx2_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_75),
.C(n_81),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_149),
.C(n_119),
.Y(n_164)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_137),
.Y(n_172)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_84),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_139),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_127),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_140),
.A2(n_143),
.B1(n_148),
.B2(n_153),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_128),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_142),
.Y(n_162)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_145),
.A2(n_151),
.B(n_154),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_126),
.A2(n_75),
.B(n_69),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_147),
.A2(n_124),
.B(n_66),
.Y(n_182)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_98),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_115),
.A2(n_94),
.B1(n_91),
.B2(n_80),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_117),
.A2(n_83),
.B1(n_96),
.B2(n_84),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_152),
.A2(n_157),
.B1(n_128),
.B2(n_122),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_127),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_113),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_155),
.B(n_2),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_113),
.A2(n_0),
.B(n_39),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_156),
.A2(n_109),
.B(n_106),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_108),
.A2(n_83),
.B1(n_95),
.B2(n_90),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_149),
.Y(n_178)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_160),
.B(n_166),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_178),
.C(n_179),
.Y(n_191)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_171),
.B(n_146),
.Y(n_194)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_173),
.Y(n_199)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_176),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_151),
.A2(n_109),
.B(n_129),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_181),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_156),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_130),
.B(n_129),
.Y(n_177)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_122),
.C(n_118),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_180),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_137),
.A2(n_124),
.B(n_118),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_66),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_135),
.B(n_3),
.Y(n_183)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_138),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_3),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_185),
.A2(n_141),
.B1(n_145),
.B2(n_147),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_197),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_160),
.A2(n_136),
.B1(n_134),
.B2(n_146),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_155),
.B1(n_143),
.B2(n_124),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_194),
.B(n_206),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_173),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_120),
.C(n_77),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_181),
.C(n_159),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_163),
.A2(n_68),
.B1(n_120),
.B2(n_100),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_198),
.A2(n_183),
.B1(n_170),
.B2(n_68),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_200),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_172),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_180),
.A2(n_176),
.B1(n_166),
.B2(n_184),
.Y(n_202)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_202),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_168),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_163),
.A2(n_68),
.B1(n_120),
.B2(n_77),
.Y(n_207)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_207),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_182),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_211),
.C(n_212),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_203),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_210),
.B(n_215),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_178),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_179),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_218),
.Y(n_234)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_217),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_172),
.C(n_159),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_219),
.A2(n_198),
.B(n_192),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_162),
.Y(n_221)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_221),
.Y(n_231)
);

MAJx2_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_171),
.C(n_175),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_222),
.A2(n_195),
.B1(n_167),
.B2(n_207),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_162),
.Y(n_223)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_225),
.A2(n_202),
.B1(n_161),
.B2(n_200),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_187),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_235),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_210),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_4),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_213),
.A2(n_201),
.B(n_189),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_232),
.A2(n_237),
.B(n_212),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_188),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_218),
.C(n_220),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_219),
.A2(n_198),
.B(n_205),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_197),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_239),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_249)
);

FAx1_ASAP7_75t_L g240 ( 
.A(n_239),
.B(n_220),
.CI(n_216),
.CON(n_240),
.SN(n_240)
);

AO22x1_ASAP7_75t_L g251 ( 
.A1(n_240),
.A2(n_243),
.B1(n_235),
.B2(n_237),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_249),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_177),
.Y(n_242)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_242),
.Y(n_253)
);

OAI21xp33_ASAP7_75t_L g243 ( 
.A1(n_226),
.A2(n_208),
.B(n_219),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_234),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_233),
.A2(n_214),
.B1(n_224),
.B2(n_222),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_250),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_247),
.A2(n_248),
.B(n_6),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_4),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_251),
.A2(n_240),
.B1(n_244),
.B2(n_229),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_257),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_227),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_255),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_236),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_240),
.C(n_244),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_251),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_258),
.Y(n_267)
);

NOR2xp67_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_243),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_263),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_264),
.B(n_254),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_259),
.A2(n_253),
.B(n_229),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_268),
.C(n_6),
.Y(n_271)
);

AOI322xp5_ASAP7_75t_L g270 ( 
.A1(n_267),
.A2(n_254),
.A3(n_259),
.B1(n_261),
.B2(n_258),
.C1(n_12),
.C2(n_13),
.Y(n_270)
);

INVxp33_ASAP7_75t_L g269 ( 
.A(n_266),
.Y(n_269)
);

AOI322xp5_ASAP7_75t_L g272 ( 
.A1(n_269),
.A2(n_270),
.A3(n_271),
.B1(n_16),
.B2(n_10),
.C1(n_11),
.C2(n_12),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_272),
.B(n_273),
.Y(n_274)
);

AOI322xp5_ASAP7_75t_L g273 ( 
.A1(n_269),
.A2(n_8),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_15),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_274),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_8),
.C(n_15),
.Y(n_276)
);


endmodule