module real_aes_8383_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_712;
wire n_183;
wire n_312;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_0), .B(n_105), .C(n_106), .Y(n_104) );
INVx1_ASAP7_75t_L g121 ( .A(n_0), .Y(n_121) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_1), .A2(n_145), .B(n_150), .C(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g257 ( .A(n_2), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_3), .A2(n_140), .B(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_4), .B(n_217), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_5), .Y(n_123) );
AOI21xp33_ASAP7_75t_L g218 ( .A1(n_6), .A2(n_140), .B(n_219), .Y(n_218) );
AND2x6_ASAP7_75t_L g145 ( .A(n_7), .B(n_146), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_8), .A2(n_139), .B(n_147), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_9), .B(n_103), .Y(n_102) );
NOR2xp33_ASAP7_75t_L g122 ( .A(n_9), .B(n_40), .Y(n_122) );
INVx1_ASAP7_75t_L g551 ( .A(n_10), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_11), .B(n_189), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_12), .B(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g224 ( .A(n_13), .Y(n_224) );
INVx1_ASAP7_75t_L g137 ( .A(n_14), .Y(n_137) );
INVx1_ASAP7_75t_L g157 ( .A(n_15), .Y(n_157) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_16), .A2(n_158), .B(n_172), .C(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_17), .B(n_217), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_18), .B(n_174), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_19), .B(n_140), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_20), .B(n_475), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_21), .A2(n_205), .B(n_231), .C(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_22), .B(n_217), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_23), .B(n_189), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g153 ( .A1(n_24), .A2(n_154), .B(n_156), .C(n_158), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_25), .B(n_189), .Y(n_448) );
CKINVDCx16_ASAP7_75t_R g479 ( .A(n_26), .Y(n_479) );
INVx1_ASAP7_75t_L g447 ( .A(n_27), .Y(n_447) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_28), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_29), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_30), .B(n_189), .Y(n_258) );
INVx1_ASAP7_75t_L g472 ( .A(n_31), .Y(n_472) );
INVx1_ASAP7_75t_L g236 ( .A(n_32), .Y(n_236) );
INVx2_ASAP7_75t_L g143 ( .A(n_33), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_34), .Y(n_504) );
A2O1A1Ixp33_ASAP7_75t_L g459 ( .A1(n_35), .A2(n_205), .B(n_225), .C(n_460), .Y(n_459) );
INVxp67_ASAP7_75t_L g473 ( .A(n_36), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g168 ( .A1(n_37), .A2(n_145), .B(n_150), .C(n_169), .Y(n_168) );
A2O1A1Ixp33_ASAP7_75t_L g445 ( .A1(n_38), .A2(n_150), .B(n_446), .C(n_451), .Y(n_445) );
CKINVDCx14_ASAP7_75t_R g458 ( .A(n_39), .Y(n_458) );
INVx1_ASAP7_75t_L g103 ( .A(n_40), .Y(n_103) );
INVx1_ASAP7_75t_L g234 ( .A(n_41), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g549 ( .A1(n_42), .A2(n_176), .B(n_222), .C(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_43), .B(n_189), .Y(n_188) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_44), .A2(n_435), .B1(n_704), .B2(n_713), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_44), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_45), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_46), .Y(n_469) );
INVx1_ASAP7_75t_L g517 ( .A(n_47), .Y(n_517) );
CKINVDCx16_ASAP7_75t_R g237 ( .A(n_48), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_49), .B(n_140), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g230 ( .A1(n_50), .A2(n_150), .B1(n_231), .B2(n_233), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_51), .Y(n_180) );
CKINVDCx16_ASAP7_75t_R g254 ( .A(n_52), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_53), .A2(n_222), .B(n_223), .C(n_225), .Y(n_221) );
CKINVDCx14_ASAP7_75t_R g548 ( .A(n_54), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g193 ( .A(n_55), .Y(n_193) );
INVx1_ASAP7_75t_L g220 ( .A(n_56), .Y(n_220) );
INVx1_ASAP7_75t_L g146 ( .A(n_57), .Y(n_146) );
INVx1_ASAP7_75t_L g136 ( .A(n_58), .Y(n_136) );
INVx1_ASAP7_75t_SL g461 ( .A(n_59), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_60), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_61), .B(n_217), .Y(n_521) );
INVx1_ASAP7_75t_L g482 ( .A(n_62), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_SL g244 ( .A1(n_63), .A2(n_174), .B(n_225), .C(n_245), .Y(n_244) );
INVxp67_ASAP7_75t_L g246 ( .A(n_64), .Y(n_246) );
AOI222xp33_ASAP7_75t_SL g124 ( .A1(n_65), .A2(n_67), .B1(n_125), .B2(n_699), .C1(n_700), .C2(n_707), .Y(n_124) );
INVx1_ASAP7_75t_L g108 ( .A(n_66), .Y(n_108) );
INVx1_ASAP7_75t_L g699 ( .A(n_67), .Y(n_699) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_68), .A2(n_140), .B(n_547), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_69), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_70), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_71), .A2(n_140), .B(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g184 ( .A(n_72), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_73), .A2(n_139), .B(n_468), .Y(n_467) );
CKINVDCx16_ASAP7_75t_R g444 ( .A(n_74), .Y(n_444) );
INVx1_ASAP7_75t_L g509 ( .A(n_75), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_76), .A2(n_100), .B1(n_109), .B2(n_716), .Y(n_99) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_77), .A2(n_145), .B(n_150), .C(n_187), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_78), .A2(n_140), .B(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g512 ( .A(n_79), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_80), .B(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g134 ( .A(n_81), .Y(n_134) );
INVx1_ASAP7_75t_L g501 ( .A(n_82), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_83), .B(n_174), .Y(n_173) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_84), .A2(n_145), .B(n_150), .C(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g105 ( .A(n_85), .Y(n_105) );
OR2x2_ASAP7_75t_L g118 ( .A(n_85), .B(n_119), .Y(n_118) );
OR2x2_ASAP7_75t_L g698 ( .A(n_85), .B(n_120), .Y(n_698) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_86), .A2(n_150), .B(n_481), .C(n_485), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_87), .B(n_133), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g261 ( .A(n_88), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_89), .A2(n_145), .B(n_150), .C(n_202), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_90), .Y(n_210) );
INVx1_ASAP7_75t_L g243 ( .A(n_91), .Y(n_243) );
CKINVDCx16_ASAP7_75t_R g148 ( .A(n_92), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_93), .B(n_171), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_94), .B(n_162), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_95), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_96), .B(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_97), .A2(n_140), .B(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g520 ( .A(n_98), .Y(n_520) );
INVx1_ASAP7_75t_L g716 ( .A(n_100), .Y(n_716) );
INVx1_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
OR2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_104), .Y(n_101) );
OR2x2_ASAP7_75t_L g434 ( .A(n_105), .B(n_120), .Y(n_434) );
NOR2x2_ASAP7_75t_L g709 ( .A(n_105), .B(n_119), .Y(n_709) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
AOI22x1_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_124), .B1(n_710), .B2(n_711), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_111), .B(n_115), .Y(n_110) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_SL g710 ( .A(n_113), .Y(n_710) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_115), .A2(n_712), .B(n_714), .Y(n_711) );
NOR2xp33_ASAP7_75t_SL g115 ( .A(n_116), .B(n_123), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_SL g715 ( .A(n_118), .Y(n_715) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_126), .A2(n_434), .B1(n_435), .B2(n_698), .Y(n_125) );
INVx2_ASAP7_75t_SL g701 ( .A(n_126), .Y(n_701) );
OR4x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_330), .C(n_389), .D(n_416), .Y(n_126) );
NAND3xp33_ASAP7_75t_SL g127 ( .A(n_128), .B(n_272), .C(n_297), .Y(n_127) );
O2A1O1Ixp33_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_195), .B(n_215), .C(n_248), .Y(n_128) );
AOI211xp5_ASAP7_75t_SL g420 ( .A1(n_129), .A2(n_421), .B(n_423), .C(n_426), .Y(n_420) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_164), .Y(n_129) );
INVx1_ASAP7_75t_L g295 ( .A(n_130), .Y(n_295) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OR2x2_ASAP7_75t_L g270 ( .A(n_131), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g302 ( .A(n_131), .Y(n_302) );
AND2x2_ASAP7_75t_L g357 ( .A(n_131), .B(n_326), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_131), .B(n_213), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_131), .B(n_214), .Y(n_415) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g276 ( .A(n_132), .Y(n_276) );
AND2x2_ASAP7_75t_L g319 ( .A(n_132), .B(n_182), .Y(n_319) );
AND2x2_ASAP7_75t_L g337 ( .A(n_132), .B(n_214), .Y(n_337) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_138), .B(n_161), .Y(n_132) );
INVx1_ASAP7_75t_L g194 ( .A(n_133), .Y(n_194) );
INVx2_ASAP7_75t_L g199 ( .A(n_133), .Y(n_199) );
O2A1O1Ixp33_ASAP7_75t_L g443 ( .A1(n_133), .A2(n_185), .B(n_444), .C(n_445), .Y(n_443) );
OA21x2_ASAP7_75t_L g545 ( .A1(n_133), .A2(n_546), .B(n_552), .Y(n_545) );
AND2x2_ASAP7_75t_SL g133 ( .A(n_134), .B(n_135), .Y(n_133) );
AND2x2_ASAP7_75t_L g163 ( .A(n_134), .B(n_135), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
BUFx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_145), .Y(n_140) );
NAND2x1p5_ASAP7_75t_L g185 ( .A(n_141), .B(n_145), .Y(n_185) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
INVx1_ASAP7_75t_L g450 ( .A(n_142), .Y(n_450) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g151 ( .A(n_143), .Y(n_151) );
INVx1_ASAP7_75t_L g232 ( .A(n_143), .Y(n_232) );
INVx1_ASAP7_75t_L g152 ( .A(n_144), .Y(n_152) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_144), .Y(n_155) );
INVx3_ASAP7_75t_L g172 ( .A(n_144), .Y(n_172) );
INVx1_ASAP7_75t_L g174 ( .A(n_144), .Y(n_174) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_144), .Y(n_189) );
INVx4_ASAP7_75t_SL g160 ( .A(n_145), .Y(n_160) );
BUFx3_ASAP7_75t_L g451 ( .A(n_145), .Y(n_451) );
O2A1O1Ixp33_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_149), .B(n_153), .C(n_160), .Y(n_147) );
O2A1O1Ixp33_ASAP7_75t_L g219 ( .A1(n_149), .A2(n_160), .B(n_220), .C(n_221), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g242 ( .A1(n_149), .A2(n_160), .B(n_243), .C(n_244), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g457 ( .A1(n_149), .A2(n_160), .B(n_458), .C(n_459), .Y(n_457) );
O2A1O1Ixp33_ASAP7_75t_SL g468 ( .A1(n_149), .A2(n_160), .B(n_469), .C(n_470), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_SL g508 ( .A1(n_149), .A2(n_160), .B(n_509), .C(n_510), .Y(n_508) );
O2A1O1Ixp33_ASAP7_75t_SL g516 ( .A1(n_149), .A2(n_160), .B(n_517), .C(n_518), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_SL g547 ( .A1(n_149), .A2(n_160), .B(n_548), .C(n_549), .Y(n_547) );
INVx5_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x6_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
BUFx3_ASAP7_75t_L g159 ( .A(n_151), .Y(n_159) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_151), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_154), .B(n_157), .Y(n_156) );
OAI22xp33_ASAP7_75t_L g471 ( .A1(n_154), .A2(n_171), .B1(n_472), .B2(n_473), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_154), .B(n_512), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_154), .B(n_520), .Y(n_519) );
INVx4_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
OAI22xp5_ASAP7_75t_SL g233 ( .A1(n_155), .A2(n_234), .B1(n_235), .B2(n_236), .Y(n_233) );
INVx2_ASAP7_75t_L g235 ( .A(n_155), .Y(n_235) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g176 ( .A(n_159), .Y(n_176) );
OAI22xp33_ASAP7_75t_L g229 ( .A1(n_160), .A2(n_185), .B1(n_230), .B2(n_237), .Y(n_229) );
INVx1_ASAP7_75t_L g485 ( .A(n_160), .Y(n_485) );
INVx4_ASAP7_75t_L g181 ( .A(n_162), .Y(n_181) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_162), .A2(n_241), .B(n_247), .Y(n_240) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_162), .Y(n_455) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g178 ( .A(n_163), .Y(n_178) );
INVx4_ASAP7_75t_L g269 ( .A(n_164), .Y(n_269) );
OAI21xp5_ASAP7_75t_L g324 ( .A1(n_164), .A2(n_325), .B(n_327), .Y(n_324) );
AND2x2_ASAP7_75t_L g405 ( .A(n_164), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g164 ( .A(n_165), .B(n_182), .Y(n_164) );
INVx1_ASAP7_75t_L g212 ( .A(n_165), .Y(n_212) );
AND2x2_ASAP7_75t_L g274 ( .A(n_165), .B(n_214), .Y(n_274) );
OR2x2_ASAP7_75t_L g303 ( .A(n_165), .B(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g317 ( .A(n_165), .Y(n_317) );
INVx3_ASAP7_75t_L g326 ( .A(n_165), .Y(n_326) );
AND2x2_ASAP7_75t_L g336 ( .A(n_165), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g369 ( .A(n_165), .B(n_275), .Y(n_369) );
AND2x2_ASAP7_75t_L g393 ( .A(n_165), .B(n_349), .Y(n_393) );
OR2x6_ASAP7_75t_L g165 ( .A(n_166), .B(n_179), .Y(n_165) );
AOI21xp5_ASAP7_75t_SL g166 ( .A1(n_167), .A2(n_168), .B(n_177), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_173), .B(n_175), .Y(n_169) );
O2A1O1Ixp33_ASAP7_75t_L g256 ( .A1(n_171), .A2(n_257), .B(n_258), .C(n_259), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_L g446 ( .A1(n_171), .A2(n_447), .B(n_448), .C(n_449), .Y(n_446) );
INVx5_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_172), .B(n_224), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_172), .B(n_246), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_172), .B(n_551), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_175), .A2(n_188), .B(n_190), .Y(n_187) );
O2A1O1Ixp33_ASAP7_75t_L g481 ( .A1(n_175), .A2(n_482), .B(n_483), .C(n_484), .Y(n_481) );
O2A1O1Ixp5_ASAP7_75t_L g500 ( .A1(n_175), .A2(n_483), .B(n_501), .C(n_502), .Y(n_500) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g191 ( .A(n_177), .Y(n_191) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_178), .A2(n_229), .B(n_238), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_178), .B(n_239), .Y(n_238) );
AO21x2_ASAP7_75t_L g252 ( .A1(n_178), .A2(n_253), .B(n_260), .Y(n_252) );
NOR2xp33_ASAP7_75t_SL g179 ( .A(n_180), .B(n_181), .Y(n_179) );
INVx3_ASAP7_75t_L g217 ( .A(n_181), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_181), .B(n_453), .Y(n_452) );
AO21x2_ASAP7_75t_L g477 ( .A1(n_181), .A2(n_478), .B(n_486), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_181), .B(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g214 ( .A(n_182), .Y(n_214) );
AND2x2_ASAP7_75t_L g429 ( .A(n_182), .B(n_271), .Y(n_429) );
AO21x2_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_191), .B(n_192), .Y(n_182) );
OAI21xp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_186), .Y(n_183) );
OAI21xp5_ASAP7_75t_L g253 ( .A1(n_185), .A2(n_254), .B(n_255), .Y(n_253) );
OAI21xp5_ASAP7_75t_L g478 ( .A1(n_185), .A2(n_479), .B(n_480), .Y(n_478) );
OAI21xp5_ASAP7_75t_L g497 ( .A1(n_185), .A2(n_498), .B(n_499), .Y(n_497) );
INVx4_ASAP7_75t_L g205 ( .A(n_189), .Y(n_205) );
INVx2_ASAP7_75t_L g222 ( .A(n_189), .Y(n_222) );
INVx1_ASAP7_75t_L g466 ( .A(n_191), .Y(n_466) );
AO21x2_ASAP7_75t_L g490 ( .A1(n_191), .A2(n_491), .B(n_492), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_194), .B(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_194), .B(n_261), .Y(n_260) );
AO21x2_ASAP7_75t_L g496 ( .A1(n_194), .A2(n_497), .B(n_503), .Y(n_496) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_211), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_197), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g349 ( .A(n_197), .B(n_337), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_197), .B(n_326), .Y(n_411) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g271 ( .A(n_198), .Y(n_271) );
AND2x2_ASAP7_75t_L g275 ( .A(n_198), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g316 ( .A(n_198), .B(n_317), .Y(n_316) );
AO21x2_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_209), .Y(n_198) );
INVx1_ASAP7_75t_L g475 ( .A(n_199), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_199), .B(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_201), .B(n_208), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_206), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_205), .B(n_461), .Y(n_460) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx3_ASAP7_75t_L g225 ( .A(n_207), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_211), .B(n_312), .Y(n_334) );
INVx1_ASAP7_75t_L g373 ( .A(n_211), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_211), .B(n_300), .Y(n_417) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
AND2x2_ASAP7_75t_L g280 ( .A(n_212), .B(n_275), .Y(n_280) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_214), .B(n_271), .Y(n_304) );
INVx1_ASAP7_75t_L g383 ( .A(n_214), .Y(n_383) );
AOI322xp5_ASAP7_75t_L g407 ( .A1(n_215), .A2(n_322), .A3(n_382), .B1(n_408), .B2(n_410), .C1(n_412), .C2(n_414), .Y(n_407) );
AND2x2_ASAP7_75t_SL g215 ( .A(n_216), .B(n_227), .Y(n_215) );
AND2x2_ASAP7_75t_L g262 ( .A(n_216), .B(n_240), .Y(n_262) );
INVx1_ASAP7_75t_SL g265 ( .A(n_216), .Y(n_265) );
AND2x2_ASAP7_75t_L g267 ( .A(n_216), .B(n_228), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_216), .B(n_284), .Y(n_290) );
INVx2_ASAP7_75t_L g309 ( .A(n_216), .Y(n_309) );
AND2x2_ASAP7_75t_L g322 ( .A(n_216), .B(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g360 ( .A(n_216), .B(n_284), .Y(n_360) );
BUFx2_ASAP7_75t_L g377 ( .A(n_216), .Y(n_377) );
AND2x2_ASAP7_75t_L g391 ( .A(n_216), .B(n_251), .Y(n_391) );
OA21x2_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B(n_226), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_227), .B(n_279), .Y(n_306) );
AND2x2_ASAP7_75t_L g433 ( .A(n_227), .B(n_309), .Y(n_433) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_240), .Y(n_227) );
OR2x2_ASAP7_75t_L g278 ( .A(n_228), .B(n_279), .Y(n_278) );
INVx3_ASAP7_75t_L g284 ( .A(n_228), .Y(n_284) );
AND2x2_ASAP7_75t_L g329 ( .A(n_228), .B(n_252), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_228), .B(n_377), .Y(n_376) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_228), .Y(n_413) );
INVx2_ASAP7_75t_L g259 ( .A(n_231), .Y(n_259) );
INVx3_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g483 ( .A(n_235), .Y(n_483) );
AND2x2_ASAP7_75t_L g264 ( .A(n_240), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g286 ( .A(n_240), .Y(n_286) );
BUFx2_ASAP7_75t_L g292 ( .A(n_240), .Y(n_292) );
AND2x2_ASAP7_75t_L g311 ( .A(n_240), .B(n_284), .Y(n_311) );
INVx3_ASAP7_75t_L g323 ( .A(n_240), .Y(n_323) );
OR2x2_ASAP7_75t_L g333 ( .A(n_240), .B(n_284), .Y(n_333) );
AOI31xp33_ASAP7_75t_SL g248 ( .A1(n_249), .A2(n_263), .A3(n_266), .B(n_268), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_262), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_250), .B(n_285), .Y(n_296) );
OR2x2_ASAP7_75t_L g320 ( .A(n_250), .B(n_290), .Y(n_320) );
INVx1_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_251), .B(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g341 ( .A(n_251), .B(n_333), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_251), .B(n_323), .Y(n_351) );
AND2x2_ASAP7_75t_L g358 ( .A(n_251), .B(n_359), .Y(n_358) );
NAND2x1_ASAP7_75t_L g386 ( .A(n_251), .B(n_322), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_251), .B(n_377), .Y(n_387) );
AND2x2_ASAP7_75t_L g399 ( .A(n_251), .B(n_284), .Y(n_399) );
INVx3_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx3_ASAP7_75t_L g279 ( .A(n_252), .Y(n_279) );
INVx1_ASAP7_75t_L g345 ( .A(n_262), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_262), .B(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_264), .B(n_340), .Y(n_374) );
AND2x4_ASAP7_75t_L g285 ( .A(n_265), .B(n_286), .Y(n_285) );
CKINVDCx16_ASAP7_75t_R g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx2_ASAP7_75t_L g364 ( .A(n_270), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_270), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g312 ( .A(n_271), .B(n_302), .Y(n_312) );
AND2x2_ASAP7_75t_L g406 ( .A(n_271), .B(n_276), .Y(n_406) );
INVx1_ASAP7_75t_L g431 ( .A(n_271), .Y(n_431) );
AOI221xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_277), .B1(n_280), .B2(n_281), .C(n_287), .Y(n_272) );
CKINVDCx14_ASAP7_75t_R g293 ( .A(n_273), .Y(n_293) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_274), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_277), .B(n_328), .Y(n_347) );
INVx3_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g396 ( .A(n_278), .B(n_292), .Y(n_396) );
AND2x2_ASAP7_75t_L g310 ( .A(n_279), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g340 ( .A(n_279), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_279), .B(n_323), .Y(n_368) );
NOR3xp33_ASAP7_75t_L g410 ( .A(n_279), .B(n_380), .C(n_411), .Y(n_410) );
AOI211xp5_ASAP7_75t_SL g343 ( .A1(n_280), .A2(n_344), .B(n_346), .C(n_354), .Y(n_343) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OAI22xp33_ASAP7_75t_L g332 ( .A1(n_282), .A2(n_333), .B1(n_334), .B2(n_335), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_283), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_283), .B(n_367), .Y(n_366) );
BUFx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g425 ( .A(n_285), .B(n_399), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_293), .B1(n_294), .B2(n_296), .Y(n_287) );
NOR2xp33_ASAP7_75t_SL g288 ( .A(n_289), .B(n_291), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_291), .B(n_340), .Y(n_371) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_294), .A2(n_386), .B1(n_417), .B2(n_424), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_305), .B1(n_307), .B2(n_312), .C(n_313), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_303), .Y(n_299) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVxp67_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OAI221xp5_ASAP7_75t_L g313 ( .A1(n_303), .A2(n_314), .B1(n_320), .B2(n_321), .C(n_324), .Y(n_313) );
INVx1_ASAP7_75t_L g356 ( .A(n_304), .Y(n_356) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx1_ASAP7_75t_SL g328 ( .A(n_309), .Y(n_328) );
OR2x2_ASAP7_75t_L g401 ( .A(n_309), .B(n_333), .Y(n_401) );
AND2x2_ASAP7_75t_L g403 ( .A(n_309), .B(n_311), .Y(n_403) );
INVx1_ASAP7_75t_L g342 ( .A(n_312), .Y(n_342) );
OR2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_318), .Y(n_314) );
AOI21xp33_ASAP7_75t_SL g372 ( .A1(n_315), .A2(n_373), .B(n_374), .Y(n_372) );
OR2x2_ASAP7_75t_L g379 ( .A(n_315), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g353 ( .A(n_316), .B(n_337), .Y(n_353) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp33_ASAP7_75t_SL g370 ( .A(n_321), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_322), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_323), .B(n_359), .Y(n_422) );
O2A1O1Ixp33_ASAP7_75t_L g338 ( .A1(n_326), .A2(n_339), .B(n_341), .C(n_342), .Y(n_338) );
NAND2x1_ASAP7_75t_SL g363 ( .A(n_326), .B(n_364), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_327), .A2(n_376), .B1(n_378), .B2(n_381), .Y(n_375) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_329), .B(n_419), .Y(n_418) );
NAND5xp2_ASAP7_75t_L g330 ( .A(n_331), .B(n_343), .C(n_361), .D(n_375), .E(n_384), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_332), .B(n_338), .Y(n_331) );
INVx1_ASAP7_75t_L g388 ( .A(n_334), .Y(n_388) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_336), .A2(n_355), .B1(n_395), .B2(n_397), .C(n_400), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_337), .B(n_431), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_340), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_340), .B(n_406), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_348), .B1(n_350), .B2(n_352), .Y(n_346) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_358), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
AND2x2_ASAP7_75t_L g428 ( .A(n_357), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AOI221xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_365), .B1(n_369), .B2(n_370), .C(n_372), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g412 ( .A(n_367), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g419 ( .A(n_377), .Y(n_419) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI21xp5_ASAP7_75t_SL g384 ( .A1(n_385), .A2(n_387), .B(n_388), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
OAI211xp5_ASAP7_75t_SL g389 ( .A1(n_390), .A2(n_392), .B(n_394), .C(n_407), .Y(n_389) );
INVx1_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
A2O1A1Ixp33_ASAP7_75t_L g416 ( .A1(n_392), .A2(n_417), .B(n_418), .C(n_420), .Y(n_416) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_396), .B(n_398), .Y(n_397) );
AOI21xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B(n_404), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AOI21xp33_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_430), .B(n_432), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g703 ( .A(n_434), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_435), .Y(n_704) );
OR3x1_ASAP7_75t_L g435 ( .A(n_436), .B(n_609), .C(n_656), .Y(n_435) );
NAND3xp33_ASAP7_75t_SL g436 ( .A(n_437), .B(n_555), .C(n_580), .Y(n_436) );
AOI221xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_495), .B1(n_522), .B2(n_525), .C(n_533), .Y(n_437) );
OAI21xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_463), .B(n_488), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_440), .B(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_440), .B(n_538), .Y(n_653) );
AND2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_454), .Y(n_440) );
AND2x2_ASAP7_75t_L g524 ( .A(n_441), .B(n_494), .Y(n_524) );
AND2x2_ASAP7_75t_L g573 ( .A(n_441), .B(n_493), .Y(n_573) );
AND2x2_ASAP7_75t_L g594 ( .A(n_441), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g599 ( .A(n_441), .B(n_566), .Y(n_599) );
OR2x2_ASAP7_75t_L g607 ( .A(n_441), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g679 ( .A(n_441), .B(n_476), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_441), .B(n_628), .Y(n_693) );
INVx3_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g539 ( .A(n_442), .B(n_454), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_442), .B(n_476), .Y(n_540) );
AND2x4_ASAP7_75t_L g561 ( .A(n_442), .B(n_494), .Y(n_561) );
AND2x2_ASAP7_75t_L g591 ( .A(n_442), .B(n_465), .Y(n_591) );
AND2x2_ASAP7_75t_L g600 ( .A(n_442), .B(n_590), .Y(n_600) );
AND2x2_ASAP7_75t_L g616 ( .A(n_442), .B(n_477), .Y(n_616) );
OR2x2_ASAP7_75t_L g625 ( .A(n_442), .B(n_608), .Y(n_625) );
AND2x2_ASAP7_75t_L g631 ( .A(n_442), .B(n_566), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_442), .B(n_637), .Y(n_636) );
OR2x2_ASAP7_75t_L g645 ( .A(n_442), .B(n_490), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_442), .B(n_535), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_442), .B(n_595), .Y(n_684) );
OR2x6_ASAP7_75t_L g442 ( .A(n_443), .B(n_452), .Y(n_442) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_450), .B(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g494 ( .A(n_454), .Y(n_494) );
AND2x2_ASAP7_75t_L g590 ( .A(n_454), .B(n_476), .Y(n_590) );
AND2x2_ASAP7_75t_L g595 ( .A(n_454), .B(n_477), .Y(n_595) );
INVx1_ASAP7_75t_L g651 ( .A(n_454), .Y(n_651) );
OA21x2_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_456), .B(n_462), .Y(n_454) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_455), .A2(n_507), .B(n_513), .Y(n_506) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_455), .A2(n_515), .B(n_521), .Y(n_514) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g560 ( .A(n_464), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_476), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_465), .B(n_524), .Y(n_523) );
BUFx3_ASAP7_75t_L g538 ( .A(n_465), .Y(n_538) );
OR2x2_ASAP7_75t_L g608 ( .A(n_465), .B(n_476), .Y(n_608) );
OR2x2_ASAP7_75t_L g669 ( .A(n_465), .B(n_576), .Y(n_669) );
OA21x2_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_467), .B(n_474), .Y(n_465) );
INVx1_ASAP7_75t_L g491 ( .A(n_467), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_474), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_476), .B(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g628 ( .A(n_476), .B(n_490), .Y(n_628) );
INVx2_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
BUFx2_ASAP7_75t_L g567 ( .A(n_477), .Y(n_567) );
INVx1_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
AOI221xp5_ASAP7_75t_L g672 ( .A1(n_489), .A2(n_673), .B1(n_677), .B2(n_680), .C(n_681), .Y(n_672) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_493), .Y(n_489) );
INVx1_ASAP7_75t_SL g536 ( .A(n_490), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_490), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g667 ( .A(n_490), .B(n_524), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_493), .B(n_538), .Y(n_659) );
AND2x2_ASAP7_75t_L g566 ( .A(n_494), .B(n_567), .Y(n_566) );
INVx1_ASAP7_75t_SL g570 ( .A(n_495), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_495), .B(n_576), .Y(n_606) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_505), .Y(n_495) );
AND2x2_ASAP7_75t_L g532 ( .A(n_496), .B(n_506), .Y(n_532) );
INVx4_ASAP7_75t_L g544 ( .A(n_496), .Y(n_544) );
BUFx3_ASAP7_75t_L g586 ( .A(n_496), .Y(n_586) );
AND3x2_ASAP7_75t_L g601 ( .A(n_496), .B(n_602), .C(n_603), .Y(n_601) );
AND2x2_ASAP7_75t_L g683 ( .A(n_505), .B(n_597), .Y(n_683) );
AND2x2_ASAP7_75t_L g691 ( .A(n_505), .B(n_576), .Y(n_691) );
INVx1_ASAP7_75t_SL g696 ( .A(n_505), .Y(n_696) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_514), .Y(n_505) );
INVx1_ASAP7_75t_SL g554 ( .A(n_506), .Y(n_554) );
AND2x2_ASAP7_75t_L g577 ( .A(n_506), .B(n_544), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_506), .B(n_528), .Y(n_579) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_506), .Y(n_619) );
OR2x2_ASAP7_75t_L g624 ( .A(n_506), .B(n_544), .Y(n_624) );
INVx2_ASAP7_75t_L g530 ( .A(n_514), .Y(n_530) );
AND2x2_ASAP7_75t_L g564 ( .A(n_514), .B(n_545), .Y(n_564) );
OR2x2_ASAP7_75t_L g584 ( .A(n_514), .B(n_545), .Y(n_584) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_514), .Y(n_604) );
INVx1_ASAP7_75t_SL g522 ( .A(n_523), .Y(n_522) );
AOI21xp33_ASAP7_75t_L g654 ( .A1(n_523), .A2(n_563), .B(n_655), .Y(n_654) );
AOI322xp5_ASAP7_75t_L g690 ( .A1(n_525), .A2(n_535), .A3(n_561), .B1(n_691), .B2(n_692), .C1(n_694), .C2(n_697), .Y(n_690) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_531), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_527), .B(n_634), .Y(n_633) );
INVx1_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_528), .B(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g553 ( .A(n_529), .B(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g621 ( .A(n_530), .B(n_544), .Y(n_621) );
AND2x2_ASAP7_75t_L g688 ( .A(n_530), .B(n_545), .Y(n_688) );
INVx1_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g629 ( .A(n_532), .B(n_583), .Y(n_629) );
AOI31xp33_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_537), .A3(n_540), .B(n_541), .Y(n_533) );
AND2x2_ASAP7_75t_L g588 ( .A(n_535), .B(n_566), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_535), .B(n_558), .Y(n_670) );
AND2x2_ASAP7_75t_L g689 ( .A(n_535), .B(n_594), .Y(n_689) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_538), .B(n_566), .Y(n_578) );
NAND2x1p5_ASAP7_75t_L g612 ( .A(n_538), .B(n_595), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g615 ( .A(n_538), .B(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_538), .B(n_679), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_539), .B(n_595), .Y(n_627) );
INVx1_ASAP7_75t_L g671 ( .A(n_539), .Y(n_671) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_553), .Y(n_542) );
INVxp67_ASAP7_75t_L g623 ( .A(n_543), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_544), .B(n_554), .Y(n_559) );
INVx1_ASAP7_75t_L g665 ( .A(n_544), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_544), .B(n_642), .Y(n_676) );
BUFx3_ASAP7_75t_L g576 ( .A(n_545), .Y(n_576) );
AND2x2_ASAP7_75t_L g602 ( .A(n_545), .B(n_554), .Y(n_602) );
INVx2_ASAP7_75t_L g642 ( .A(n_545), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g674 ( .A(n_553), .B(n_675), .Y(n_674) );
AOI211xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_560), .B(n_562), .C(n_571), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AOI21xp33_ASAP7_75t_L g605 ( .A1(n_557), .A2(n_606), .B(n_607), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_558), .B(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_558), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OR2x2_ASAP7_75t_L g638 ( .A(n_559), .B(n_584), .Y(n_638) );
INVx3_ASAP7_75t_L g569 ( .A(n_561), .Y(n_569) );
OAI22xp5_ASAP7_75t_SL g562 ( .A1(n_563), .A2(n_565), .B1(n_568), .B2(n_570), .Y(n_562) );
OAI21xp5_ASAP7_75t_SL g587 ( .A1(n_564), .A2(n_588), .B(n_589), .Y(n_587) );
AND2x2_ASAP7_75t_L g613 ( .A(n_564), .B(n_577), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_564), .B(n_665), .Y(n_664) );
INVxp67_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g568 ( .A(n_567), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g637 ( .A(n_567), .Y(n_637) );
OAI21xp5_ASAP7_75t_SL g581 ( .A1(n_568), .A2(n_582), .B(n_587), .Y(n_581) );
OAI22xp33_ASAP7_75t_SL g571 ( .A1(n_572), .A2(n_574), .B1(n_578), .B2(n_579), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_573), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
INVx1_ASAP7_75t_L g597 ( .A(n_576), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_576), .B(n_619), .Y(n_618) );
NOR3xp33_ASAP7_75t_L g580 ( .A(n_581), .B(n_592), .C(n_605), .Y(n_580) );
OAI22xp5_ASAP7_75t_SL g647 ( .A1(n_582), .A2(n_648), .B1(n_652), .B2(n_653), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_583), .B(n_585), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g652 ( .A(n_584), .B(n_585), .Y(n_652) );
AND2x2_ASAP7_75t_L g660 ( .A(n_585), .B(n_641), .Y(n_660) );
CKINVDCx16_ASAP7_75t_R g585 ( .A(n_586), .Y(n_585) );
O2A1O1Ixp33_ASAP7_75t_SL g668 ( .A1(n_586), .A2(n_669), .B(n_670), .C(n_671), .Y(n_668) );
OR2x2_ASAP7_75t_L g695 ( .A(n_586), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
OAI21xp33_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_596), .B(n_598), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
O2A1O1Ixp33_ASAP7_75t_L g630 ( .A1(n_594), .A2(n_631), .B(n_632), .C(n_635), .Y(n_630) );
OAI21xp33_ASAP7_75t_SL g598 ( .A1(n_599), .A2(n_600), .B(n_601), .Y(n_598) );
AND2x2_ASAP7_75t_L g663 ( .A(n_602), .B(n_621), .Y(n_663) );
INVxp67_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g641 ( .A(n_604), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g646 ( .A(n_606), .Y(n_646) );
NAND3xp33_ASAP7_75t_SL g609 ( .A(n_610), .B(n_630), .C(n_643), .Y(n_609) );
AOI211xp5_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_613), .B(n_614), .C(n_622), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_617), .Y(n_614) );
INVx1_ASAP7_75t_L g680 ( .A(n_617), .Y(n_680) );
OR2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
INVx1_ASAP7_75t_L g640 ( .A(n_619), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_619), .B(n_688), .Y(n_687) );
INVxp67_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
A2O1A1Ixp33_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_624), .B(n_625), .C(n_626), .Y(n_622) );
INVx2_ASAP7_75t_SL g634 ( .A(n_624), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_625), .A2(n_636), .B1(n_638), .B2(n_639), .Y(n_635) );
OAI21xp33_ASAP7_75t_SL g626 ( .A1(n_627), .A2(n_628), .B(n_629), .Y(n_626) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
AOI211xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_646), .B(n_647), .C(n_654), .Y(n_643) );
INVx1_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
INVxp33_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g697 ( .A(n_651), .Y(n_697) );
NAND4xp25_ASAP7_75t_L g656 ( .A(n_657), .B(n_672), .C(n_685), .D(n_690), .Y(n_656) );
AOI211xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_660), .B(n_661), .C(n_668), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AOI21xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_664), .B(n_666), .Y(n_661) );
AOI21xp33_ASAP7_75t_L g681 ( .A1(n_662), .A2(n_682), .B(n_684), .Y(n_681) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_669), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_689), .Y(n_685) );
INVxp67_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g706 ( .A(n_698), .Y(n_706) );
OAI22xp5_ASAP7_75t_SL g700 ( .A1(n_701), .A2(n_702), .B1(n_704), .B2(n_705), .Y(n_700) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVx3_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
endmodule