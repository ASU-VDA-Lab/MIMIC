module fake_netlist_6_4204_n_191 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_191);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_191;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_63;
wire n_39;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_184;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_160;
wire n_90;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_188;
wire n_102;
wire n_186;
wire n_87;
wire n_189;
wire n_32;
wire n_66;
wire n_130;
wire n_85;
wire n_78;
wire n_84;
wire n_99;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_181;
wire n_76;
wire n_36;
wire n_182;
wire n_124;
wire n_55;
wire n_126;
wire n_94;
wire n_97;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_190;
wire n_123;
wire n_136;
wire n_72;
wire n_187;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_35;
wire n_183;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_171;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx2_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_30),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_23),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_28),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

BUFx8_ASAP7_75t_SL g54 ( 
.A(n_52),
.Y(n_54)
);

INVxp33_ASAP7_75t_SL g55 ( 
.A(n_51),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

AO22x2_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_53),
.B(n_2),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_3),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_4),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx8_ASAP7_75t_SL g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_37),
.B(n_5),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g73 ( 
.A(n_37),
.B(n_5),
.C(n_6),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

CKINVDCx11_ASAP7_75t_R g76 ( 
.A(n_54),
.Y(n_76)
);

AOI211xp5_ASAP7_75t_L g77 ( 
.A1(n_59),
.A2(n_46),
.B(n_40),
.C(n_49),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_71),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_55),
.B(n_33),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_49),
.B1(n_48),
.B2(n_46),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_33),
.Y(n_82)
);

AND2x6_ASAP7_75t_SL g83 ( 
.A(n_61),
.B(n_48),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

AND2x4_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_45),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

BUFx8_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_62),
.B(n_43),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_44),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

OAI21x1_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_66),
.B(n_63),
.Y(n_93)
);

AO21x2_ASAP7_75t_L g94 ( 
.A1(n_91),
.A2(n_66),
.B(n_41),
.Y(n_94)
);

AO31x2_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_68),
.A3(n_65),
.B(n_64),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_68),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_53),
.B1(n_72),
.B2(n_73),
.Y(n_97)
);

OAI21x1_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_63),
.B(n_65),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_68),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_76),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_73),
.B(n_65),
.C(n_64),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_72),
.B1(n_57),
.B2(n_50),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_77),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_101),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_88),
.Y(n_106)
);

AOI21x1_ASAP7_75t_SL g107 ( 
.A1(n_96),
.A2(n_87),
.B(n_57),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_SL g108 ( 
.A1(n_103),
.A2(n_45),
.B(n_88),
.C(n_41),
.Y(n_108)
);

BUFx8_ASAP7_75t_SL g109 ( 
.A(n_92),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_79),
.Y(n_111)
);

AND2x4_ASAP7_75t_SL g112 ( 
.A(n_106),
.B(n_100),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_94),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_92),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

NOR2x1_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_111),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_111),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_114),
.Y(n_123)
);

AND2x4_ASAP7_75t_SL g124 ( 
.A(n_120),
.B(n_117),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_113),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_104),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_104),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_111),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_105),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_112),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_112),
.Y(n_134)
);

AOI222xp33_ASAP7_75t_L g135 ( 
.A1(n_129),
.A2(n_97),
.B1(n_89),
.B2(n_90),
.C1(n_103),
.C2(n_57),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_104),
.Y(n_136)
);

AOI31xp33_ASAP7_75t_L g137 ( 
.A1(n_130),
.A2(n_105),
.A3(n_102),
.B(n_70),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_133),
.A2(n_108),
.B(n_118),
.C(n_47),
.Y(n_139)
);

XOR2x2_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_83),
.Y(n_140)
);

OAI322xp33_ASAP7_75t_L g141 ( 
.A1(n_127),
.A2(n_74),
.A3(n_69),
.B1(n_47),
.B2(n_56),
.C1(n_58),
.C2(n_60),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_134),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_125),
.Y(n_143)
);

AOI211xp5_ASAP7_75t_SL g144 ( 
.A1(n_137),
.A2(n_128),
.B(n_134),
.C(n_126),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_89),
.B1(n_126),
.B2(n_128),
.Y(n_145)
);

AOI211xp5_ASAP7_75t_L g146 ( 
.A1(n_141),
.A2(n_108),
.B(n_74),
.C(n_58),
.Y(n_146)
);

AOI221xp5_ASAP7_75t_L g147 ( 
.A1(n_141),
.A2(n_57),
.B1(n_86),
.B2(n_85),
.C(n_81),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_93),
.B(n_131),
.Y(n_149)
);

AOI32xp33_ASAP7_75t_L g150 ( 
.A1(n_136),
.A2(n_57),
.A3(n_39),
.B1(n_89),
.B2(n_60),
.Y(n_150)
);

AOI221xp5_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_86),
.B1(n_85),
.B2(n_43),
.C(n_83),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_136),
.A2(n_132),
.B1(n_124),
.B2(n_138),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_151),
.B(n_140),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_94),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_89),
.C(n_87),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_144),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_124),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_146),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_64),
.Y(n_162)
);

NAND4xp75_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_147),
.C(n_150),
.D(n_9),
.Y(n_163)
);

AND2x4_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_17),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_15),
.Y(n_165)
);

AND2x4_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_24),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_93),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

AOI221xp5_ASAP7_75t_L g169 ( 
.A1(n_160),
.A2(n_87),
.B1(n_8),
.B2(n_11),
.C(n_12),
.Y(n_169)
);

NAND3xp33_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_87),
.C(n_100),
.Y(n_170)
);

OAI221xp5_ASAP7_75t_SL g171 ( 
.A1(n_169),
.A2(n_159),
.B1(n_154),
.B2(n_11),
.C(n_13),
.Y(n_171)
);

OAI221xp5_ASAP7_75t_SL g172 ( 
.A1(n_165),
.A2(n_7),
.B1(n_8),
.B2(n_14),
.C(n_109),
.Y(n_172)
);

AND2x4_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_14),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_SL g174 ( 
.A(n_170),
.B(n_118),
.C(n_117),
.Y(n_174)
);

OAI221xp5_ASAP7_75t_L g175 ( 
.A1(n_162),
.A2(n_75),
.B1(n_78),
.B2(n_84),
.C(n_100),
.Y(n_175)
);

NAND3xp33_ASAP7_75t_SL g176 ( 
.A(n_167),
.B(n_26),
.C(n_29),
.Y(n_176)
);

OAI211xp5_ASAP7_75t_SL g177 ( 
.A1(n_163),
.A2(n_84),
.B(n_96),
.C(n_99),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_168),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_173),
.B(n_164),
.Y(n_179)
);

NAND2x1p5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_163),
.Y(n_180)
);

AO21x1_ASAP7_75t_L g181 ( 
.A1(n_172),
.A2(n_93),
.B(n_98),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_31),
.Y(n_182)
);

OA21x2_ASAP7_75t_L g183 ( 
.A1(n_175),
.A2(n_98),
.B(n_84),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_176),
.A2(n_75),
.B1(n_100),
.B2(n_110),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_180),
.A2(n_100),
.B1(n_110),
.B2(n_107),
.Y(n_185)
);

AO22x2_ASAP7_75t_L g186 ( 
.A1(n_184),
.A2(n_107),
.B1(n_110),
.B2(n_99),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_181),
.A2(n_95),
.B1(n_110),
.B2(n_178),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_179),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_187),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_186),
.A2(n_182),
.B(n_183),
.Y(n_190)
);

AOI221xp5_ASAP7_75t_L g191 ( 
.A1(n_189),
.A2(n_95),
.B1(n_185),
.B2(n_186),
.C(n_190),
.Y(n_191)
);


endmodule