module real_aes_6664_n_383 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_383);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_383;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_635;
wire n_792;
wire n_673;
wire n_386;
wire n_503;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_991;
wire n_667;
wire n_1114;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_841;
wire n_718;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_852;
wire n_766;
wire n_1113;
wire n_974;
wire n_919;
wire n_1089;
wire n_857;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_1123;
wire n_952;
wire n_429;
wire n_1110;
wire n_1137;
wire n_448;
wire n_545;
wire n_556;
wire n_752;
wire n_593;
wire n_460;
wire n_937;
wire n_989;
wire n_773;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_537;
wire n_884;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_1146;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_1147;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_677;
wire n_958;
wire n_1021;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1140;
wire n_1099;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_1108;
wire n_966;
wire n_1160;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_1078;
wire n_994;
wire n_1072;
wire n_384;
wire n_744;
wire n_938;
wire n_1128;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_951;
wire n_875;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_962;
wire n_693;
wire n_1082;
wire n_468;
wire n_746;
wire n_656;
wire n_532;
wire n_755;
wire n_1025;
wire n_1148;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_874;
wire n_796;
wire n_1152;
wire n_801;
wire n_1126;
wire n_529;
wire n_1115;
wire n_455;
wire n_960;
wire n_504;
wire n_725;
wire n_671;
wire n_1084;
wire n_973;
wire n_1081;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1121;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_936;
wire n_610;
wire n_581;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_1135;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_1100;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_449;
wire n_754;
wire n_607;
wire n_417;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_1142;
wire n_1141;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_1149;
wire n_405;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_617;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1103;
wire n_1031;
wire n_1037;
wire n_1131;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1154;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_1145;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_501;
wire n_488;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_1163;
wire n_945;
wire n_604;
wire n_898;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_713;
wire n_598;
wire n_404;
wire n_735;
wire n_728;
wire n_756;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1105;
wire n_1132;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_1003;
wire n_533;
wire n_1000;
wire n_1028;
wire n_1014;
wire n_727;
wire n_1083;
wire n_397;
wire n_749;
wire n_385;
wire n_663;
wire n_1056;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_915;
wire n_1002;
wire n_1155;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_1043;
wire n_850;
wire n_1136;
wire n_720;
wire n_972;
wire n_1127;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_831;
wire n_487;
wire n_653;
wire n_526;
wire n_928;
wire n_637;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_922;
wire n_520;
wire n_482;
wire n_633;
wire n_926;
wire n_679;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_1130;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_1090;
wire n_1133;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_1162;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_698;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_823;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1150;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_1161;
wire n_1143;
wire n_929;
wire n_686;
wire n_776;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_1159;
wire n_1156;
wire n_829;
wire n_1030;
wire n_1088;
wire n_988;
wire n_1055;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1151;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_968;
wire n_650;
wire n_646;
wire n_710;
wire n_743;
wire n_393;
wire n_1040;
wire n_703;
wire n_652;
wire n_500;
wire n_601;
wire n_1097;
wire n_661;
wire n_463;
wire n_1076;
wire n_396;
wire n_804;
wire n_1101;
wire n_447;
wire n_1102;
wire n_603;
wire n_403;
wire n_854;
wire n_1119;
wire n_424;
wire n_1039;
wire n_802;
wire n_868;
wire n_877;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_1144;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_1153;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_0), .A2(n_197), .B1(n_680), .B2(n_681), .Y(n_679) );
INVx1_ASAP7_75t_L g817 ( .A(n_1), .Y(n_817) );
AOI22xp33_ASAP7_75t_SL g1102 ( .A1(n_2), .A2(n_248), .B1(n_617), .B2(n_1103), .Y(n_1102) );
AOI222xp33_ASAP7_75t_L g899 ( .A1(n_3), .A2(n_187), .B1(n_334), .B2(n_471), .C1(n_478), .C2(n_524), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_4), .A2(n_259), .B1(n_537), .B2(n_557), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_5), .A2(n_109), .B1(n_687), .B2(n_700), .Y(n_699) );
AOI221xp5_ASAP7_75t_L g854 ( .A1(n_6), .A2(n_328), .B1(n_455), .B2(n_687), .C(n_855), .Y(n_854) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_7), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_8), .A2(n_83), .B1(n_524), .B2(n_1003), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_9), .A2(n_243), .B1(n_621), .B2(n_922), .Y(n_921) );
AO22x2_ASAP7_75t_L g408 ( .A1(n_10), .A2(n_232), .B1(n_409), .B2(n_410), .Y(n_408) );
INVx1_ASAP7_75t_L g1120 ( .A(n_10), .Y(n_1120) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_11), .A2(n_179), .B1(n_452), .B2(n_872), .Y(n_892) );
AOI22xp33_ASAP7_75t_SL g574 ( .A1(n_12), .A2(n_357), .B1(n_520), .B2(n_575), .Y(n_574) );
CKINVDCx20_ASAP7_75t_R g932 ( .A(n_13), .Y(n_932) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_14), .A2(n_168), .B1(n_456), .B2(n_561), .Y(n_652) );
CKINVDCx20_ASAP7_75t_R g608 ( .A(n_15), .Y(n_608) );
CKINVDCx20_ASAP7_75t_R g627 ( .A(n_16), .Y(n_627) );
INVx1_ASAP7_75t_L g764 ( .A(n_17), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_18), .A2(n_200), .B1(n_579), .B2(n_735), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_19), .A2(n_255), .B1(n_447), .B2(n_456), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_20), .A2(n_113), .B1(n_687), .B2(n_709), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_21), .A2(n_322), .B1(n_708), .B2(n_709), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g977 ( .A(n_22), .Y(n_977) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_23), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_24), .A2(n_323), .B1(n_429), .B2(n_436), .Y(n_428) );
AOI22xp33_ASAP7_75t_SL g737 ( .A1(n_25), .A2(n_312), .B1(n_455), .B2(n_540), .Y(n_737) );
AOI222xp33_ASAP7_75t_L g883 ( .A1(n_26), .A2(n_70), .B1(n_285), .B2(n_520), .C1(n_610), .C2(n_884), .Y(n_883) );
AOI22xp5_ASAP7_75t_SL g559 ( .A1(n_27), .A2(n_253), .B1(n_560), .B2(n_561), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g638 ( .A(n_28), .Y(n_638) );
AOI221xp5_ASAP7_75t_L g859 ( .A1(n_29), .A2(n_40), .B1(n_713), .B2(n_735), .C(n_860), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g1105 ( .A1(n_30), .A2(n_258), .B1(n_452), .B2(n_537), .Y(n_1105) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_31), .A2(n_364), .B1(n_430), .B2(n_654), .Y(n_653) );
CKINVDCx20_ASAP7_75t_R g934 ( .A(n_32), .Y(n_934) );
CKINVDCx20_ASAP7_75t_R g596 ( .A(n_33), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_34), .A2(n_251), .B1(n_535), .B2(n_872), .Y(n_1070) );
AO22x2_ASAP7_75t_L g412 ( .A1(n_35), .A2(n_128), .B1(n_409), .B2(n_413), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_36), .A2(n_182), .B1(n_437), .B2(n_448), .Y(n_1074) );
CKINVDCx20_ASAP7_75t_R g885 ( .A(n_37), .Y(n_885) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_38), .A2(n_664), .B1(n_690), .B2(n_691), .Y(n_663) );
INVx1_ASAP7_75t_L g691 ( .A(n_38), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_39), .A2(n_57), .B1(n_532), .B2(n_535), .Y(n_531) );
AOI22xp33_ASAP7_75t_SL g1073 ( .A1(n_41), .A2(n_64), .B1(n_452), .B2(n_550), .Y(n_1073) );
INVx1_ASAP7_75t_L g795 ( .A(n_42), .Y(n_795) );
AOI22xp5_ASAP7_75t_L g1063 ( .A1(n_43), .A2(n_295), .B1(n_524), .B2(n_1064), .Y(n_1063) );
AOI22xp5_ASAP7_75t_L g824 ( .A1(n_44), .A2(n_65), .B1(n_454), .B2(n_656), .Y(n_824) );
INVx1_ASAP7_75t_L g1138 ( .A(n_45), .Y(n_1138) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_46), .A2(n_175), .B1(n_545), .B2(n_872), .Y(n_1023) );
INVx1_ASAP7_75t_L g857 ( .A(n_47), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_48), .A2(n_308), .B1(n_617), .B2(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g1019 ( .A(n_49), .Y(n_1019) );
AOI22xp5_ASAP7_75t_L g793 ( .A1(n_50), .A2(n_220), .B1(n_485), .B2(n_572), .Y(n_793) );
AOI222xp33_ASAP7_75t_L g863 ( .A1(n_51), .A2(n_146), .B1(n_155), .B2(n_478), .C1(n_483), .C2(n_518), .Y(n_863) );
AOI22xp5_ASAP7_75t_SL g556 ( .A1(n_52), .A2(n_318), .B1(n_557), .B2(n_558), .Y(n_556) );
AOI222xp33_ASAP7_75t_L g715 ( .A1(n_53), .A2(n_303), .B1(n_321), .B2(n_523), .C1(n_594), .C2(n_716), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g900 ( .A(n_54), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_55), .A2(n_129), .B1(n_532), .B2(n_913), .Y(n_912) );
AOI22xp5_ASAP7_75t_SL g823 ( .A1(n_56), .A2(n_231), .B1(n_456), .B2(n_558), .Y(n_823) );
INVx1_ASAP7_75t_L g773 ( .A(n_58), .Y(n_773) );
CKINVDCx20_ASAP7_75t_R g605 ( .A(n_59), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_60), .A2(n_185), .B1(n_436), .B2(n_549), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_61), .A2(n_329), .B1(n_731), .B2(n_878), .Y(n_877) );
CKINVDCx16_ASAP7_75t_R g591 ( .A(n_62), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_63), .A2(n_306), .B1(n_601), .B2(n_675), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_66), .B(n_523), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g1075 ( .A(n_67), .Y(n_1075) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_68), .A2(n_362), .B1(n_421), .B2(n_683), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_69), .A2(n_277), .B1(n_603), .B2(n_727), .Y(n_771) );
AOI22xp5_ASAP7_75t_L g1020 ( .A1(n_71), .A2(n_98), .B1(n_524), .B2(n_731), .Y(n_1020) );
AOI22xp5_ASAP7_75t_L g1123 ( .A1(n_72), .A2(n_1124), .B1(n_1148), .B2(n_1149), .Y(n_1123) );
CKINVDCx20_ASAP7_75t_R g1148 ( .A(n_72), .Y(n_1148) );
INVx1_ASAP7_75t_L g815 ( .A(n_73), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_74), .A2(n_158), .B1(n_543), .B2(n_547), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g805 ( .A(n_75), .B(n_565), .Y(n_805) );
CKINVDCx20_ASAP7_75t_R g668 ( .A(n_76), .Y(n_668) );
AOI22xp33_ASAP7_75t_SL g1099 ( .A1(n_77), .A2(n_211), .B1(n_922), .B2(n_1100), .Y(n_1099) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_78), .A2(n_99), .B1(n_779), .B2(n_919), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_79), .A2(n_228), .B1(n_579), .B2(n_582), .Y(n_578) );
CKINVDCx20_ASAP7_75t_R g650 ( .A(n_80), .Y(n_650) );
INVx1_ASAP7_75t_L g1091 ( .A(n_81), .Y(n_1091) );
INVx1_ASAP7_75t_L g769 ( .A(n_82), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_84), .A2(n_102), .B1(n_537), .B2(n_538), .Y(n_536) );
AOI22xp5_ASAP7_75t_SL g826 ( .A1(n_85), .A2(n_103), .B1(n_535), .B2(n_749), .Y(n_826) );
INVx1_ASAP7_75t_L g1146 ( .A(n_86), .Y(n_1146) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_87), .A2(n_161), .B1(n_543), .B2(n_960), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_88), .A2(n_167), .B1(n_621), .B2(n_984), .Y(n_1134) );
AO22x2_ASAP7_75t_L g418 ( .A1(n_89), .A2(n_266), .B1(n_409), .B2(n_410), .Y(n_418) );
INVx1_ASAP7_75t_L g1117 ( .A(n_89), .Y(n_1117) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_90), .A2(n_276), .B1(n_430), .B2(n_437), .Y(n_882) );
AOI22xp33_ASAP7_75t_SL g1098 ( .A1(n_91), .A2(n_92), .B1(n_779), .B2(n_919), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_93), .A2(n_353), .B1(n_610), .B2(n_645), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_94), .A2(n_350), .B1(n_545), .B2(n_660), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_95), .A2(n_369), .B1(n_549), .B2(n_551), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_96), .A2(n_299), .B1(n_598), .B2(n_673), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_97), .A2(n_225), .B1(n_523), .B2(n_670), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_100), .A2(n_314), .B1(n_656), .B2(n_658), .Y(n_655) );
OA22x2_ASAP7_75t_L g695 ( .A1(n_101), .A2(n_696), .B1(n_697), .B2(n_717), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_101), .Y(n_696) );
AOI22xp33_ASAP7_75t_SL g827 ( .A1(n_104), .A2(n_213), .B1(n_565), .B2(n_617), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g1024 ( .A1(n_105), .A2(n_122), .B1(n_535), .B2(n_881), .Y(n_1024) );
INVx1_ASAP7_75t_L g1137 ( .A(n_106), .Y(n_1137) );
AOI22xp33_ASAP7_75t_SL g1066 ( .A1(n_107), .A2(n_115), .B1(n_575), .B2(n_716), .Y(n_1066) );
INVx1_ASAP7_75t_L g820 ( .A(n_108), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_110), .A2(n_244), .B1(n_984), .B2(n_986), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_111), .A2(n_137), .B1(n_683), .B2(n_684), .Y(n_682) );
INVx1_ASAP7_75t_L g1127 ( .A(n_112), .Y(n_1127) );
AOI22xp33_ASAP7_75t_SL g732 ( .A1(n_114), .A2(n_222), .B1(n_713), .B2(n_733), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_116), .Y(n_569) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_117), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_118), .B(n_1015), .Y(n_1014) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_119), .Y(n_796) );
AOI22xp5_ASAP7_75t_L g782 ( .A1(n_120), .A2(n_250), .B1(n_430), .B2(n_783), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g947 ( .A(n_121), .Y(n_947) );
AOI22xp5_ASAP7_75t_L g1005 ( .A1(n_123), .A2(n_284), .B1(n_558), .B2(n_874), .Y(n_1005) );
INVx1_ASAP7_75t_L g1132 ( .A(n_124), .Y(n_1132) );
CKINVDCx20_ASAP7_75t_R g978 ( .A(n_125), .Y(n_978) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_126), .Y(n_745) );
INVx1_ASAP7_75t_L g1001 ( .A(n_127), .Y(n_1001) );
INVx1_ASAP7_75t_L g1121 ( .A(n_128), .Y(n_1121) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_130), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g917 ( .A(n_131), .Y(n_917) );
AOI22xp5_ASAP7_75t_L g999 ( .A1(n_132), .A2(n_208), .B1(n_576), .B2(n_607), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_133), .A2(n_141), .B1(n_617), .B2(n_986), .Y(n_1027) );
CKINVDCx20_ASAP7_75t_R g419 ( .A(n_134), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g1082 ( .A1(n_135), .A2(n_1083), .B1(n_1084), .B2(n_1085), .Y(n_1082) );
INVx1_ASAP7_75t_L g1083 ( .A(n_135), .Y(n_1083) );
CKINVDCx20_ASAP7_75t_R g951 ( .A(n_136), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_138), .A2(n_212), .B1(n_913), .B2(n_956), .Y(n_955) );
CKINVDCx20_ASAP7_75t_R g830 ( .A(n_139), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_140), .A2(n_267), .B1(n_601), .B2(n_675), .Y(n_928) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_142), .Y(n_460) );
AOI211xp5_ASAP7_75t_L g593 ( .A1(n_143), .A2(n_594), .B(n_595), .C(n_604), .Y(n_593) );
INVx1_ASAP7_75t_L g1009 ( .A(n_144), .Y(n_1009) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_145), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g946 ( .A(n_147), .Y(n_946) );
CKINVDCx20_ASAP7_75t_R g911 ( .A(n_148), .Y(n_911) );
INVx1_ASAP7_75t_L g1028 ( .A(n_149), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_150), .A2(n_338), .B1(n_615), .B2(n_618), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g1071 ( .A1(n_151), .A2(n_181), .B1(n_778), .B2(n_881), .Y(n_1071) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_152), .A2(n_264), .B1(n_603), .B2(n_727), .Y(n_835) );
AOI22xp33_ASAP7_75t_SL g738 ( .A1(n_153), .A2(n_230), .B1(n_446), .B2(n_660), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_154), .Y(n_747) );
AOI211xp5_ASAP7_75t_L g739 ( .A1(n_156), .A2(n_683), .B(n_740), .C(n_746), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g1017 ( .A1(n_157), .A2(n_360), .B1(n_520), .B2(n_575), .Y(n_1017) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_159), .Y(n_465) );
CKINVDCx16_ASAP7_75t_R g1158 ( .A(n_160), .Y(n_1158) );
AOI22xp5_ASAP7_75t_L g1162 ( .A1(n_160), .A2(n_1124), .B1(n_1149), .B2(n_1158), .Y(n_1162) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_162), .A2(n_194), .B1(n_437), .B2(n_550), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_163), .A2(n_359), .B1(n_600), .B2(n_601), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_164), .A2(n_279), .B1(n_572), .B2(n_600), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_165), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_166), .A2(n_242), .B1(n_621), .B2(n_689), .Y(n_688) );
AND2x6_ASAP7_75t_L g386 ( .A(n_169), .B(n_387), .Y(n_386) );
HB1xp67_ASAP7_75t_L g1114 ( .A(n_169), .Y(n_1114) );
AOI22xp33_ASAP7_75t_L g1130 ( .A1(n_170), .A2(n_310), .B1(n_564), .B2(n_617), .Y(n_1130) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_171), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_172), .Y(n_798) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_173), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_174), .A2(n_265), .B1(n_483), .B2(n_670), .Y(n_975) );
AOI22xp33_ASAP7_75t_SL g1026 ( .A1(n_176), .A2(n_355), .B1(n_540), .B2(n_550), .Y(n_1026) );
AOI22xp5_ASAP7_75t_L g571 ( .A1(n_177), .A2(n_247), .B1(n_524), .B2(n_572), .Y(n_571) );
AO22x1_ASAP7_75t_L g851 ( .A1(n_178), .A2(n_190), .B1(n_852), .B2(n_853), .Y(n_851) );
AOI221xp5_ASAP7_75t_L g850 ( .A1(n_180), .A2(n_337), .B1(n_537), .B2(n_557), .C(n_851), .Y(n_850) );
AOI22xp5_ASAP7_75t_L g1002 ( .A1(n_183), .A2(n_379), .B1(n_484), .B2(n_1003), .Y(n_1002) );
INVx1_ASAP7_75t_L g971 ( .A(n_184), .Y(n_971) );
INVx1_ASAP7_75t_L g1095 ( .A(n_186), .Y(n_1095) );
INVx1_ASAP7_75t_L g1142 ( .A(n_188), .Y(n_1142) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_189), .Y(n_450) );
AOI22xp33_ASAP7_75t_SL g1006 ( .A1(n_191), .A2(n_195), .B1(n_547), .B2(n_986), .Y(n_1006) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_192), .Y(n_526) );
AO22x2_ASAP7_75t_L g416 ( .A1(n_193), .A2(n_254), .B1(n_409), .B2(n_413), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g1118 ( .A(n_193), .B(n_1119), .Y(n_1118) );
CKINVDCx20_ASAP7_75t_R g640 ( .A(n_196), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_198), .A2(n_256), .B1(n_656), .B2(n_778), .Y(n_889) );
AOI22xp33_ASAP7_75t_SL g1007 ( .A1(n_199), .A2(n_348), .B1(n_456), .B2(n_778), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1092 ( .A1(n_201), .A2(n_382), .B1(n_520), .B2(n_727), .Y(n_1092) );
INVx1_ASAP7_75t_L g1088 ( .A(n_202), .Y(n_1088) );
AOI22xp33_ASAP7_75t_SL g777 ( .A1(n_203), .A2(n_336), .B1(n_778), .B2(n_779), .Y(n_777) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_204), .Y(n_728) );
INVx1_ASAP7_75t_L g1094 ( .A(n_205), .Y(n_1094) );
AOI22xp5_ASAP7_75t_SL g563 ( .A1(n_206), .A2(n_280), .B1(n_564), .B2(n_565), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g1046 ( .A(n_207), .Y(n_1046) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_209), .A2(n_245), .B1(n_660), .B2(n_872), .Y(n_871) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_210), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g1055 ( .A1(n_214), .A2(n_343), .B1(n_437), .B2(n_615), .Y(n_1055) );
CKINVDCx20_ASAP7_75t_R g974 ( .A(n_215), .Y(n_974) );
CKINVDCx20_ASAP7_75t_R g1056 ( .A(n_216), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_217), .B(n_897), .Y(n_896) );
AOI22xp33_ASAP7_75t_SL g730 ( .A1(n_218), .A2(n_352), .B1(n_600), .B2(n_731), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g399 ( .A1(n_219), .A2(n_400), .B1(n_500), .B2(n_501), .Y(n_399) );
INVx1_ASAP7_75t_L g500 ( .A(n_219), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g926 ( .A(n_221), .Y(n_926) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_223), .Y(n_516) );
AOI22xp33_ASAP7_75t_SL g1054 ( .A1(n_224), .A2(n_372), .B1(n_558), .B2(n_687), .Y(n_1054) );
CKINVDCx20_ASAP7_75t_R g623 ( .A(n_226), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g846 ( .A1(n_227), .A2(n_847), .B1(n_848), .B2(n_864), .Y(n_846) );
INVx1_ASAP7_75t_L g864 ( .A(n_227), .Y(n_864) );
CKINVDCx20_ASAP7_75t_R g642 ( .A(n_229), .Y(n_642) );
CKINVDCx20_ASAP7_75t_R g927 ( .A(n_233), .Y(n_927) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_234), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_235), .A2(n_246), .B1(n_452), .B2(n_455), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g909 ( .A(n_236), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_237), .A2(n_356), .B1(n_615), .B2(n_618), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_238), .B(n_735), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_239), .A2(n_301), .B1(n_601), .B2(n_675), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_240), .A2(n_367), .B1(n_547), .B2(n_660), .Y(n_893) );
CKINVDCx20_ASAP7_75t_R g583 ( .A(n_241), .Y(n_583) );
AND2x2_ASAP7_75t_L g390 ( .A(n_249), .B(n_391), .Y(n_390) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_252), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_257), .A2(n_272), .B1(n_557), .B2(n_874), .Y(n_873) );
OA22x2_ASAP7_75t_L g758 ( .A1(n_260), .A2(n_759), .B1(n_760), .B2(n_761), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_260), .Y(n_759) );
AOI22xp33_ASAP7_75t_SL g786 ( .A1(n_261), .A2(n_291), .B1(n_551), .B2(n_658), .Y(n_786) );
AOI22xp5_ASAP7_75t_L g903 ( .A1(n_262), .A2(n_904), .B1(n_935), .B2(n_936), .Y(n_903) );
INVx1_ASAP7_75t_L g935 ( .A(n_262), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_263), .A2(n_317), .B1(n_447), .B2(n_881), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_268), .A2(n_316), .B1(n_620), .B2(n_621), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_269), .A2(n_361), .B1(n_779), .B2(n_989), .Y(n_988) );
AOI211xp5_ASAP7_75t_L g383 ( .A1(n_270), .A2(n_384), .B(n_392), .C(n_1122), .Y(n_383) );
INVx1_ASAP7_75t_L g792 ( .A(n_271), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_273), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_274), .A2(n_381), .B1(n_703), .B2(n_705), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_275), .A2(n_349), .B1(n_681), .B2(n_982), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_278), .A2(n_320), .B1(n_673), .B2(n_713), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_281), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_282), .A2(n_332), .B1(n_532), .B2(n_962), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_283), .A2(n_365), .B1(n_598), .B2(n_735), .Y(n_876) );
CKINVDCx20_ASAP7_75t_R g832 ( .A(n_286), .Y(n_832) );
INVx1_ASAP7_75t_L g409 ( .A(n_287), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_287), .Y(n_411) );
INVx1_ASAP7_75t_L g1089 ( .A(n_288), .Y(n_1089) );
INVx1_ASAP7_75t_L g1041 ( .A(n_289), .Y(n_1041) );
INVx1_ASAP7_75t_L g1140 ( .A(n_290), .Y(n_1140) );
AOI22xp5_ASAP7_75t_L g942 ( .A1(n_292), .A2(n_943), .B1(n_963), .B2(n_964), .Y(n_942) );
CKINVDCx20_ASAP7_75t_R g963 ( .A(n_292), .Y(n_963) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_293), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_294), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g807 ( .A(n_296), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g811 ( .A(n_297), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g861 ( .A(n_298), .Y(n_861) );
AOI22xp5_ASAP7_75t_L g1008 ( .A1(n_300), .A2(n_340), .B1(n_618), .B2(n_881), .Y(n_1008) );
INVx1_ASAP7_75t_L g1039 ( .A(n_302), .Y(n_1039) );
INVx1_ASAP7_75t_L g1133 ( .A(n_304), .Y(n_1133) );
CKINVDCx20_ASAP7_75t_R g839 ( .A(n_305), .Y(n_839) );
INVx1_ASAP7_75t_L g972 ( .A(n_307), .Y(n_972) );
CKINVDCx20_ASAP7_75t_R g931 ( .A(n_309), .Y(n_931) );
CKINVDCx20_ASAP7_75t_R g950 ( .A(n_311), .Y(n_950) );
CKINVDCx20_ASAP7_75t_R g647 ( .A(n_313), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_315), .A2(n_341), .B1(n_575), .B2(n_603), .Y(n_898) );
AO22x2_ASAP7_75t_L g634 ( .A1(n_319), .A2(n_635), .B1(n_661), .B2(n_662), .Y(n_634) );
CKINVDCx20_ASAP7_75t_R g662 ( .A(n_319), .Y(n_662) );
INVx1_ASAP7_75t_L g391 ( .A(n_324), .Y(n_391) );
AOI22xp5_ASAP7_75t_SL g967 ( .A1(n_325), .A2(n_968), .B1(n_990), .B2(n_991), .Y(n_967) );
INVx1_ASAP7_75t_L g991 ( .A(n_325), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g1143 ( .A(n_326), .B(n_1144), .Y(n_1143) );
INVx1_ASAP7_75t_L g387 ( .A(n_327), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_330), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g1016 ( .A(n_331), .B(n_897), .Y(n_1016) );
INVx1_ASAP7_75t_L g1147 ( .A(n_333), .Y(n_1147) );
INVx1_ASAP7_75t_L g818 ( .A(n_335), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_339), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g774 ( .A(n_342), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g920 ( .A(n_344), .Y(n_920) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_345), .Y(n_808) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_346), .Y(n_834) );
CKINVDCx20_ASAP7_75t_R g895 ( .A(n_347), .Y(n_895) );
CKINVDCx20_ASAP7_75t_R g1047 ( .A(n_351), .Y(n_1047) );
INVx1_ASAP7_75t_L g629 ( .A(n_354), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_358), .B(n_897), .Y(n_997) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_363), .Y(n_625) );
INVx1_ASAP7_75t_L g766 ( .A(n_366), .Y(n_766) );
INVx1_ASAP7_75t_L g856 ( .A(n_368), .Y(n_856) );
XNOR2xp5_ASAP7_75t_L g719 ( .A(n_370), .B(n_720), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g952 ( .A(n_371), .Y(n_952) );
INVx1_ASAP7_75t_L g1129 ( .A(n_373), .Y(n_1129) );
CKINVDCx20_ASAP7_75t_R g1043 ( .A(n_374), .Y(n_1043) );
OA22x2_ASAP7_75t_L g503 ( .A1(n_375), .A2(n_504), .B1(n_505), .B2(n_552), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_375), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g862 ( .A(n_376), .Y(n_862) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_377), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_378), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g1062 ( .A(n_380), .Y(n_1062) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_388), .Y(n_385) );
HB1xp67_ASAP7_75t_L g1113 ( .A(n_387), .Y(n_1113) );
OAI21xp5_ASAP7_75t_L g1156 ( .A1(n_388), .A2(n_1112), .B(n_1157), .Y(n_1156) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_389), .Y(n_388) );
INVxp67_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_841), .B1(n_1107), .B2(n_1108), .C(n_1109), .Y(n_392) );
INVx1_ASAP7_75t_L g1107 ( .A(n_393), .Y(n_1107) );
XOR2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_754), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_397), .B1(n_585), .B2(n_586), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
XOR2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_502), .Y(n_397) );
BUFx3_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g501 ( .A(n_400), .Y(n_501) );
AND2x2_ASAP7_75t_SL g400 ( .A(n_401), .B(n_458), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_402), .B(n_440), .Y(n_401) );
OAI221xp5_ASAP7_75t_SL g402 ( .A1(n_403), .A2(n_419), .B1(n_420), .B2(n_427), .C(n_428), .Y(n_402) );
INVx3_ASAP7_75t_L g557 ( .A(n_403), .Y(n_557) );
INVx2_ASAP7_75t_SL g709 ( .A(n_403), .Y(n_709) );
INVx4_ASAP7_75t_L g749 ( .A(n_403), .Y(n_749) );
INVx11_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx11_ASAP7_75t_L g546 ( .A(n_404), .Y(n_546) );
AND2x6_ASAP7_75t_L g404 ( .A(n_405), .B(n_414), .Y(n_404) );
AND2x4_ASAP7_75t_L g581 ( .A(n_405), .B(n_449), .Y(n_581) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g463 ( .A(n_406), .B(n_464), .Y(n_463) );
OR2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_412), .Y(n_406) );
AND2x2_ASAP7_75t_L g425 ( .A(n_407), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g435 ( .A(n_407), .B(n_412), .Y(n_435) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g475 ( .A(n_408), .B(n_416), .Y(n_475) );
AND2x2_ASAP7_75t_L g480 ( .A(n_408), .B(n_412), .Y(n_480) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_411), .Y(n_413) );
INVx2_ASAP7_75t_L g426 ( .A(n_412), .Y(n_426) );
INVx1_ASAP7_75t_L g439 ( .A(n_412), .Y(n_439) );
AND2x2_ASAP7_75t_L g443 ( .A(n_414), .B(n_425), .Y(n_443) );
AND2x4_ASAP7_75t_L g454 ( .A(n_414), .B(n_435), .Y(n_454) );
AND2x6_ASAP7_75t_L g479 ( .A(n_414), .B(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_417), .Y(n_414) );
AND2x2_ASAP7_75t_L g449 ( .A(n_415), .B(n_418), .Y(n_449) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_416), .B(n_418), .Y(n_424) );
AND2x2_ASAP7_75t_L g433 ( .A(n_416), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g434 ( .A(n_418), .Y(n_434) );
INVx1_ASAP7_75t_L g474 ( .A(n_418), .Y(n_474) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
HB1xp67_ASAP7_75t_L g853 ( .A(n_421), .Y(n_853) );
BUFx3_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx3_ASAP7_75t_L g535 ( .A(n_422), .Y(n_535) );
BUFx3_ASAP7_75t_L g564 ( .A(n_422), .Y(n_564) );
BUFx2_ASAP7_75t_L g618 ( .A(n_422), .Y(n_618) );
BUFx3_ASAP7_75t_L g660 ( .A(n_422), .Y(n_660) );
BUFx2_ASAP7_75t_SL g681 ( .A(n_422), .Y(n_681) );
INVx1_ASAP7_75t_L g812 ( .A(n_422), .Y(n_812) );
BUFx2_ASAP7_75t_SL g919 ( .A(n_422), .Y(n_919) );
AND2x4_ASAP7_75t_L g422 ( .A(n_423), .B(n_425), .Y(n_422) );
AND2x2_ASAP7_75t_L g565 ( .A(n_423), .B(n_492), .Y(n_565) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OR2x6_ASAP7_75t_L g438 ( .A(n_424), .B(n_439), .Y(n_438) );
AND2x4_ASAP7_75t_L g448 ( .A(n_425), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g457 ( .A(n_425), .B(n_433), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_425), .B(n_433), .Y(n_632) );
AND2x2_ASAP7_75t_L g473 ( .A(n_426), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g492 ( .A(n_426), .Y(n_492) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx5_ASAP7_75t_L g550 ( .A(n_431), .Y(n_550) );
INVx3_ASAP7_75t_L g558 ( .A(n_431), .Y(n_558) );
INVx1_ASAP7_75t_L g620 ( .A(n_431), .Y(n_620) );
INVx4_ASAP7_75t_L g704 ( .A(n_431), .Y(n_704) );
BUFx3_ASAP7_75t_L g985 ( .A(n_431), .Y(n_985) );
INVx8_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_435), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g742 ( .A(n_433), .B(n_435), .Y(n_742) );
INVx1_ASAP7_75t_L g499 ( .A(n_434), .Y(n_499) );
NAND2x1p5_ASAP7_75t_L g468 ( .A(n_435), .B(n_449), .Y(n_468) );
AND2x6_ASAP7_75t_L g582 ( .A(n_435), .B(n_449), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g858 ( .A(n_436), .Y(n_858) );
BUFx4f_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
BUFx2_ASAP7_75t_L g654 ( .A(n_437), .Y(n_654) );
BUFx2_ASAP7_75t_L g705 ( .A(n_437), .Y(n_705) );
BUFx2_ASAP7_75t_L g1100 ( .A(n_437), .Y(n_1100) );
INVx6_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g551 ( .A(n_438), .Y(n_551) );
INVx1_ASAP7_75t_SL g621 ( .A(n_438), .Y(n_621) );
INVx1_ASAP7_75t_SL g986 ( .A(n_438), .Y(n_986) );
INVx1_ASAP7_75t_L g577 ( .A(n_439), .Y(n_577) );
OAI221xp5_ASAP7_75t_SL g440 ( .A1(n_441), .A2(n_444), .B1(n_445), .B2(n_450), .C(n_451), .Y(n_440) );
INVx2_ASAP7_75t_L g989 ( .A(n_441), .Y(n_989) );
INVx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx6f_ASAP7_75t_L g537 ( .A(n_442), .Y(n_537) );
BUFx3_ASAP7_75t_L g708 ( .A(n_442), .Y(n_708) );
BUFx3_ASAP7_75t_L g913 ( .A(n_442), .Y(n_913) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx2_ASAP7_75t_SL g560 ( .A(n_443), .Y(n_560) );
INVx2_ASAP7_75t_L g657 ( .A(n_443), .Y(n_657) );
BUFx2_ASAP7_75t_SL g683 ( .A(n_443), .Y(n_683) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx3_ASAP7_75t_L g547 ( .A(n_448), .Y(n_547) );
BUFx6f_ASAP7_75t_L g617 ( .A(n_448), .Y(n_617) );
BUFx3_ASAP7_75t_L g658 ( .A(n_448), .Y(n_658) );
INVx2_ASAP7_75t_L g803 ( .A(n_448), .Y(n_803) );
INVx1_ASAP7_75t_L g464 ( .A(n_449), .Y(n_464) );
INVx3_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_453), .A2(n_623), .B1(n_624), .B2(n_625), .Y(n_622) );
INVx2_ASAP7_75t_L g687 ( .A(n_453), .Y(n_687) );
OAI22xp5_ASAP7_75t_SL g806 ( .A1(n_453), .A2(n_657), .B1(n_807), .B2(n_808), .Y(n_806) );
INVx2_ASAP7_75t_L g874 ( .A(n_453), .Y(n_874) );
INVx2_ASAP7_75t_L g960 ( .A(n_453), .Y(n_960) );
OAI221xp5_ASAP7_75t_SL g1131 ( .A1(n_453), .A2(n_630), .B1(n_1132), .B2(n_1133), .C(n_1134), .Y(n_1131) );
INVx6_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx3_ASAP7_75t_L g540 ( .A(n_454), .Y(n_540) );
BUFx3_ASAP7_75t_L g561 ( .A(n_454), .Y(n_561) );
BUFx3_ASAP7_75t_L g785 ( .A(n_454), .Y(n_785) );
BUFx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g701 ( .A(n_456), .Y(n_701) );
BUFx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx3_ASAP7_75t_L g534 ( .A(n_457), .Y(n_534) );
BUFx3_ASAP7_75t_L g684 ( .A(n_457), .Y(n_684) );
BUFx3_ASAP7_75t_L g872 ( .A(n_457), .Y(n_872) );
NOR3xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_469), .C(n_488), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B1(n_465), .B2(n_466), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_461), .A2(n_508), .B1(n_509), .B2(n_510), .Y(n_507) );
OAI221xp5_ASAP7_75t_SL g925 ( .A1(n_461), .A2(n_767), .B1(n_926), .B2(n_927), .C(n_928), .Y(n_925) );
OAI22xp5_ASAP7_75t_L g970 ( .A1(n_461), .A2(n_512), .B1(n_971), .B2(n_972), .Y(n_970) );
OAI22xp5_ASAP7_75t_L g1087 ( .A1(n_461), .A2(n_767), .B1(n_1088), .B2(n_1089), .Y(n_1087) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g639 ( .A(n_462), .Y(n_639) );
INVx1_ASAP7_75t_SL g1040 ( .A(n_462), .Y(n_1040) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx6f_ASAP7_75t_L g765 ( .A(n_463), .Y(n_765) );
OAI21xp5_ASAP7_75t_L g791 ( .A1(n_463), .A2(n_792), .B(n_793), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_466), .A2(n_638), .B1(n_639), .B2(n_640), .Y(n_637) );
OAI22xp5_ASAP7_75t_SL g829 ( .A1(n_466), .A2(n_830), .B1(n_831), .B2(n_832), .Y(n_829) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx3_ASAP7_75t_L g512 ( .A(n_468), .Y(n_512) );
OAI222xp33_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_476), .B1(n_477), .B2(n_481), .C1(n_482), .C2(n_487), .Y(n_469) );
OAI222xp33_ASAP7_75t_L g949 ( .A1(n_470), .A2(n_482), .B1(n_667), .B2(n_950), .C1(n_951), .C2(n_952), .Y(n_949) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_471), .Y(n_470) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_472), .Y(n_520) );
BUFx6f_ASAP7_75t_L g607 ( .A(n_472), .Y(n_607) );
BUFx2_ASAP7_75t_L g645 ( .A(n_472), .Y(n_645) );
BUFx4f_ASAP7_75t_SL g716 ( .A(n_472), .Y(n_716) );
AND2x4_ASAP7_75t_L g472 ( .A(n_473), .B(n_475), .Y(n_472) );
INVx1_ASAP7_75t_L g486 ( .A(n_474), .Y(n_486) );
AND2x4_ASAP7_75t_L g485 ( .A(n_475), .B(n_486), .Y(n_485) );
NAND2x1p5_ASAP7_75t_L g491 ( .A(n_475), .B(n_492), .Y(n_491) );
AND2x4_ASAP7_75t_L g576 ( .A(n_475), .B(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_SL g770 ( .A(n_478), .Y(n_770) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx4_ASAP7_75t_L g515 ( .A(n_479), .Y(n_515) );
INVx2_ASAP7_75t_L g570 ( .A(n_479), .Y(n_570) );
BUFx3_ASAP7_75t_L g594 ( .A(n_479), .Y(n_594) );
INVx2_ASAP7_75t_L g667 ( .A(n_479), .Y(n_667) );
INVx2_ASAP7_75t_SL g799 ( .A(n_479), .Y(n_799) );
INVx1_ASAP7_75t_L g497 ( .A(n_480), .Y(n_497) );
AND2x4_ASAP7_75t_L g572 ( .A(n_480), .B(n_499), .Y(n_572) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g933 ( .A(n_484), .Y(n_933) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx12f_ASAP7_75t_L g524 ( .A(n_485), .Y(n_524) );
BUFx6f_ASAP7_75t_L g727 ( .A(n_485), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B1(n_493), .B2(n_494), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_490), .A2(n_526), .B1(n_527), .B2(n_528), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g976 ( .A1(n_490), .A2(n_977), .B1(n_978), .B2(n_979), .Y(n_976) );
BUFx3_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx4_ASAP7_75t_L g649 ( .A(n_491), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_491), .A2(n_606), .B1(n_773), .B2(n_774), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g794 ( .A1(n_491), .A2(n_512), .B1(n_795), .B2(n_796), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g860 ( .A1(n_491), .A2(n_494), .B1(n_861), .B2(n_862), .Y(n_860) );
HB1xp67_ASAP7_75t_L g1048 ( .A(n_491), .Y(n_1048) );
OAI22xp5_ASAP7_75t_L g1093 ( .A1(n_491), .A2(n_528), .B1(n_1094), .B2(n_1095), .Y(n_1093) );
OAI22xp5_ASAP7_75t_L g1145 ( .A1(n_494), .A2(n_648), .B1(n_1146), .B2(n_1147), .Y(n_1145) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g979 ( .A(n_495), .Y(n_979) );
CKINVDCx16_ASAP7_75t_R g495 ( .A(n_496), .Y(n_495) );
BUFx2_ASAP7_75t_L g528 ( .A(n_496), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_496), .A2(n_647), .B1(n_648), .B2(n_650), .Y(n_646) );
OR2x6_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_553), .B1(n_554), .B2(n_584), .Y(n_502) );
INVx1_ASAP7_75t_L g584 ( .A(n_503), .Y(n_584) );
INVx1_ASAP7_75t_L g552 ( .A(n_505), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_529), .Y(n_505) );
NOR3xp33_ASAP7_75t_L g506 ( .A(n_507), .B(n_513), .C(n_525), .Y(n_506) );
OAI211xp5_ASAP7_75t_L g595 ( .A1(n_510), .A2(n_596), .B(n_597), .C(n_599), .Y(n_595) );
OAI221xp5_ASAP7_75t_L g945 ( .A1(n_510), .A2(n_639), .B1(n_946), .B2(n_947), .C(n_948), .Y(n_945) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx3_ASAP7_75t_L g767 ( .A(n_512), .Y(n_767) );
OA211x2_ASAP7_75t_L g894 ( .A1(n_512), .A2(n_895), .B(n_896), .C(n_898), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g1038 ( .A1(n_512), .A2(n_1039), .B1(n_1040), .B2(n_1041), .Y(n_1038) );
OAI22xp5_ASAP7_75t_L g1136 ( .A1(n_512), .A2(n_1040), .B1(n_1137), .B2(n_1138), .Y(n_1136) );
OAI221xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_516), .B1(n_517), .B2(n_521), .C(n_522), .Y(n_513) );
BUFx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OAI22xp5_ASAP7_75t_SL g836 ( .A1(n_515), .A2(n_837), .B1(n_838), .B2(n_839), .Y(n_836) );
INVx4_ASAP7_75t_L g884 ( .A(n_515), .Y(n_884) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g797 ( .A1(n_519), .A2(n_798), .B1(n_799), .B2(n_800), .Y(n_797) );
INVx4_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g838 ( .A(n_520), .Y(n_838) );
BUFx4f_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g611 ( .A(n_524), .Y(n_611) );
NOR2xp67_ASAP7_75t_L g529 ( .A(n_530), .B(n_541), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_536), .Y(n_530) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
BUFx4f_ASAP7_75t_SL g779 ( .A(n_534), .Y(n_779) );
BUFx2_ASAP7_75t_L g962 ( .A(n_535), .Y(n_962) );
INVx1_ASAP7_75t_SL g628 ( .A(n_537), .Y(n_628) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_548), .Y(n_541) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g680 ( .A(n_546), .Y(n_680) );
INVx5_ASAP7_75t_SL g778 ( .A(n_546), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g816 ( .A(n_546), .B(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g908 ( .A(n_546), .Y(n_908) );
BUFx2_ASAP7_75t_L g852 ( .A(n_547), .Y(n_852) );
BUFx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
BUFx6f_ASAP7_75t_L g689 ( .A(n_550), .Y(n_689) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
XOR2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_583), .Y(n_554) );
NAND4xp75_ASAP7_75t_SL g555 ( .A(n_556), .B(n_559), .C(n_562), .D(n_567), .Y(n_555) );
INVx1_ASAP7_75t_L g624 ( .A(n_557), .Y(n_624) );
INVx1_ASAP7_75t_L g910 ( .A(n_561), .Y(n_910) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_566), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_568), .B(n_573), .Y(n_567) );
OAI21xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_570), .B(n_571), .Y(n_568) );
OAI222xp33_ASAP7_75t_L g722 ( .A1(n_570), .A2(n_723), .B1(n_724), .B2(n_725), .C1(n_726), .C2(n_728), .Y(n_722) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_572), .Y(n_603) );
BUFx3_ASAP7_75t_L g731 ( .A(n_572), .Y(n_731) );
BUFx2_ASAP7_75t_SL g1003 ( .A(n_572), .Y(n_1003) );
BUFx2_ASAP7_75t_SL g1064 ( .A(n_572), .Y(n_1064) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_578), .Y(n_573) );
BUFx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
BUFx2_ASAP7_75t_L g600 ( .A(n_576), .Y(n_600) );
INVx1_ASAP7_75t_L g676 ( .A(n_576), .Y(n_676) );
BUFx2_ASAP7_75t_L g878 ( .A(n_576), .Y(n_878) );
BUFx6f_ASAP7_75t_L g713 ( .A(n_579), .Y(n_713) );
INVx5_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g598 ( .A(n_580), .Y(n_598) );
INVx2_ASAP7_75t_L g897 ( .A(n_580), .Y(n_897) );
INVx4_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
BUFx2_ASAP7_75t_L g673 ( .A(n_582), .Y(n_673) );
BUFx4f_ASAP7_75t_L g735 ( .A(n_582), .Y(n_735) );
BUFx2_ASAP7_75t_L g1015 ( .A(n_582), .Y(n_1015) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OAI22xp5_ASAP7_75t_SL g586 ( .A1(n_587), .A2(n_693), .B1(n_694), .B2(n_753), .Y(n_586) );
INVx2_ASAP7_75t_SL g753 ( .A(n_587), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B1(n_633), .B2(n_692), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_589), .A2(n_590), .B1(n_719), .B2(n_750), .Y(n_718) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
XNOR2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_612), .Y(n_592) );
INVx3_ASAP7_75t_L g643 ( .A(n_594), .Y(n_643) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_606), .B1(n_608), .B2(n_609), .Y(n_604) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_607), .Y(n_670) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx3_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NOR3xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_622), .C(n_626), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_619), .Y(n_613) );
INVx3_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx4_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_628), .B1(n_629), .B2(n_630), .Y(n_626) );
OAI221xp5_ASAP7_75t_SL g1126 ( .A1(n_628), .A2(n_1127), .B1(n_1128), .B2(n_1129), .C(n_1130), .Y(n_1126) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g814 ( .A(n_632), .B(n_815), .Y(n_814) );
INVx2_ASAP7_75t_L g692 ( .A(n_633), .Y(n_692) );
XNOR2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_663), .Y(n_633) );
INVx1_ASAP7_75t_SL g661 ( .A(n_635), .Y(n_661) );
AND2x2_ASAP7_75t_SL g635 ( .A(n_636), .B(n_651), .Y(n_635) );
NOR3xp33_ASAP7_75t_L g636 ( .A(n_637), .B(n_641), .C(n_646), .Y(n_636) );
OAI21xp33_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_643), .B(n_644), .Y(n_641) );
OAI21xp33_ASAP7_75t_L g973 ( .A1(n_643), .A2(n_974), .B(n_975), .Y(n_973) );
INVx1_ASAP7_75t_L g1141 ( .A(n_645), .Y(n_1141) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx3_ASAP7_75t_SL g831 ( .A(n_649), .Y(n_831) );
AND4x1_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .C(n_655), .D(n_659), .Y(n_651) );
INVx3_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx3_ASAP7_75t_L g881 ( .A(n_657), .Y(n_881) );
BUFx2_ASAP7_75t_L g916 ( .A(n_658), .Y(n_916) );
INVx2_ASAP7_75t_SL g690 ( .A(n_664), .Y(n_690) );
AND2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_677), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_666), .B(n_671), .Y(n_665) );
OAI21xp5_ASAP7_75t_SL g666 ( .A1(n_667), .A2(n_668), .B(n_669), .Y(n_666) );
OAI21xp5_ASAP7_75t_L g1000 ( .A1(n_667), .A2(n_1001), .B(n_1002), .Y(n_1000) );
OAI21xp5_ASAP7_75t_SL g1018 ( .A1(n_667), .A2(n_1019), .B(n_1020), .Y(n_1018) );
OAI21xp5_ASAP7_75t_L g1061 ( .A1(n_667), .A2(n_1062), .B(n_1063), .Y(n_1061) );
INVx2_ASAP7_75t_SL g724 ( .A(n_670), .Y(n_724) );
NAND2xp5_ASAP7_75t_SL g671 ( .A(n_672), .B(n_674), .Y(n_671) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_678), .B(n_685), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_679), .B(n_682), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_688), .Y(n_685) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_718), .B1(n_751), .B2(n_752), .Y(n_694) );
INVx1_ASAP7_75t_L g752 ( .A(n_695), .Y(n_752) );
INVx1_ASAP7_75t_SL g717 ( .A(n_697), .Y(n_717) );
NAND4xp75_ASAP7_75t_L g697 ( .A(n_698), .B(n_706), .C(n_711), .D(n_715), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_702), .Y(n_698) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
BUFx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g923 ( .A(n_704), .Y(n_923) );
INVx1_ASAP7_75t_L g744 ( .A(n_705), .Y(n_744) );
AND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_710), .Y(n_706) );
INVx1_ASAP7_75t_L g1128 ( .A(n_709), .Y(n_1128) );
AND2x2_ASAP7_75t_SL g711 ( .A(n_712), .B(n_714), .Y(n_711) );
INVx1_ASAP7_75t_L g930 ( .A(n_716), .Y(n_930) );
INVx1_ASAP7_75t_L g751 ( .A(n_718), .Y(n_751) );
INVx1_ASAP7_75t_L g750 ( .A(n_719), .Y(n_750) );
NAND3x1_ASAP7_75t_L g720 ( .A(n_721), .B(n_736), .C(n_739), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_729), .Y(n_721) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
BUFx4f_ASAP7_75t_L g1144 ( .A(n_727), .Y(n_1144) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_732), .Y(n_729) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .Y(n_736) );
OAI22xp5_ASAP7_75t_SL g740 ( .A1(n_741), .A2(n_743), .B1(n_744), .B2(n_745), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g855 ( .A1(n_741), .A2(n_856), .B1(n_857), .B2(n_858), .Y(n_855) );
BUFx2_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g810 ( .A1(n_742), .A2(n_811), .B1(n_812), .B2(n_813), .Y(n_810) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
AO22x2_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_758), .B1(n_787), .B2(n_840), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g761 ( .A(n_762), .B(n_775), .Y(n_761) );
NOR3xp33_ASAP7_75t_L g762 ( .A(n_763), .B(n_768), .C(n_772), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_765), .B1(n_766), .B2(n_767), .Y(n_763) );
OAI21xp5_ASAP7_75t_SL g833 ( .A1(n_765), .A2(n_834), .B(n_835), .Y(n_833) );
OAI21xp33_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_770), .B(n_771), .Y(n_768) );
OAI21xp33_ASAP7_75t_L g1042 ( .A1(n_770), .A2(n_1043), .B(n_1044), .Y(n_1042) );
OAI21xp33_ASAP7_75t_SL g1090 ( .A1(n_770), .A2(n_1091), .B(n_1092), .Y(n_1090) );
OAI221xp5_ASAP7_75t_SL g1139 ( .A1(n_770), .A2(n_1140), .B1(n_1141), .B2(n_1142), .C(n_1143), .Y(n_1139) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_776), .B(n_781), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_777), .B(n_780), .Y(n_776) );
INVx1_ASAP7_75t_L g1104 ( .A(n_778), .Y(n_1104) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_782), .B(n_786), .Y(n_781) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx3_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx2_ASAP7_75t_L g840 ( .A(n_787), .Y(n_840) );
XOR2x2_ASAP7_75t_L g787 ( .A(n_788), .B(n_819), .Y(n_787) );
XNOR2x1_ASAP7_75t_L g788 ( .A(n_789), .B(n_818), .Y(n_788) );
AND3x2_ASAP7_75t_L g789 ( .A(n_790), .B(n_801), .C(n_809), .Y(n_789) );
NOR3xp33_ASAP7_75t_L g790 ( .A(n_791), .B(n_794), .C(n_797), .Y(n_790) );
OAI222xp33_ASAP7_75t_L g929 ( .A1(n_799), .A2(n_930), .B1(n_931), .B2(n_932), .C1(n_933), .C2(n_934), .Y(n_929) );
NOR2xp33_ASAP7_75t_L g801 ( .A(n_802), .B(n_806), .Y(n_801) );
OAI21xp5_ASAP7_75t_SL g802 ( .A1(n_803), .A2(n_804), .B(n_805), .Y(n_802) );
INVx1_ASAP7_75t_L g956 ( .A(n_803), .Y(n_956) );
INVx2_ASAP7_75t_L g982 ( .A(n_803), .Y(n_982) );
NOR3xp33_ASAP7_75t_L g809 ( .A(n_810), .B(n_814), .C(n_816), .Y(n_809) );
XNOR2xp5_ASAP7_75t_L g819 ( .A(n_820), .B(n_821), .Y(n_819) );
NAND3x1_ASAP7_75t_SL g821 ( .A(n_822), .B(n_825), .C(n_828), .Y(n_821) );
AND2x2_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .Y(n_822) );
AND2x2_ASAP7_75t_L g825 ( .A(n_826), .B(n_827), .Y(n_825) );
NOR3xp33_ASAP7_75t_L g828 ( .A(n_829), .B(n_833), .C(n_836), .Y(n_828) );
INVx1_ASAP7_75t_L g1108 ( .A(n_841), .Y(n_1108) );
XNOR2xp5_ASAP7_75t_L g841 ( .A(n_842), .B(n_938), .Y(n_841) );
HB1xp67_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
XNOR2xp5_ASAP7_75t_SL g843 ( .A(n_844), .B(n_865), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx2_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
AND4x1_ASAP7_75t_L g849 ( .A(n_850), .B(n_854), .C(n_859), .D(n_863), .Y(n_849) );
AOI22xp5_ASAP7_75t_L g865 ( .A1(n_866), .A2(n_867), .B1(n_903), .B2(n_937), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
AO22x1_ASAP7_75t_SL g867 ( .A1(n_868), .A2(n_886), .B1(n_901), .B2(n_902), .Y(n_867) );
INVx2_ASAP7_75t_SL g901 ( .A(n_868), .Y(n_901) );
XOR2x2_ASAP7_75t_L g868 ( .A(n_869), .B(n_885), .Y(n_868) );
NAND4xp75_ASAP7_75t_L g869 ( .A(n_870), .B(n_875), .C(n_879), .D(n_883), .Y(n_869) );
AND2x2_ASAP7_75t_L g870 ( .A(n_871), .B(n_873), .Y(n_870) );
AND2x2_ASAP7_75t_SL g875 ( .A(n_876), .B(n_877), .Y(n_875) );
AND2x2_ASAP7_75t_L g879 ( .A(n_880), .B(n_882), .Y(n_879) );
INVx2_ASAP7_75t_SL g902 ( .A(n_886), .Y(n_902) );
XOR2x2_ASAP7_75t_L g886 ( .A(n_887), .B(n_900), .Y(n_886) );
NAND4xp75_ASAP7_75t_L g887 ( .A(n_888), .B(n_891), .C(n_894), .D(n_899), .Y(n_887) );
AND2x2_ASAP7_75t_L g888 ( .A(n_889), .B(n_890), .Y(n_888) );
AND2x2_ASAP7_75t_L g891 ( .A(n_892), .B(n_893), .Y(n_891) );
INVx1_ASAP7_75t_L g937 ( .A(n_903), .Y(n_937) );
INVx1_ASAP7_75t_L g936 ( .A(n_904), .Y(n_936) );
AND2x2_ASAP7_75t_L g904 ( .A(n_905), .B(n_924), .Y(n_904) );
NOR2xp33_ASAP7_75t_L g905 ( .A(n_906), .B(n_914), .Y(n_905) );
OAI221xp5_ASAP7_75t_SL g906 ( .A1(n_907), .A2(n_909), .B1(n_910), .B2(n_911), .C(n_912), .Y(n_906) );
INVx2_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
OAI221xp5_ASAP7_75t_SL g914 ( .A1(n_915), .A2(n_917), .B1(n_918), .B2(n_920), .C(n_921), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
INVx3_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
NOR2xp33_ASAP7_75t_SL g924 ( .A(n_925), .B(n_929), .Y(n_924) );
OAI22xp5_ASAP7_75t_L g1045 ( .A1(n_930), .A2(n_1046), .B1(n_1047), .B2(n_1048), .Y(n_1045) );
AOI22xp5_ASAP7_75t_SL g938 ( .A1(n_939), .A2(n_1078), .B1(n_1079), .B2(n_1106), .Y(n_938) );
INVx1_ASAP7_75t_L g1106 ( .A(n_939), .Y(n_1106) );
AOI22xp5_ASAP7_75t_L g939 ( .A1(n_940), .A2(n_941), .B1(n_965), .B2(n_1077), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
INVx1_ASAP7_75t_SL g964 ( .A(n_943), .Y(n_964) );
AND2x2_ASAP7_75t_L g943 ( .A(n_944), .B(n_953), .Y(n_943) );
NOR2xp33_ASAP7_75t_SL g944 ( .A(n_945), .B(n_949), .Y(n_944) );
NOR2xp33_ASAP7_75t_L g953 ( .A(n_954), .B(n_958), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_955), .B(n_957), .Y(n_954) );
NAND2xp5_ASAP7_75t_SL g958 ( .A(n_959), .B(n_961), .Y(n_958) );
INVx1_ASAP7_75t_L g1077 ( .A(n_965), .Y(n_1077) );
XOR2xp5_ASAP7_75t_L g965 ( .A(n_966), .B(n_1031), .Y(n_965) );
OA22x2_ASAP7_75t_L g966 ( .A1(n_967), .A2(n_992), .B1(n_1029), .B2(n_1030), .Y(n_966) );
INVx1_ASAP7_75t_L g1029 ( .A(n_967), .Y(n_1029) );
INVx2_ASAP7_75t_SL g990 ( .A(n_968), .Y(n_990) );
AND2x2_ASAP7_75t_SL g968 ( .A(n_969), .B(n_980), .Y(n_968) );
NOR3xp33_ASAP7_75t_L g969 ( .A(n_970), .B(n_973), .C(n_976), .Y(n_969) );
AND4x1_ASAP7_75t_L g980 ( .A(n_981), .B(n_983), .C(n_987), .D(n_988), .Y(n_980) );
INVx3_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
INVx1_ASAP7_75t_L g1030 ( .A(n_992), .Y(n_1030) );
XOR2x2_ASAP7_75t_L g992 ( .A(n_993), .B(n_1010), .Y(n_992) );
OA22x2_ASAP7_75t_L g1031 ( .A1(n_993), .A2(n_1032), .B1(n_1033), .B2(n_1076), .Y(n_1031) );
INVx1_ASAP7_75t_L g1032 ( .A(n_993), .Y(n_1032) );
XOR2x2_ASAP7_75t_L g993 ( .A(n_994), .B(n_1009), .Y(n_993) );
NAND4xp75_ASAP7_75t_SL g994 ( .A(n_995), .B(n_1004), .C(n_1007), .D(n_1008), .Y(n_994) );
NOR2xp67_ASAP7_75t_SL g995 ( .A(n_996), .B(n_1000), .Y(n_995) );
NAND3xp33_ASAP7_75t_L g996 ( .A(n_997), .B(n_998), .C(n_999), .Y(n_996) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1006), .Y(n_1004) );
XOR2x2_ASAP7_75t_SL g1010 ( .A(n_1011), .B(n_1028), .Y(n_1010) );
NAND2x1p5_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1021), .Y(n_1011) );
NOR2xp33_ASAP7_75t_L g1012 ( .A(n_1013), .B(n_1018), .Y(n_1012) );
NAND3xp33_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1016), .C(n_1017), .Y(n_1013) );
NOR2x1_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1025), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1024), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1027), .Y(n_1025) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1033), .Y(n_1076) );
OAI22xp5_ASAP7_75t_L g1033 ( .A1(n_1034), .A2(n_1035), .B1(n_1057), .B2(n_1058), .Y(n_1033) );
INVx1_ASAP7_75t_SL g1034 ( .A(n_1035), .Y(n_1034) );
XNOR2x1_ASAP7_75t_L g1035 ( .A(n_1036), .B(n_1056), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_1037), .B(n_1049), .Y(n_1036) );
NOR3xp33_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1042), .C(n_1045), .Y(n_1037) );
NOR2xp33_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1053), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g1050 ( .A(n_1051), .B(n_1052), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1055), .Y(n_1053) );
AO22x1_ASAP7_75t_L g1080 ( .A1(n_1057), .A2(n_1058), .B1(n_1081), .B2(n_1082), .Y(n_1080) );
INVx3_ASAP7_75t_SL g1057 ( .A(n_1058), .Y(n_1057) );
XOR2x2_ASAP7_75t_L g1058 ( .A(n_1059), .B(n_1075), .Y(n_1058) );
NAND2xp5_ASAP7_75t_SL g1059 ( .A(n_1060), .B(n_1068), .Y(n_1059) );
NOR2xp33_ASAP7_75t_L g1060 ( .A(n_1061), .B(n_1065), .Y(n_1060) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_1066), .B(n_1067), .Y(n_1065) );
NOR2xp33_ASAP7_75t_L g1068 ( .A(n_1069), .B(n_1072), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1071), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_1073), .B(n_1074), .Y(n_1072) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
BUFx2_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
INVx1_ASAP7_75t_SL g1084 ( .A(n_1085), .Y(n_1084) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1096), .Y(n_1085) );
NOR3xp33_ASAP7_75t_L g1086 ( .A(n_1087), .B(n_1090), .C(n_1093), .Y(n_1086) );
NOR2xp33_ASAP7_75t_L g1096 ( .A(n_1097), .B(n_1101), .Y(n_1096) );
NAND2xp5_ASAP7_75t_L g1097 ( .A(n_1098), .B(n_1099), .Y(n_1097) );
NAND2xp5_ASAP7_75t_L g1101 ( .A(n_1102), .B(n_1105), .Y(n_1101) );
INVx2_ASAP7_75t_L g1103 ( .A(n_1104), .Y(n_1103) );
INVx1_ASAP7_75t_SL g1109 ( .A(n_1110), .Y(n_1109) );
NOR2x1_ASAP7_75t_L g1110 ( .A(n_1111), .B(n_1115), .Y(n_1110) );
OR2x2_ASAP7_75t_SL g1163 ( .A(n_1111), .B(n_1116), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1111 ( .A(n_1112), .B(n_1114), .Y(n_1111) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
HB1xp67_ASAP7_75t_L g1150 ( .A(n_1113), .Y(n_1150) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1113), .B(n_1154), .Y(n_1157) );
CKINVDCx16_ASAP7_75t_R g1154 ( .A(n_1114), .Y(n_1154) );
CKINVDCx20_ASAP7_75t_R g1115 ( .A(n_1116), .Y(n_1115) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_1117), .B(n_1118), .Y(n_1116) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1121), .Y(n_1119) );
OAI322xp33_ASAP7_75t_L g1122 ( .A1(n_1123), .A2(n_1150), .A3(n_1151), .B1(n_1155), .B2(n_1158), .C1(n_1159), .C2(n_1163), .Y(n_1122) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1124), .Y(n_1149) );
AND2x2_ASAP7_75t_SL g1124 ( .A(n_1125), .B(n_1135), .Y(n_1124) );
NOR2xp33_ASAP7_75t_L g1125 ( .A(n_1126), .B(n_1131), .Y(n_1125) );
NOR3xp33_ASAP7_75t_L g1135 ( .A(n_1136), .B(n_1139), .C(n_1145), .Y(n_1135) );
BUFx2_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
HB1xp67_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
CKINVDCx16_ASAP7_75t_R g1155 ( .A(n_1156), .Y(n_1155) );
INVx1_ASAP7_75t_SL g1159 ( .A(n_1160), .Y(n_1159) );
BUFx2_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
endmodule