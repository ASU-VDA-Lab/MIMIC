module fake_jpeg_28935_n_129 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_129);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_121;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_59),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_46),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_1),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_62),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_54),
.A2(n_23),
.B1(n_41),
.B2(n_40),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_63),
.B1(n_55),
.B2(n_4),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_1),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_46),
.Y(n_70)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_70),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_48),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_55),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_75),
.Y(n_81)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NAND3xp33_ASAP7_75t_SL g75 ( 
.A(n_61),
.B(n_46),
.C(n_44),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

AO21x1_ASAP7_75t_L g83 ( 
.A1(n_77),
.A2(n_56),
.B(n_6),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_69),
.B(n_53),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_82),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_3),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_83),
.A2(n_13),
.B1(n_19),
.B2(n_20),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_77),
.A2(n_56),
.B1(n_51),
.B2(n_50),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_77),
.A2(n_49),
.B1(n_43),
.B2(n_5),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_92),
.B(n_22),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_5),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_91),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_7),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_89),
.B(n_27),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_7),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_9),
.B(n_10),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_80),
.B(n_11),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_96),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_88),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_95),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_79),
.B(n_12),
.Y(n_96)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_66),
.B(n_16),
.Y(n_97)
);

NAND3xp33_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_98),
.C(n_100),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_85),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_84),
.Y(n_101)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_104),
.C(n_106),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_26),
.Y(n_104)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_28),
.C(n_29),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_107),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_84),
.B(n_34),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_109),
.C(n_110),
.Y(n_113)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_35),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_111),
.A2(n_110),
.B1(n_104),
.B2(n_42),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_121),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

NAND3xp33_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_122),
.C(n_97),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_102),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_113),
.C(n_99),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_123),
.C(n_112),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_126),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_127),
.A2(n_122),
.B(n_118),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_117),
.Y(n_129)
);


endmodule