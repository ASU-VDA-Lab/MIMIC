module fake_jpeg_13448_n_179 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_179);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_19),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_12),
.B(n_44),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_6),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_34),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_6),
.B(n_3),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx6_ASAP7_75t_SL g69 ( 
.A(n_35),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_36),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_9),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_0),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_14),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_50),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_10),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_83),
.Y(n_92)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_67),
.B(n_0),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_56),
.Y(n_84)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_88),
.Y(n_97)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx4_ASAP7_75t_SL g88 ( 
.A(n_60),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_52),
.B(n_1),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_71),
.Y(n_103)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_76),
.B1(n_51),
.B2(n_75),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_99),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_84),
.A2(n_74),
.B1(n_75),
.B2(n_82),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_94),
.A2(n_73),
.B(n_62),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_76),
.B1(n_51),
.B2(n_74),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_84),
.B(n_56),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_72),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_89),
.B1(n_65),
.B2(n_55),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_62),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_91),
.A2(n_65),
.B1(n_55),
.B2(n_64),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_105),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_88),
.B(n_59),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_108),
.A2(n_125),
.B1(n_61),
.B2(n_54),
.Y(n_140)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_112),
.B(n_118),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_100),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_116),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_97),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_103),
.A2(n_94),
.B(n_92),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_57),
.C(n_63),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_79),
.Y(n_118)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_122),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_121),
.A2(n_4),
.B(n_5),
.Y(n_145)
);

BUFx24_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_124),
.Y(n_134)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_114),
.A2(n_72),
.B1(n_58),
.B2(n_77),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_127),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_146)
);

AND2x4_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_78),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_145),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_135),
.A2(n_137),
.B(n_18),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_70),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_143),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_SL g137 ( 
.A1(n_113),
.A2(n_29),
.B(n_48),
.C(n_46),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_121),
.B(n_120),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_138),
.B(n_141),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_140),
.A2(n_142),
.B1(n_24),
.B2(n_25),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_53),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_2),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_134),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_149),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_128),
.A2(n_27),
.B1(n_40),
.B2(n_39),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_148),
.A2(n_157),
.B(n_139),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_126),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_7),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_154),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_138),
.A2(n_8),
.B1(n_11),
.B2(n_15),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_155),
.A2(n_159),
.B(n_137),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_16),
.Y(n_156)
);

A2O1A1O1Ixp25_ASAP7_75t_L g166 ( 
.A1(n_156),
.A2(n_30),
.B(n_31),
.C(n_32),
.D(n_33),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_130),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_41),
.C(n_21),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_160),
.C(n_137),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_164),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_165),
.B(n_166),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_157),
.C(n_150),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_170),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_152),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_171),
.A2(n_167),
.B(n_161),
.C(n_168),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_172),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_158),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_151),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_161),
.C(n_148),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_177),
.A2(n_133),
.B1(n_144),
.B2(n_150),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_146),
.Y(n_179)
);


endmodule