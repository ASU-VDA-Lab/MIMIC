module fake_jpeg_691_n_184 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_184);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_31),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx11_ASAP7_75t_SL g57 ( 
.A(n_10),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx11_ASAP7_75t_SL g60 ( 
.A(n_44),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_12),
.Y(n_66)
);

CKINVDCx9p33_ASAP7_75t_R g67 ( 
.A(n_57),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_SL g68 ( 
.A1(n_61),
.A2(n_46),
.B(n_43),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_59),
.Y(n_78)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_0),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_53),
.Y(n_79)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_73),
.A2(n_59),
.B1(n_65),
.B2(n_48),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_54),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_74),
.B(n_71),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_61),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_83),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_73),
.A2(n_53),
.B1(n_65),
.B2(n_62),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_77),
.A2(n_81),
.B(n_69),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_84),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_79),
.B(n_69),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_72),
.A2(n_58),
.B1(n_62),
.B2(n_51),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_56),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_74),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_89),
.A2(n_81),
.B1(n_69),
.B2(n_72),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_82),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_90),
.B(n_82),
.Y(n_107)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_98),
.Y(n_110)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx3_ASAP7_75t_SL g97 ( 
.A(n_80),
.Y(n_97)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_76),
.B(n_50),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_100),
.Y(n_120)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_102),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_55),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_104),
.Y(n_115)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_105),
.A2(n_119),
.B1(n_28),
.B2(n_41),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_47),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_113),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_107),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_63),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_108),
.B(n_6),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_68),
.B(n_73),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_27),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_54),
.B(n_48),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_52),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_35),
.Y(n_128)
);

NAND2xp33_ASAP7_75t_SL g116 ( 
.A(n_96),
.B(n_100),
.Y(n_116)
);

NAND3xp33_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_7),
.C(n_8),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_92),
.A2(n_51),
.B1(n_49),
.B2(n_2),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_117),
.A2(n_121),
.B1(n_4),
.B2(n_5),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_97),
.A2(n_49),
.B1(n_1),
.B2(n_2),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_127),
.B1(n_13),
.B2(n_14),
.Y(n_153)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_128),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_42),
.B1(n_40),
.B2(n_38),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_34),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_141),
.Y(n_154)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_133),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_112),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_138),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_135),
.A2(n_136),
.B1(n_119),
.B2(n_14),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_110),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_137),
.A2(n_121),
.B(n_20),
.Y(n_148)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_26),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_142),
.A2(n_143),
.B(n_144),
.Y(n_151)
);

OAI32xp33_ASAP7_75t_L g143 ( 
.A1(n_106),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_11),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_SL g147 ( 
.A1(n_126),
.A2(n_116),
.B(n_113),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_150),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_148),
.B(n_153),
.Y(n_164)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_21),
.C(n_23),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_126),
.A2(n_140),
.B1(n_124),
.B2(n_127),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_157),
.A2(n_128),
.B1(n_135),
.B2(n_131),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_161),
.A2(n_166),
.B1(n_154),
.B2(n_152),
.Y(n_169)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_145),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_163),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_151),
.A2(n_143),
.B(n_136),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_146),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_165),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_149),
.B(n_15),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_159),
.Y(n_168)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_168),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_169),
.A2(n_171),
.B(n_158),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_147),
.B1(n_159),
.B2(n_158),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_173),
.A2(n_168),
.B1(n_171),
.B2(n_167),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_167),
.C(n_156),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_174),
.B(n_170),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_176),
.A2(n_177),
.B1(n_175),
.B2(n_164),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_155),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_179),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_180),
.B(n_16),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_17),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_18),
.C(n_24),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_18),
.Y(n_184)
);


endmodule