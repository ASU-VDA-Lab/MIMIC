module fake_jpeg_1647_n_462 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_462);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_462;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_387;
wire n_270;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_15),
.B(n_9),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_53),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_54),
.B(n_66),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_55),
.B(n_56),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_26),
.B(n_0),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_57),
.Y(n_154)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_58),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_60),
.Y(n_140)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g177 ( 
.A(n_63),
.Y(n_177)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_64),
.Y(n_164)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_24),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_67),
.B(n_68),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_42),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_0),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_69),
.B(n_70),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_34),
.B(n_1),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_22),
.B(n_41),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_71),
.B(n_76),
.Y(n_162)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g174 ( 
.A(n_72),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_42),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_73),
.B(n_80),
.Y(n_121)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_74),
.Y(n_168)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_22),
.B(n_1),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_37),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_81),
.Y(n_169)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_83),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_37),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_84),
.B(n_102),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g182 ( 
.A(n_85),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_87),
.Y(n_124)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_88),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_35),
.B(n_3),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_89),
.B(n_107),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_47),
.Y(n_90)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx4_ASAP7_75t_SL g91 ( 
.A(n_47),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_91),
.Y(n_178)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_93),
.Y(n_152)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_97),
.Y(n_159)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_98),
.Y(n_179)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_100),
.Y(n_175)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_32),
.Y(n_101)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_101),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_36),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

BUFx2_ASAP7_75t_SL g163 ( 
.A(n_104),
.Y(n_163)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_32),
.Y(n_106)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_37),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_109),
.Y(n_165)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_21),
.Y(n_110)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_110),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_45),
.Y(n_111)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_111),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_46),
.Y(n_112)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_112),
.Y(n_181)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_113),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_59),
.A2(n_46),
.B1(n_43),
.B2(n_38),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_118),
.A2(n_157),
.B1(n_12),
.B2(n_13),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_81),
.A2(n_41),
.B1(n_49),
.B2(n_46),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_126),
.A2(n_131),
.B1(n_136),
.B2(n_146),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_58),
.B(n_36),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_129),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_60),
.A2(n_49),
.B1(n_20),
.B2(n_39),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_61),
.A2(n_39),
.B1(n_38),
.B2(n_31),
.Y(n_135)
);

AO21x1_ASAP7_75t_L g186 ( 
.A1(n_135),
.A2(n_153),
.B(n_160),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_78),
.A2(n_43),
.B1(n_50),
.B2(n_51),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_91),
.A2(n_51),
.B1(n_50),
.B2(n_33),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_83),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_151),
.B(n_158),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_92),
.A2(n_25),
.B1(n_31),
.B2(n_29),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_85),
.A2(n_19),
.B1(n_29),
.B2(n_20),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_62),
.B(n_33),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_86),
.A2(n_21),
.B1(n_25),
.B2(n_19),
.Y(n_160)
);

AND2x2_ASAP7_75t_SL g161 ( 
.A(n_101),
.B(n_17),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_161),
.Y(n_243)
);

AOI21xp33_ASAP7_75t_L g170 ( 
.A1(n_63),
.A2(n_17),
.B(n_27),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_4),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_90),
.A2(n_27),
.B1(n_17),
.B2(n_5),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_171),
.A2(n_172),
.B1(n_176),
.B2(n_184),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_98),
.A2(n_27),
.B1(n_4),
.B2(n_5),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_74),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_113),
.B(n_3),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_180),
.B(n_129),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_99),
.A2(n_97),
.B1(n_100),
.B2(n_75),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_104),
.Y(n_185)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_187),
.Y(n_261)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_188),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_189),
.Y(n_256)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_190),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_191),
.B(n_195),
.Y(n_287)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_130),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_192),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_193),
.B(n_209),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_117),
.B(n_64),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_165),
.Y(n_196)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_196),
.Y(n_285)
);

O2A1O1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_118),
.A2(n_95),
.B(n_77),
.C(n_63),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_198),
.A2(n_179),
.B(n_174),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_121),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_199),
.B(n_206),
.Y(n_257)
);

OAI32xp33_ASAP7_75t_L g200 ( 
.A1(n_138),
.A2(n_57),
.A3(n_112),
.B1(n_111),
.B2(n_109),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_200),
.A2(n_239),
.B(n_172),
.Y(n_252)
);

AND2x2_ASAP7_75t_SL g201 ( 
.A(n_116),
.B(n_79),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_201),
.Y(n_253)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_114),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_202),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_115),
.B(n_79),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_203),
.B(n_215),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_139),
.A2(n_108),
.B1(n_96),
.B2(n_7),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_204),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_147),
.B(n_4),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_205),
.B(n_213),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_162),
.B(n_6),
.Y(n_206)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_130),
.Y(n_208)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_208),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_114),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_210),
.Y(n_249)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_127),
.Y(n_211)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_211),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_150),
.B(n_6),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_212),
.B(n_222),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_6),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_139),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_214),
.A2(n_237),
.B1(n_238),
.B2(n_241),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_166),
.B(n_8),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_181),
.Y(n_216)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_216),
.Y(n_266)
);

BUFx12f_ASAP7_75t_SL g217 ( 
.A(n_174),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_217),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_140),
.Y(n_218)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_218),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_161),
.B(n_8),
.Y(n_219)
);

AND2x2_ASAP7_75t_SL g264 ( 
.A(n_219),
.B(n_122),
.Y(n_264)
);

OR2x4_ASAP7_75t_L g220 ( 
.A(n_137),
.B(n_72),
.Y(n_220)
);

A2O1A1Ixp33_ASAP7_75t_L g272 ( 
.A1(n_220),
.A2(n_174),
.B(n_163),
.C(n_143),
.Y(n_272)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_175),
.Y(n_221)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_221),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_119),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_152),
.B(n_11),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_223),
.B(n_235),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_224),
.A2(n_176),
.B1(n_171),
.B2(n_184),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_154),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_225),
.B(n_232),
.Y(n_260)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_156),
.Y(n_228)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_228),
.Y(n_273)
);

AO22x2_ASAP7_75t_L g229 ( 
.A1(n_159),
.A2(n_72),
.B1(n_133),
.B2(n_134),
.Y(n_229)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_229),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_168),
.Y(n_230)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_230),
.Y(n_282)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_142),
.Y(n_231)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_231),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_177),
.Y(n_232)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_120),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_233),
.Y(n_276)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_173),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_234),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_123),
.B(n_145),
.Y(n_235)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_140),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_236),
.B(n_240),
.Y(n_280)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_132),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_144),
.Y(n_238)
);

NAND2xp33_ASAP7_75t_SL g239 ( 
.A(n_159),
.B(n_133),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_141),
.B(n_124),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_168),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_128),
.B(n_148),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_242),
.B(n_244),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_177),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_154),
.B(n_164),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_245),
.B(n_201),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_246),
.A2(n_247),
.B1(n_250),
.B2(n_254),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_224),
.A2(n_136),
.B1(n_169),
.B2(n_183),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_207),
.A2(n_183),
.B1(n_146),
.B2(n_169),
.Y(n_250)
);

AO21x1_ASAP7_75t_L g321 ( 
.A1(n_252),
.A2(n_272),
.B(n_232),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_200),
.A2(n_182),
.B1(n_144),
.B2(n_125),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_264),
.B(n_201),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_243),
.A2(n_125),
.B1(n_155),
.B2(n_182),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_265),
.A2(n_271),
.B1(n_286),
.B2(n_253),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_197),
.A2(n_155),
.B1(n_179),
.B2(n_164),
.Y(n_271)
);

OAI21xp33_ASAP7_75t_SL g297 ( 
.A1(n_278),
.A2(n_239),
.B(n_220),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_283),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_223),
.B(n_219),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_219),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_282),
.Y(n_291)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_291),
.Y(n_344)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_292),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_294),
.B(n_295),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_262),
.Y(n_295)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_258),
.Y(n_296)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_296),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_297),
.B(n_319),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_299),
.Y(n_333)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_289),
.Y(n_300)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_300),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_213),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_301),
.B(n_303),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_274),
.B(n_205),
.Y(n_302)
);

AOI21xp33_ASAP7_75t_L g353 ( 
.A1(n_302),
.A2(n_325),
.B(n_249),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_227),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_289),
.Y(n_304)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_304),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_305),
.A2(n_308),
.B1(n_309),
.B2(n_313),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_226),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_306),
.B(n_315),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_268),
.A2(n_198),
.B1(n_221),
.B2(n_190),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_307),
.A2(n_316),
.B(n_320),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_254),
.A2(n_186),
.B1(n_229),
.B2(n_216),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_277),
.A2(n_229),
.B1(n_187),
.B2(n_210),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_253),
.B(n_194),
.C(n_231),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_310),
.B(n_317),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_252),
.A2(n_186),
.B1(n_229),
.B2(n_236),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_311),
.A2(n_314),
.B1(n_324),
.B2(n_265),
.Y(n_328)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_251),
.Y(n_312)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_312),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_250),
.A2(n_208),
.B1(n_192),
.B2(n_218),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_277),
.A2(n_238),
.B1(n_196),
.B2(n_233),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_259),
.B(n_202),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_272),
.A2(n_217),
.B(n_189),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_275),
.B(n_280),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_260),
.Y(n_318)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_318),
.Y(n_349)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_251),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_255),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_321),
.A2(n_322),
.B(n_264),
.Y(n_342)
);

AO21x1_ASAP7_75t_L g322 ( 
.A1(n_278),
.A2(n_244),
.B(n_209),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_247),
.A2(n_188),
.B1(n_230),
.B2(n_246),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_323),
.A2(n_290),
.B1(n_281),
.B2(n_264),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_280),
.A2(n_230),
.B1(n_283),
.B2(n_274),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_287),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_311),
.A2(n_286),
.B1(n_263),
.B2(n_268),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_326),
.A2(n_342),
.B(n_346),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_328),
.A2(n_338),
.B1(n_340),
.B2(n_297),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_298),
.A2(n_271),
.B1(n_263),
.B2(n_287),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_331),
.A2(n_339),
.B1(n_343),
.B2(n_351),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_317),
.B(n_275),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_332),
.B(n_350),
.C(n_310),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_298),
.A2(n_263),
.B1(n_281),
.B2(n_276),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_323),
.A2(n_264),
.B1(n_257),
.B2(n_288),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_308),
.A2(n_276),
.B1(n_248),
.B2(n_273),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_321),
.A2(n_288),
.B(n_273),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_293),
.B(n_269),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_324),
.A2(n_248),
.B1(n_269),
.B2(n_258),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_353),
.B(n_299),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_354),
.B(n_350),
.Y(n_377)
);

AOI21xp33_ASAP7_75t_L g396 ( 
.A1(n_356),
.A2(n_373),
.B(n_302),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_346),
.B(n_322),
.Y(n_357)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_357),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_332),
.B(n_306),
.C(n_294),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_358),
.B(n_370),
.C(n_371),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_295),
.Y(n_359)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_359),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_349),
.B(n_320),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_360),
.B(n_363),
.Y(n_380)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_330),
.Y(n_361)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_361),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_341),
.A2(n_321),
.B(n_322),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_362),
.A2(n_368),
.B(n_327),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_348),
.B(n_301),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_364),
.A2(n_357),
.B1(n_339),
.B2(n_368),
.Y(n_382)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_330),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_365),
.B(n_369),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_342),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_367),
.B(n_372),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_341),
.A2(n_316),
.B(n_307),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_348),
.B(n_303),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_337),
.B(n_292),
.C(n_291),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_337),
.B(n_315),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_347),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_352),
.B(n_319),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_328),
.A2(n_305),
.B1(n_309),
.B2(n_313),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_374),
.A2(n_376),
.B1(n_329),
.B2(n_351),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_352),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_375),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_331),
.A2(n_291),
.B1(n_314),
.B2(n_312),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_377),
.B(n_386),
.C(n_393),
.Y(n_397)
);

BUFx24_ASAP7_75t_SL g378 ( 
.A(n_369),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_378),
.B(n_396),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_371),
.B(n_333),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_381),
.B(n_373),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_382),
.A2(n_362),
.B1(n_357),
.B2(n_376),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_383),
.A2(n_388),
.B(n_366),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_384),
.A2(n_387),
.B1(n_390),
.B2(n_364),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_370),
.B(n_333),
.C(n_327),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_355),
.A2(n_338),
.B1(n_340),
.B2(n_327),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_355),
.A2(n_326),
.B1(n_344),
.B2(n_345),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_376),
.A2(n_343),
.B1(n_345),
.B2(n_336),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_370),
.B(n_336),
.C(n_335),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_385),
.B(n_354),
.C(n_371),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_398),
.B(n_401),
.C(n_403),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_399),
.A2(n_408),
.B1(n_395),
.B2(n_390),
.Y(n_418)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_389),
.Y(n_400)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_400),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_385),
.B(n_354),
.C(n_358),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_377),
.B(n_358),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_402),
.B(n_407),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_393),
.B(n_386),
.C(n_381),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_404),
.A2(n_405),
.B1(n_406),
.B2(n_399),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_384),
.A2(n_364),
.B1(n_375),
.B2(n_357),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_387),
.A2(n_362),
.B1(n_356),
.B2(n_363),
.Y(n_406)
);

INVxp33_ASAP7_75t_SL g407 ( 
.A(n_391),
.Y(n_407)
);

CKINVDCx14_ASAP7_75t_R g408 ( 
.A(n_380),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_383),
.A2(n_366),
.B(n_360),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_409),
.A2(n_410),
.B(n_388),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_412),
.B(n_392),
.C(n_372),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_416),
.B(n_417),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_418),
.A2(n_374),
.B1(n_410),
.B2(n_344),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_419),
.A2(n_409),
.B1(n_404),
.B2(n_405),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_397),
.B(n_379),
.C(n_389),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_420),
.B(n_422),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_400),
.A2(n_380),
.B1(n_359),
.B2(n_379),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_421),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_397),
.B(n_394),
.C(n_365),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_398),
.B(n_394),
.C(n_361),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_423),
.B(n_422),
.C(n_403),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_401),
.B(n_335),
.C(n_334),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_424),
.B(n_412),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_427),
.A2(n_431),
.B1(n_433),
.B2(n_414),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_420),
.B(n_402),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_428),
.B(n_413),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_429),
.B(n_430),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_415),
.A2(n_411),
.B1(n_406),
.B2(n_374),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_417),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_432),
.B(n_296),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_435),
.B(n_438),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_434),
.B(n_423),
.Y(n_436)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_436),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_437),
.A2(n_258),
.B1(n_270),
.B2(n_256),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_429),
.B(n_413),
.C(n_334),
.Y(n_438)
);

OAI321xp33_ASAP7_75t_L g440 ( 
.A1(n_426),
.A2(n_411),
.A3(n_304),
.B1(n_300),
.B2(n_267),
.C(n_296),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_440),
.B(n_270),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_441),
.A2(n_425),
.B(n_427),
.Y(n_445)
);

A2O1A1Ixp33_ASAP7_75t_L g442 ( 
.A1(n_426),
.A2(n_249),
.B(n_266),
.C(n_267),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_442),
.A2(n_256),
.B(n_266),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_439),
.A2(n_433),
.B1(n_425),
.B2(n_428),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_443),
.B(n_445),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_446),
.B(n_448),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_449),
.B(n_442),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_447),
.B(n_438),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_450),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_451),
.Y(n_454)
);

OAI32xp33_ASAP7_75t_L g455 ( 
.A1(n_453),
.A2(n_444),
.A3(n_449),
.B1(n_261),
.B2(n_285),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_455),
.A2(n_261),
.B(n_285),
.Y(n_458)
);

OAI21xp33_ASAP7_75t_L g457 ( 
.A1(n_456),
.A2(n_452),
.B(n_451),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_457),
.Y(n_459)
);

BUFx24_ASAP7_75t_SL g460 ( 
.A(n_459),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_460),
.B(n_454),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_461),
.B(n_458),
.Y(n_462)
);


endmodule