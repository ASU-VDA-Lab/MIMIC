module real_aes_8802_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_756;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g548 ( .A1(n_0), .A2(n_174), .B(n_549), .C(n_552), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_1), .B(n_499), .Y(n_553) );
INVx1_ASAP7_75t_L g108 ( .A(n_2), .Y(n_108) );
INVx1_ASAP7_75t_L g186 ( .A(n_3), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_4), .B(n_146), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_5), .A2(n_472), .B(n_493), .Y(n_492) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_6), .A2(n_166), .B(n_502), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_7), .A2(n_38), .B1(n_140), .B2(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_8), .B(n_166), .Y(n_175) );
AND2x6_ASAP7_75t_L g158 ( .A(n_9), .B(n_159), .Y(n_158) );
A2O1A1Ixp33_ASAP7_75t_L g561 ( .A1(n_10), .A2(n_158), .B(n_477), .C(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_11), .B(n_114), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_11), .B(n_39), .Y(n_434) );
INVx1_ASAP7_75t_L g136 ( .A(n_12), .Y(n_136) );
INVx1_ASAP7_75t_L g179 ( .A(n_13), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_14), .B(n_144), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_15), .B(n_146), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_16), .B(n_132), .Y(n_250) );
AO32x2_ASAP7_75t_L g192 ( .A1(n_17), .A2(n_131), .A3(n_157), .B1(n_166), .B2(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_18), .B(n_140), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_19), .B(n_132), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_20), .A2(n_55), .B1(n_140), .B2(n_195), .Y(n_196) );
AOI22xp33_ASAP7_75t_SL g234 ( .A1(n_21), .A2(n_82), .B1(n_140), .B2(n_144), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_22), .B(n_140), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_23), .A2(n_157), .B(n_477), .C(n_526), .Y(n_525) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_24), .A2(n_61), .B1(n_122), .B2(n_123), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_24), .Y(n_122) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_25), .A2(n_157), .B(n_477), .C(n_505), .Y(n_504) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_26), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_27), .B(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_28), .B(n_439), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_29), .A2(n_472), .B(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_30), .B(n_161), .Y(n_209) );
INVx2_ASAP7_75t_L g142 ( .A(n_31), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_32), .A2(n_475), .B(n_485), .C(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_33), .B(n_140), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_34), .B(n_161), .Y(n_220) );
XNOR2x2_ASAP7_75t_SL g119 ( .A(n_35), .B(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_36), .B(n_216), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g453 ( .A1(n_37), .A2(n_86), .B1(n_454), .B2(n_455), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_37), .Y(n_454) );
INVx1_ASAP7_75t_L g114 ( .A(n_39), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_40), .B(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_41), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_42), .B(n_146), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_43), .B(n_472), .Y(n_503) );
A2O1A1Ixp33_ASAP7_75t_L g474 ( .A1(n_44), .A2(n_475), .B(n_479), .C(n_485), .Y(n_474) );
OAI321xp33_ASAP7_75t_L g118 ( .A1(n_45), .A2(n_119), .A3(n_428), .B1(n_435), .B2(n_436), .C(n_438), .Y(n_118) );
INVx1_ASAP7_75t_L g435 ( .A(n_45), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_46), .A2(n_105), .B1(n_115), .B2(n_768), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_47), .B(n_140), .Y(n_169) );
INVx1_ASAP7_75t_L g550 ( .A(n_48), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_49), .A2(n_92), .B1(n_195), .B2(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g480 ( .A(n_50), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_51), .B(n_140), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_52), .B(n_140), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_53), .B(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_54), .B(n_152), .Y(n_173) );
AOI22xp33_ASAP7_75t_SL g248 ( .A1(n_56), .A2(n_62), .B1(n_140), .B2(n_144), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_57), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_58), .B(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_59), .B(n_140), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_60), .B(n_140), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_61), .Y(n_123) );
OAI22xp5_ASAP7_75t_SL g460 ( .A1(n_61), .A2(n_123), .B1(n_124), .B2(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g159 ( .A(n_63), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_64), .B(n_472), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_65), .B(n_499), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_66), .A2(n_152), .B(n_182), .C(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_67), .B(n_140), .Y(n_187) );
INVx1_ASAP7_75t_L g135 ( .A(n_68), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_69), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_70), .B(n_146), .Y(n_517) );
AO32x2_ASAP7_75t_L g230 ( .A1(n_71), .A2(n_157), .A3(n_166), .B1(n_231), .B2(n_235), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_72), .B(n_147), .Y(n_563) );
INVx1_ASAP7_75t_L g150 ( .A(n_73), .Y(n_150) );
INVx1_ASAP7_75t_L g204 ( .A(n_74), .Y(n_204) );
CKINVDCx16_ASAP7_75t_R g547 ( .A(n_75), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_76), .B(n_482), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g536 ( .A1(n_77), .A2(n_477), .B(n_485), .C(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_78), .B(n_144), .Y(n_205) );
CKINVDCx16_ASAP7_75t_R g494 ( .A(n_79), .Y(n_494) );
INVx1_ASAP7_75t_L g112 ( .A(n_80), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_81), .B(n_481), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_83), .B(n_195), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_84), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_85), .B(n_144), .Y(n_208) );
INVx1_ASAP7_75t_L g455 ( .A(n_86), .Y(n_455) );
INVx2_ASAP7_75t_L g133 ( .A(n_87), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_88), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_89), .B(n_156), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_90), .B(n_144), .Y(n_170) );
INVx2_ASAP7_75t_L g109 ( .A(n_91), .Y(n_109) );
OR2x2_ASAP7_75t_L g431 ( .A(n_91), .B(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g459 ( .A(n_91), .B(n_433), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_93), .A2(n_103), .B1(n_144), .B2(n_145), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_94), .B(n_472), .Y(n_513) );
INVx1_ASAP7_75t_L g516 ( .A(n_95), .Y(n_516) );
INVxp67_ASAP7_75t_L g497 ( .A(n_96), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_97), .B(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_98), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g538 ( .A(n_99), .Y(n_538) );
INVx1_ASAP7_75t_L g559 ( .A(n_100), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_101), .A2(n_451), .B1(n_452), .B2(n_453), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_101), .Y(n_451) );
AND2x2_ASAP7_75t_L g487 ( .A(n_102), .B(n_161), .Y(n_487) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
HB1xp67_ASAP7_75t_L g768 ( .A(n_106), .Y(n_768) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_113), .Y(n_106) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_108), .B(n_109), .C(n_110), .Y(n_107) );
AND2x2_ASAP7_75t_L g433 ( .A(n_108), .B(n_434), .Y(n_433) );
NOR2x2_ASAP7_75t_L g447 ( .A(n_109), .B(n_432), .Y(n_447) );
OR2x2_ASAP7_75t_L g464 ( .A(n_109), .B(n_433), .Y(n_464) );
OA211x2_ASAP7_75t_L g115 ( .A1(n_110), .A2(n_116), .B(n_118), .C(n_442), .Y(n_115) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g443 ( .A(n_117), .Y(n_443) );
NAND2x1p5_ASAP7_75t_L g436 ( .A(n_119), .B(n_437), .Y(n_436) );
XNOR2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_124), .Y(n_120) );
INVx1_ASAP7_75t_SL g461 ( .A(n_124), .Y(n_461) );
OR3x1_ASAP7_75t_L g124 ( .A(n_125), .B(n_356), .C(n_405), .Y(n_124) );
NAND5xp2_ASAP7_75t_L g125 ( .A(n_126), .B(n_271), .C(n_299), .D(n_329), .E(n_343), .Y(n_125) );
AOI221xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_189), .B1(n_221), .B2(n_226), .C(n_237), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_128), .B(n_162), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_128), .B(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g251 ( .A(n_129), .Y(n_251) );
AND2x2_ASAP7_75t_L g259 ( .A(n_129), .B(n_165), .Y(n_259) );
AND2x2_ASAP7_75t_L g282 ( .A(n_129), .B(n_164), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_129), .B(n_176), .Y(n_297) );
OR2x2_ASAP7_75t_L g306 ( .A(n_129), .B(n_244), .Y(n_306) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_129), .Y(n_309) );
AND2x2_ASAP7_75t_L g417 ( .A(n_129), .B(n_244), .Y(n_417) );
OA21x2_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_137), .B(n_160), .Y(n_129) );
OA21x2_ASAP7_75t_L g176 ( .A1(n_130), .A2(n_177), .B(n_188), .Y(n_176) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_131), .B(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_132), .Y(n_166) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
AND2x2_ASAP7_75t_SL g161 ( .A(n_133), .B(n_134), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
OAI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_149), .B(n_157), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_143), .B(n_146), .Y(n_138) );
INVx3_ASAP7_75t_L g203 ( .A(n_140), .Y(n_203) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_140), .Y(n_540) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g195 ( .A(n_141), .Y(n_195) );
BUFx3_ASAP7_75t_L g233 ( .A(n_141), .Y(n_233) );
AND2x6_ASAP7_75t_L g477 ( .A(n_141), .B(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g145 ( .A(n_142), .Y(n_145) );
INVx1_ASAP7_75t_L g153 ( .A(n_142), .Y(n_153) );
INVx2_ASAP7_75t_L g180 ( .A(n_144), .Y(n_180) );
INVx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_146), .A2(n_169), .B(n_170), .Y(n_168) );
INVx2_ASAP7_75t_L g174 ( .A(n_146), .Y(n_174) );
O2A1O1Ixp5_ASAP7_75t_SL g202 ( .A1(n_146), .A2(n_203), .B(n_204), .C(n_205), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_146), .B(n_497), .Y(n_496) );
INVx5_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
OAI22xp5_ASAP7_75t_SL g231 ( .A1(n_147), .A2(n_156), .B1(n_232), .B2(n_234), .Y(n_231) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_148), .Y(n_156) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_148), .Y(n_184) );
INVx1_ASAP7_75t_L g216 ( .A(n_148), .Y(n_216) );
AND2x2_ASAP7_75t_L g473 ( .A(n_148), .B(n_153), .Y(n_473) );
INVx1_ASAP7_75t_L g478 ( .A(n_148), .Y(n_478) );
O2A1O1Ixp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_154), .C(n_155), .Y(n_149) );
O2A1O1Ixp33_ASAP7_75t_L g185 ( .A1(n_151), .A2(n_174), .B(n_186), .C(n_187), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_151), .A2(n_527), .B(n_528), .Y(n_526) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_155), .A2(n_218), .B(n_219), .Y(n_217) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
OAI22xp5_ASAP7_75t_L g193 ( .A1(n_156), .A2(n_174), .B1(n_194), .B2(n_196), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_156), .A2(n_174), .B1(n_247), .B2(n_248), .Y(n_246) );
INVx4_ASAP7_75t_L g551 ( .A(n_156), .Y(n_551) );
NAND3xp33_ASAP7_75t_L g270 ( .A(n_157), .B(n_245), .C(n_246), .Y(n_270) );
BUFx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
OAI21xp5_ASAP7_75t_L g167 ( .A1(n_158), .A2(n_168), .B(n_171), .Y(n_167) );
OAI21xp5_ASAP7_75t_L g177 ( .A1(n_158), .A2(n_178), .B(n_185), .Y(n_177) );
OAI21xp5_ASAP7_75t_L g201 ( .A1(n_158), .A2(n_202), .B(n_206), .Y(n_201) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_158), .A2(n_212), .B(n_217), .Y(n_211) );
AND2x4_ASAP7_75t_L g472 ( .A(n_158), .B(n_473), .Y(n_472) );
INVx4_ASAP7_75t_SL g486 ( .A(n_158), .Y(n_486) );
NAND2x1p5_ASAP7_75t_L g560 ( .A(n_158), .B(n_473), .Y(n_560) );
OA21x2_ASAP7_75t_L g200 ( .A1(n_161), .A2(n_201), .B(n_209), .Y(n_200) );
OA21x2_ASAP7_75t_L g210 ( .A1(n_161), .A2(n_211), .B(n_220), .Y(n_210) );
INVx2_ASAP7_75t_L g235 ( .A(n_161), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_161), .A2(n_471), .B(n_474), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_161), .A2(n_513), .B(n_514), .Y(n_512) );
INVx1_ASAP7_75t_L g532 ( .A(n_161), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_162), .B(n_309), .Y(n_365) );
INVx2_ASAP7_75t_SL g162 ( .A(n_163), .Y(n_162) );
OAI311xp33_ASAP7_75t_L g307 ( .A1(n_163), .A2(n_308), .A3(n_309), .B1(n_310), .C1(n_325), .Y(n_307) );
AND2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_176), .Y(n_163) );
AND2x2_ASAP7_75t_L g268 ( .A(n_164), .B(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g275 ( .A(n_164), .Y(n_275) );
AND2x2_ASAP7_75t_L g396 ( .A(n_164), .B(n_225), .Y(n_396) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_165), .B(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g252 ( .A(n_165), .B(n_176), .Y(n_252) );
AND2x2_ASAP7_75t_L g304 ( .A(n_165), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g318 ( .A(n_165), .B(n_251), .Y(n_318) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_175), .Y(n_165) );
INVx4_ASAP7_75t_L g245 ( .A(n_166), .Y(n_245) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_166), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_166), .A2(n_503), .B(n_504), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_174), .Y(n_171) );
INVx2_ASAP7_75t_L g225 ( .A(n_176), .Y(n_225) );
AND2x2_ASAP7_75t_L g267 ( .A(n_176), .B(n_251), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_181), .C(n_182), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_180), .A2(n_506), .B(n_507), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_180), .A2(n_563), .B(n_564), .Y(n_562) );
O2A1O1Ixp33_ASAP7_75t_L g537 ( .A1(n_182), .A2(n_538), .B(n_539), .C(n_540), .Y(n_537) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_183), .A2(n_207), .B(n_208), .Y(n_206) );
INVx4_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g482 ( .A(n_184), .Y(n_482) );
AND2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_197), .Y(n_189) );
OR2x2_ASAP7_75t_L g362 ( .A(n_190), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_190), .B(n_368), .Y(n_379) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_191), .B(n_375), .Y(n_374) );
BUFx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g236 ( .A(n_192), .Y(n_236) );
AND2x2_ASAP7_75t_L g303 ( .A(n_192), .B(n_230), .Y(n_303) );
AND2x2_ASAP7_75t_L g314 ( .A(n_192), .B(n_210), .Y(n_314) );
AND2x2_ASAP7_75t_L g323 ( .A(n_192), .B(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_197), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_197), .B(n_264), .Y(n_308) );
INVx2_ASAP7_75t_SL g197 ( .A(n_198), .Y(n_197) );
OR2x2_ASAP7_75t_L g295 ( .A(n_198), .B(n_254), .Y(n_295) );
OR2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_210), .Y(n_198) );
INVx2_ASAP7_75t_L g228 ( .A(n_199), .Y(n_228) );
AND2x2_ASAP7_75t_L g322 ( .A(n_199), .B(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g240 ( .A(n_200), .Y(n_240) );
OR2x2_ASAP7_75t_L g339 ( .A(n_200), .B(n_340), .Y(n_339) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_200), .Y(n_402) );
AND2x2_ASAP7_75t_L g241 ( .A(n_210), .B(n_236), .Y(n_241) );
INVx1_ASAP7_75t_L g262 ( .A(n_210), .Y(n_262) );
AND2x2_ASAP7_75t_L g283 ( .A(n_210), .B(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g324 ( .A(n_210), .Y(n_324) );
INVx1_ASAP7_75t_L g340 ( .A(n_210), .Y(n_340) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_210), .Y(n_415) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_215), .Y(n_212) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVxp67_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_223), .B(n_328), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g371 ( .A1(n_223), .A2(n_313), .B1(n_362), .B2(n_372), .Y(n_371) );
INVx1_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
OAI211xp5_ASAP7_75t_SL g405 ( .A1(n_224), .A2(n_406), .B(n_408), .C(n_426), .Y(n_405) );
INVx2_ASAP7_75t_L g258 ( .A(n_225), .Y(n_258) );
AND2x2_ASAP7_75t_L g316 ( .A(n_225), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g327 ( .A(n_225), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_226), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_229), .Y(n_226) );
AND2x2_ASAP7_75t_L g300 ( .A(n_227), .B(n_264), .Y(n_300) );
BUFx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g332 ( .A(n_228), .B(n_323), .Y(n_332) );
AND2x2_ASAP7_75t_L g351 ( .A(n_228), .B(n_265), .Y(n_351) );
AND2x4_ASAP7_75t_L g287 ( .A(n_229), .B(n_261), .Y(n_287) );
AND2x2_ASAP7_75t_L g425 ( .A(n_229), .B(n_401), .Y(n_425) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_236), .Y(n_229) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_230), .Y(n_254) );
INVx1_ASAP7_75t_L g265 ( .A(n_230), .Y(n_265) );
INVx1_ASAP7_75t_L g364 ( .A(n_230), .Y(n_364) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_233), .Y(n_484) );
INVx2_ASAP7_75t_L g552 ( .A(n_233), .Y(n_552) );
INVx1_ASAP7_75t_L g529 ( .A(n_235), .Y(n_529) );
OR2x2_ASAP7_75t_L g255 ( .A(n_236), .B(n_240), .Y(n_255) );
AND2x2_ASAP7_75t_L g264 ( .A(n_236), .B(n_265), .Y(n_264) );
NOR2xp67_ASAP7_75t_L g284 ( .A(n_236), .B(n_285), .Y(n_284) );
OAI221xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_242), .B1(n_253), .B2(n_256), .C(n_260), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_239), .A2(n_261), .B(n_263), .C(n_266), .Y(n_260) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
INVx1_ASAP7_75t_L g285 ( .A(n_240), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_240), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_SL g368 ( .A(n_240), .B(n_262), .Y(n_368) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_240), .Y(n_375) );
AND2x2_ASAP7_75t_L g293 ( .A(n_241), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g330 ( .A(n_241), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_252), .Y(n_242) );
INVx2_ASAP7_75t_L g321 ( .A(n_243), .Y(n_321) );
AOI222xp33_ASAP7_75t_L g370 ( .A1(n_243), .A2(n_254), .B1(n_371), .B2(n_373), .C1(n_374), .C2(n_376), .Y(n_370) );
AND2x2_ASAP7_75t_L g427 ( .A(n_243), .B(n_396), .Y(n_427) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_251), .Y(n_243) );
INVx1_ASAP7_75t_L g317 ( .A(n_244), .Y(n_317) );
AO21x1_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_246), .B(n_249), .Y(n_244) );
INVx3_ASAP7_75t_L g499 ( .A(n_245), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_245), .B(n_519), .Y(n_518) );
AO21x2_ASAP7_75t_L g534 ( .A1(n_245), .A2(n_535), .B(n_542), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_245), .B(n_543), .Y(n_542) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_245), .A2(n_558), .B(n_565), .Y(n_557) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x4_ASAP7_75t_L g269 ( .A(n_250), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g355 ( .A(n_252), .B(n_289), .Y(n_355) );
AOI21xp33_ASAP7_75t_L g366 ( .A1(n_253), .A2(n_367), .B(n_369), .Y(n_366) );
OR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
INVx2_ASAP7_75t_L g294 ( .A(n_254), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_254), .B(n_261), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_254), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_SL g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx3_ASAP7_75t_L g320 ( .A(n_258), .Y(n_320) );
OR2x2_ASAP7_75t_L g372 ( .A(n_258), .B(n_294), .Y(n_372) );
AND2x2_ASAP7_75t_L g288 ( .A(n_259), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g326 ( .A(n_259), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_259), .B(n_320), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_259), .B(n_316), .Y(n_342) );
AND2x2_ASAP7_75t_L g346 ( .A(n_259), .B(n_328), .Y(n_346) );
INVxp67_ASAP7_75t_L g278 ( .A(n_261), .Y(n_278) );
BUFx3_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_263), .A2(n_336), .B1(n_341), .B2(n_342), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_263), .B(n_368), .Y(n_398) );
INVx1_ASAP7_75t_SL g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g384 ( .A(n_264), .B(n_375), .Y(n_384) );
AND2x2_ASAP7_75t_L g413 ( .A(n_264), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g418 ( .A(n_264), .B(n_368), .Y(n_418) );
INVx1_ASAP7_75t_L g331 ( .A(n_265), .Y(n_331) );
BUFx2_ASAP7_75t_L g337 ( .A(n_265), .Y(n_337) );
INVx1_ASAP7_75t_L g422 ( .A(n_266), .Y(n_422) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
NAND2x1p5_ASAP7_75t_L g273 ( .A(n_267), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g298 ( .A(n_268), .Y(n_298) );
NOR2x1_ASAP7_75t_L g274 ( .A(n_269), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g281 ( .A(n_269), .B(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g290 ( .A(n_269), .Y(n_290) );
INVx3_ASAP7_75t_L g328 ( .A(n_269), .Y(n_328) );
OR2x2_ASAP7_75t_L g394 ( .A(n_269), .B(n_395), .Y(n_394) );
AOI211xp5_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_276), .B(n_279), .C(n_291), .Y(n_271) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_272), .A2(n_409), .B1(n_416), .B2(n_418), .C(n_419), .Y(n_408) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_280), .B(n_286), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_282), .B(n_320), .Y(n_334) );
AND2x2_ASAP7_75t_L g376 ( .A(n_282), .B(n_316), .Y(n_376) );
INVx1_ASAP7_75t_SL g389 ( .A(n_283), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_283), .B(n_337), .Y(n_392) );
INVx1_ASAP7_75t_L g410 ( .A(n_284), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
AOI221xp5_ASAP7_75t_L g377 ( .A1(n_288), .A2(n_378), .B1(n_380), .B2(n_384), .C(n_385), .Y(n_377) );
AND2x2_ASAP7_75t_L g404 ( .A(n_289), .B(n_396), .Y(n_404) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g388 ( .A(n_290), .Y(n_388) );
AOI21xp33_ASAP7_75t_SL g291 ( .A1(n_292), .A2(n_295), .B(n_296), .Y(n_291) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g359 ( .A(n_294), .B(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g345 ( .A(n_295), .Y(n_345) );
INVx1_ASAP7_75t_L g373 ( .A(n_296), .Y(n_373) );
OR2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
O2A1O1Ixp33_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_301), .B(n_304), .C(n_307), .Y(n_299) );
OAI31xp33_ASAP7_75t_L g426 ( .A1(n_300), .A2(n_338), .A3(n_425), .B(n_427), .Y(n_426) );
INVxp67_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g400 ( .A(n_303), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_SL g421 ( .A(n_303), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_305), .B(n_320), .Y(n_348) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g423 ( .A(n_306), .B(n_320), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_315), .B1(n_319), .B2(n_322), .Y(n_310) );
NAND2xp33_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_314), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g350 ( .A(n_314), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g353 ( .A(n_314), .B(n_337), .Y(n_353) );
AND2x2_ASAP7_75t_L g407 ( .A(n_314), .B(n_402), .Y(n_407) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
INVx1_ASAP7_75t_L g382 ( .A(n_318), .Y(n_382) );
NOR2xp67_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
OAI32xp33_ASAP7_75t_L g385 ( .A1(n_320), .A2(n_354), .A3(n_386), .B1(n_388), .B2(n_389), .Y(n_385) );
INVx1_ASAP7_75t_L g360 ( .A(n_323), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_323), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g383 ( .A(n_327), .Y(n_383) );
O2A1O1Ixp33_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_332), .B(n_333), .C(n_335), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_331), .B(n_368), .Y(n_367) );
AOI221xp5_ASAP7_75t_L g343 ( .A1(n_332), .A2(n_344), .B1(n_345), .B2(n_346), .C(n_347), .Y(n_343) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g344 ( .A(n_342), .Y(n_344) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_349), .B1(n_352), .B2(n_354), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND4xp25_ASAP7_75t_SL g409 ( .A(n_352), .B(n_410), .C(n_411), .D(n_412), .Y(n_409) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
NAND4xp25_ASAP7_75t_SL g356 ( .A(n_357), .B(n_370), .C(n_377), .D(n_390), .Y(n_356) );
O2A1O1Ixp33_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_361), .B(n_365), .C(n_366), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g387 ( .A(n_363), .Y(n_387) );
INVx2_ASAP7_75t_L g411 ( .A(n_368), .Y(n_411) );
OR2x2_ASAP7_75t_L g420 ( .A(n_375), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_393), .B(n_397), .Y(n_390) );
INVxp67_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g416 ( .A(n_396), .B(n_417), .Y(n_416) );
AOI21xp33_ASAP7_75t_SL g397 ( .A1(n_398), .A2(n_399), .B(n_403), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
CKINVDCx16_ASAP7_75t_R g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_422), .B1(n_423), .B2(n_424), .Y(n_419) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g437 ( .A(n_430), .Y(n_437) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_SL g441 ( .A(n_431), .Y(n_441) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NAND4xp25_ASAP7_75t_SL g442 ( .A(n_438), .B(n_443), .C(n_444), .D(n_448), .Y(n_442) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
INVx3_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_450), .B1(n_456), .B2(n_763), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_460), .B1(n_462), .B2(n_465), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g764 ( .A(n_458), .Y(n_764) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g765 ( .A(n_460), .Y(n_765) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g766 ( .A(n_463), .Y(n_766) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx4_ASAP7_75t_L g767 ( .A(n_465), .Y(n_767) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OR5x1_ASAP7_75t_L g466 ( .A(n_467), .B(n_636), .C(n_714), .D(n_738), .E(n_755), .Y(n_466) );
OAI211xp5_ASAP7_75t_SL g467 ( .A1(n_468), .A2(n_508), .B(n_554), .C(n_613), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_488), .Y(n_468) );
AND2x2_ASAP7_75t_L g567 ( .A(n_469), .B(n_490), .Y(n_567) );
INVx5_ASAP7_75t_SL g595 ( .A(n_469), .Y(n_595) );
AND2x2_ASAP7_75t_L g631 ( .A(n_469), .B(n_616), .Y(n_631) );
OR2x2_ASAP7_75t_L g670 ( .A(n_469), .B(n_489), .Y(n_670) );
OR2x2_ASAP7_75t_L g701 ( .A(n_469), .B(n_592), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_469), .B(n_605), .Y(n_737) );
AND2x2_ASAP7_75t_L g749 ( .A(n_469), .B(n_592), .Y(n_749) );
OR2x6_ASAP7_75t_L g469 ( .A(n_470), .B(n_487), .Y(n_469) );
BUFx2_ASAP7_75t_L g524 ( .A(n_472), .Y(n_524) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_476), .A2(n_486), .B(n_494), .C(n_495), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_SL g546 ( .A1(n_476), .A2(n_486), .B(n_547), .C(n_548), .Y(n_546) );
INVx5_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B(n_483), .C(n_484), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g515 ( .A1(n_481), .A2(n_484), .B(n_516), .C(n_517), .Y(n_515) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g748 ( .A(n_488), .B(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
OR2x2_ASAP7_75t_L g611 ( .A(n_489), .B(n_612), .Y(n_611) );
OR2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_500), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_490), .B(n_592), .Y(n_591) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_490), .Y(n_604) );
INVx3_ASAP7_75t_L g619 ( .A(n_490), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_490), .B(n_500), .Y(n_643) );
OR2x2_ASAP7_75t_L g652 ( .A(n_490), .B(n_595), .Y(n_652) );
AND2x2_ASAP7_75t_L g656 ( .A(n_490), .B(n_616), .Y(n_656) );
AND2x2_ASAP7_75t_L g662 ( .A(n_490), .B(n_663), .Y(n_662) );
INVxp67_ASAP7_75t_L g699 ( .A(n_490), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_490), .B(n_557), .Y(n_713) );
OA21x2_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_492), .B(n_498), .Y(n_490) );
OA21x2_ASAP7_75t_L g544 ( .A1(n_499), .A2(n_545), .B(n_553), .Y(n_544) );
OR2x2_ASAP7_75t_L g605 ( .A(n_500), .B(n_557), .Y(n_605) );
AND2x2_ASAP7_75t_L g616 ( .A(n_500), .B(n_592), .Y(n_616) );
AND2x2_ASAP7_75t_L g628 ( .A(n_500), .B(n_619), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_500), .B(n_557), .Y(n_651) );
INVx1_ASAP7_75t_SL g663 ( .A(n_500), .Y(n_663) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g556 ( .A(n_501), .B(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_501), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_520), .Y(n_509) );
AND2x2_ASAP7_75t_L g576 ( .A(n_510), .B(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_510), .B(n_533), .Y(n_580) );
AND2x2_ASAP7_75t_L g583 ( .A(n_510), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_510), .B(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g608 ( .A(n_510), .B(n_599), .Y(n_608) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_510), .Y(n_627) );
AND2x2_ASAP7_75t_L g648 ( .A(n_510), .B(n_649), .Y(n_648) );
OR2x2_ASAP7_75t_L g658 ( .A(n_510), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g704 ( .A(n_510), .B(n_587), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_510), .B(n_610), .Y(n_731) );
INVx5_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx2_ASAP7_75t_L g601 ( .A(n_511), .Y(n_601) );
AND2x2_ASAP7_75t_L g667 ( .A(n_511), .B(n_599), .Y(n_667) );
AND2x2_ASAP7_75t_L g751 ( .A(n_511), .B(n_619), .Y(n_751) );
OR2x6_ASAP7_75t_L g511 ( .A(n_512), .B(n_518), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_520), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g740 ( .A(n_520), .Y(n_740) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_533), .Y(n_520) );
AND2x2_ASAP7_75t_L g570 ( .A(n_521), .B(n_571), .Y(n_570) );
AND2x4_ASAP7_75t_L g579 ( .A(n_521), .B(n_577), .Y(n_579) );
INVx5_ASAP7_75t_L g587 ( .A(n_521), .Y(n_587) );
AND2x2_ASAP7_75t_L g610 ( .A(n_521), .B(n_544), .Y(n_610) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_521), .Y(n_647) );
OR2x6_ASAP7_75t_L g521 ( .A(n_522), .B(n_530), .Y(n_521) );
AOI21xp5_ASAP7_75t_SL g522 ( .A1(n_523), .A2(n_525), .B(n_529), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
INVx1_ASAP7_75t_L g688 ( .A(n_533), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_533), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g721 ( .A(n_533), .B(n_587), .Y(n_721) );
A2O1A1Ixp33_ASAP7_75t_L g750 ( .A1(n_533), .A2(n_644), .B(n_751), .C(n_752), .Y(n_750) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_544), .Y(n_533) );
BUFx2_ASAP7_75t_L g571 ( .A(n_534), .Y(n_571) );
INVx2_ASAP7_75t_L g575 ( .A(n_534), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_541), .Y(n_535) );
INVx2_ASAP7_75t_L g577 ( .A(n_544), .Y(n_577) );
AND2x2_ASAP7_75t_L g584 ( .A(n_544), .B(n_575), .Y(n_584) );
AND2x2_ASAP7_75t_L g675 ( .A(n_544), .B(n_587), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
AOI211x1_ASAP7_75t_SL g554 ( .A1(n_555), .A2(n_568), .B(n_581), .C(n_606), .Y(n_554) );
INVx1_ASAP7_75t_L g672 ( .A(n_555), .Y(n_672) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_567), .Y(n_555) );
INVx5_ASAP7_75t_SL g592 ( .A(n_557), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_557), .B(n_662), .Y(n_661) );
AOI311xp33_ASAP7_75t_L g680 ( .A1(n_557), .A2(n_681), .A3(n_683), .B(n_684), .C(n_690), .Y(n_680) );
A2O1A1Ixp33_ASAP7_75t_L g715 ( .A1(n_557), .A2(n_628), .B(n_716), .C(n_719), .Y(n_715) );
OAI21xp5_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_560), .B(n_561), .Y(n_558) );
INVxp67_ASAP7_75t_L g635 ( .A(n_567), .Y(n_635) );
NAND4xp25_ASAP7_75t_SL g568 ( .A(n_569), .B(n_572), .C(n_578), .D(n_580), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_569), .B(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g626 ( .A(n_570), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_576), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_573), .B(n_579), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_573), .B(n_586), .Y(n_706) );
BUFx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_574), .B(n_587), .Y(n_724) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g599 ( .A(n_575), .Y(n_599) );
INVxp67_ASAP7_75t_L g634 ( .A(n_576), .Y(n_634) );
AND2x4_ASAP7_75t_L g586 ( .A(n_577), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g660 ( .A(n_577), .B(n_599), .Y(n_660) );
INVx1_ASAP7_75t_L g687 ( .A(n_577), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_577), .B(n_674), .Y(n_734) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_578), .B(n_648), .Y(n_668) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_579), .B(n_601), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_579), .B(n_648), .Y(n_747) );
INVx1_ASAP7_75t_L g758 ( .A(n_580), .Y(n_758) );
A2O1A1Ixp33_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_585), .B(n_588), .C(n_596), .Y(n_581) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g600 ( .A(n_584), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g638 ( .A(n_584), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g620 ( .A(n_585), .Y(n_620) );
AND2x2_ASAP7_75t_L g597 ( .A(n_586), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_586), .B(n_648), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_586), .B(n_667), .Y(n_691) );
OR2x2_ASAP7_75t_L g607 ( .A(n_587), .B(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g639 ( .A(n_587), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_587), .B(n_599), .Y(n_654) );
AND2x2_ASAP7_75t_L g711 ( .A(n_587), .B(n_667), .Y(n_711) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_587), .Y(n_718) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_589), .A2(n_601), .B1(n_723), .B2(n_725), .C(n_728), .Y(n_722) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_593), .Y(n_589) );
INVx1_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g612 ( .A(n_592), .B(n_595), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_592), .B(n_662), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_592), .B(n_619), .Y(n_727) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g712 ( .A(n_594), .B(n_713), .Y(n_712) );
OR2x2_ASAP7_75t_L g726 ( .A(n_594), .B(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_595), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g623 ( .A(n_595), .B(n_616), .Y(n_623) );
AND2x2_ASAP7_75t_L g693 ( .A(n_595), .B(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_595), .B(n_642), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_595), .B(n_743), .Y(n_742) );
OAI21xp5_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_600), .B(n_602), .Y(n_596) );
INVx2_ASAP7_75t_L g629 ( .A(n_597), .Y(n_629) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g649 ( .A(n_599), .Y(n_649) );
OR2x2_ASAP7_75t_L g653 ( .A(n_601), .B(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g756 ( .A(n_601), .B(n_724), .Y(n_756) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
AOI21xp33_ASAP7_75t_SL g606 ( .A1(n_607), .A2(n_609), .B(n_611), .Y(n_606) );
INVx1_ASAP7_75t_L g760 ( .A(n_607), .Y(n_760) );
INVx2_ASAP7_75t_SL g674 ( .A(n_608), .Y(n_674) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
A2O1A1Ixp33_ASAP7_75t_L g755 ( .A1(n_611), .A2(n_692), .B(n_756), .C(n_757), .Y(n_755) );
OAI322xp33_ASAP7_75t_SL g624 ( .A1(n_612), .A2(n_625), .A3(n_628), .B1(n_629), .B2(n_630), .C1(n_632), .C2(n_635), .Y(n_624) );
INVx2_ASAP7_75t_L g644 ( .A(n_612), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_620), .B1(n_621), .B2(n_623), .C(n_624), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OAI22xp33_ASAP7_75t_SL g690 ( .A1(n_615), .A2(n_691), .B1(n_692), .B2(n_695), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_616), .B(n_619), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_616), .B(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g689 ( .A(n_618), .B(n_651), .Y(n_689) );
INVx1_ASAP7_75t_L g679 ( .A(n_619), .Y(n_679) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AOI21xp5_ASAP7_75t_L g732 ( .A1(n_623), .A2(n_733), .B(n_735), .Y(n_732) );
AOI21xp33_ASAP7_75t_L g657 ( .A1(n_625), .A2(n_658), .B(n_661), .Y(n_657) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NOR2xp67_ASAP7_75t_SL g686 ( .A(n_627), .B(n_687), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_627), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_SL g743 ( .A(n_628), .Y(n_743) );
INVx1_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND4xp25_ASAP7_75t_L g636 ( .A(n_637), .B(n_664), .C(n_680), .D(n_696), .Y(n_636) );
AOI211xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_640), .B(n_645), .C(n_657), .Y(n_637) );
INVx1_ASAP7_75t_L g729 ( .A(n_638), .Y(n_729) );
AND2x2_ASAP7_75t_L g677 ( .A(n_639), .B(n_660), .Y(n_677) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
INVx1_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_644), .B(n_679), .Y(n_678) );
OAI22xp33_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_650), .B1(n_653), .B2(n_655), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_647), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g695 ( .A(n_648), .Y(n_695) );
O2A1O1Ixp33_ASAP7_75t_L g709 ( .A1(n_648), .A2(n_687), .B(n_710), .C(n_712), .Y(n_709) );
OR2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVx1_ASAP7_75t_L g694 ( .A(n_651), .Y(n_694) );
INVx1_ASAP7_75t_L g754 ( .A(n_652), .Y(n_754) );
NAND2xp33_ASAP7_75t_SL g744 ( .A(n_653), .B(n_745), .Y(n_744) );
INVx1_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g683 ( .A(n_662), .Y(n_683) );
O2A1O1Ixp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_668), .B(n_669), .C(n_671), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .B1(n_676), .B2(n_678), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_674), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_679), .B(n_700), .Y(n_762) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AOI21xp33_ASAP7_75t_SL g684 ( .A1(n_685), .A2(n_688), .B(n_689), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_702), .B1(n_705), .B2(n_707), .C(n_709), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
INVx1_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVxp67_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_712), .A2(n_729), .B1(n_730), .B2(n_731), .Y(n_728) );
NAND3xp33_ASAP7_75t_SL g714 ( .A(n_715), .B(n_722), .C(n_732), .Y(n_714) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
CKINVDCx16_ASAP7_75t_R g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVxp67_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
OAI211xp5_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_740), .B(n_741), .C(n_750), .Y(n_738) );
INVx1_ASAP7_75t_L g759 ( .A(n_739), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_744), .B1(n_746), .B2(n_748), .Y(n_741) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
AOI22xp5_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_759), .B1(n_760), .B2(n_761), .Y(n_757) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
OAI22x1_ASAP7_75t_SL g763 ( .A1(n_764), .A2(n_765), .B1(n_766), .B2(n_767), .Y(n_763) );
endmodule