module real_jpeg_14300_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_33;
wire n_38;
wire n_50;
wire n_35;
wire n_29;
wire n_55;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_51;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_39;
wire n_36;
wire n_40;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_48;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

BUFx10_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g12 ( 
.A1(n_3),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_12)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_3),
.A2(n_15),
.B1(n_46),
.B2(n_48),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_4),
.A2(n_13),
.B1(n_16),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_5),
.A2(n_13),
.B1(n_16),
.B2(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_6),
.B(n_17),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_6),
.B(n_28),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_6),
.A2(n_20),
.B1(n_46),
.B2(n_48),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_6),
.A2(n_31),
.B(n_48),
.C(n_54),
.Y(n_53)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_33),
.Y(n_8)
);

AOI21xp5_ASAP7_75t_L g9 ( 
.A1(n_10),
.A2(n_23),
.B(n_32),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_11),
.B(n_21),
.Y(n_10)
);

AOI22xp5_ASAP7_75t_SL g11 ( 
.A1(n_12),
.A2(n_17),
.B1(n_18),
.B2(n_20),
.Y(n_11)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_12),
.A2(n_17),
.B1(n_18),
.B2(n_25),
.Y(n_24)
);

INVx3_ASAP7_75t_SL g16 ( 
.A(n_13),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_13),
.B(n_22),
.Y(n_21)
);

OA22x2_ASAP7_75t_L g29 ( 
.A1(n_13),
.A2(n_16),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

OAI21xp33_ASAP7_75t_L g54 ( 
.A1(n_16),
.A2(n_20),
.B(n_30),
.Y(n_54)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_19),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_27),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_24),
.B(n_27),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_28),
.A2(n_45),
.B1(n_49),
.B2(n_51),
.Y(n_44)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_30),
.A2(n_31),
.B1(n_46),
.B2(n_48),
.Y(n_50)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_55),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_42),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_36),
.B(n_42),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_52),
.B2(n_53),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);


endmodule