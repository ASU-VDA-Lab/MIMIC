module real_jpeg_29774_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_258;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_70;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_216;
wire n_167;
wire n_128;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_0),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_0),
.A2(n_29),
.B1(n_33),
.B2(n_36),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_0),
.A2(n_29),
.B1(n_80),
.B2(n_81),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_0),
.A2(n_29),
.B1(n_49),
.B2(n_50),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_1),
.B(n_36),
.Y(n_65)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_1),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_2),
.A2(n_49),
.B1(n_50),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_2),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_2),
.A2(n_27),
.B1(n_30),
.B2(n_59),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_2),
.A2(n_33),
.B1(n_36),
.B2(n_59),
.Y(n_120)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_3),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_4),
.A2(n_80),
.B1(n_81),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_4),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_4),
.A2(n_49),
.B1(n_50),
.B2(n_152),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_4),
.A2(n_27),
.B1(n_30),
.B2(n_152),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_4),
.A2(n_33),
.B1(n_36),
.B2(n_152),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_6),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_6),
.B(n_83),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_6),
.B(n_49),
.Y(n_191)
);

AOI21xp33_ASAP7_75t_L g195 ( 
.A1(n_6),
.A2(n_49),
.B(n_191),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_6),
.A2(n_27),
.B1(n_30),
.B2(n_150),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_6),
.A2(n_11),
.B(n_33),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_6),
.B(n_100),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_6),
.A2(n_64),
.B1(n_66),
.B2(n_239),
.Y(n_241)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_7),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_8),
.A2(n_49),
.B1(n_50),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_8),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_8),
.A2(n_27),
.B1(n_30),
.B2(n_57),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_8),
.A2(n_33),
.B1(n_36),
.B2(n_57),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_9),
.A2(n_80),
.B1(n_81),
.B2(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_9),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_9),
.A2(n_49),
.B1(n_50),
.B2(n_107),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_9),
.A2(n_27),
.B1(n_30),
.B2(n_107),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_9),
.A2(n_33),
.B1(n_36),
.B2(n_107),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_10),
.A2(n_80),
.B1(n_81),
.B2(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_10),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_10),
.A2(n_49),
.B1(n_50),
.B2(n_132),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_10),
.A2(n_27),
.B1(n_30),
.B2(n_132),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_10),
.A2(n_33),
.B1(n_36),
.B2(n_132),
.Y(n_231)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_12),
.A2(n_27),
.B1(n_30),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_12),
.A2(n_43),
.B1(n_80),
.B2(n_81),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_12),
.A2(n_33),
.B1(n_36),
.B2(n_43),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_12),
.A2(n_43),
.B1(n_49),
.B2(n_50),
.Y(n_102)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_15),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_134),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_133),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_110),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_20),
.B(n_110),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_89),
.B2(n_109),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_61),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_44),
.B(n_60),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_24),
.B(n_44),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_38),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_25),
.A2(n_40),
.B(n_199),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_26),
.Y(n_143)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_27),
.A2(n_30),
.B1(n_35),
.B2(n_37),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_27),
.A2(n_30),
.B1(n_48),
.B2(n_54),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g192 ( 
.A(n_27),
.B(n_47),
.Y(n_192)
);

A2O1A1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_27),
.A2(n_35),
.B(n_150),
.C(n_218),
.Y(n_217)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI32xp33_ASAP7_75t_L g189 ( 
.A1(n_30),
.A2(n_50),
.A3(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_31),
.B(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_32),
.A2(n_40),
.B1(n_72),
.B2(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_32),
.A2(n_38),
.B(n_98),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_32),
.A2(n_40),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_32),
.A2(n_40),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_32),
.A2(n_40),
.B1(n_198),
.B2(n_216),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_32),
.B(n_150),
.Y(n_237)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_32)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_36),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_42),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_40),
.A2(n_72),
.B(n_73),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_40),
.A2(n_73),
.B(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_53),
.B1(n_55),
.B2(n_58),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_45),
.B(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_45),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_45),
.A2(n_53),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_45),
.A2(n_53),
.B1(n_146),
.B2(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_45),
.A2(n_53),
.B1(n_176),
.B2(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_53),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_46)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_47),
.Y(n_190)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_49),
.A2(n_50),
.B1(n_78),
.B2(n_79),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_49),
.B(n_78),
.Y(n_164)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_50),
.A2(n_82),
.B1(n_149),
.B2(n_164),
.Y(n_163)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_52),
.Y(n_54)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_53),
.B(n_102),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_53),
.B(n_127),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_56),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_74),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_71),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_63),
.A2(n_75),
.B1(n_76),
.B2(n_88),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_63),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_63),
.A2(n_71),
.B1(n_88),
.B2(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_66),
.B(n_69),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_64),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_64),
.A2(n_120),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_64),
.A2(n_95),
.B(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_64),
.A2(n_68),
.B1(n_231),
.B2(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_93),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_65),
.A2(n_70),
.B(n_122),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_65),
.A2(n_96),
.B1(n_230),
.B2(n_232),
.Y(n_229)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx5_ASAP7_75t_SL g167 ( 
.A(n_67),
.Y(n_167)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_68),
.B(n_94),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_68),
.B(n_150),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_71),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_84),
.B(n_85),
.Y(n_76)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_77),
.A2(n_83),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_80),
.B(n_82),
.C(n_83),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_80),
.Y(n_82)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

HAxp5_ASAP7_75t_SL g149 ( 
.A(n_80),
.B(n_150),
.CON(n_149),
.SN(n_149)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_83),
.B(n_84),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_86),
.A2(n_105),
.B1(n_106),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_86),
.A2(n_105),
.B1(n_131),
.B2(n_157),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_89),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_99),
.C(n_103),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_97),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_91),
.B(n_97),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_92),
.A2(n_166),
.B(n_180),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_99),
.A2(n_103),
.B1(n_104),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_99),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_106),
.B(n_108),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.C(n_117),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_115),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_117),
.B(n_279),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_124),
.C(n_129),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_118),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_123),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_124),
.A2(n_129),
.B1(n_130),
.B2(n_272),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_124),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B(n_128),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_125),
.A2(n_160),
.B(n_161),
.Y(n_159)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_276),
.B(n_281),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_181),
.B(n_262),
.C(n_275),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_168),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_137),
.B(n_168),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_153),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_139),
.B(n_140),
.C(n_153),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.C(n_148),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_141),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_148),
.B(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_151),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_162),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_158),
.B2(n_159),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_155),
.B(n_159),
.C(n_162),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_165),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.C(n_174),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_169),
.A2(n_170),
.B1(n_257),
.B2(n_259),
.Y(n_256)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_174),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.C(n_179),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_179),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_261),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_254),
.B(n_260),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_209),
.B(n_253),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_200),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_185),
.B(n_200),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_193),
.C(n_196),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_186),
.A2(n_187),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_189),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_193),
.A2(n_194),
.B1(n_196),
.B2(n_197),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_205),
.B2(n_206),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_201),
.B(n_207),
.C(n_208),
.Y(n_255)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_247),
.B(n_252),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_227),
.B(n_246),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_219),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_212),
.B(n_219),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_213),
.A2(n_214),
.B1(n_217),
.B2(n_234),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_217),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_225),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_224),
.C(n_225),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_226),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_235),
.B(n_245),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_233),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_229),
.B(n_233),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_240),
.B(n_244),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_237),
.B(n_238),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_248),
.B(n_249),
.Y(n_252)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_255),
.B(n_256),
.Y(n_260)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_257),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_263),
.B(n_264),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_273),
.B2(n_274),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_270),
.C(n_274),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_273),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_277),
.B(n_278),
.Y(n_281)
);


endmodule