module fake_jpeg_13888_n_368 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_368);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_368;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_21),
.B(n_8),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_77),
.Y(n_98)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_49),
.Y(n_139)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_20),
.B(n_8),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_52),
.B(n_71),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_53),
.Y(n_131)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_54),
.Y(n_140)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_60),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_63),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_68),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_69),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_70),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_20),
.B(n_36),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

BUFx4f_ASAP7_75t_SL g141 ( 
.A(n_75),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g133 ( 
.A(n_76),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_79),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_84),
.Y(n_100)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_82),
.Y(n_114)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_16),
.Y(n_83)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_36),
.B(n_15),
.Y(n_84)
);

BUFx4f_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_85),
.Y(n_135)
);

AOI21xp33_ASAP7_75t_L g86 ( 
.A1(n_37),
.A2(n_7),
.B(n_14),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_86),
.B(n_0),
.C(n_1),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_16),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_87),
.B(n_88),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_89),
.B(n_92),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_93),
.Y(n_118)
);

CKINVDCx9p33_ASAP7_75t_R g91 ( 
.A(n_41),
.Y(n_91)
);

INVx2_ASAP7_75t_R g116 ( 
.A(n_91),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_17),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_17),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_95),
.Y(n_120)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_27),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_60),
.A2(n_61),
.B1(n_59),
.B2(n_53),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_103),
.A2(n_104),
.B1(n_113),
.B2(n_117),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_47),
.A2(n_32),
.B1(n_45),
.B2(n_31),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_52),
.A2(n_37),
.B1(n_43),
.B2(n_31),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_75),
.A2(n_43),
.B1(n_27),
.B2(n_23),
.Y(n_117)
);

CKINVDCx12_ASAP7_75t_R g122 ( 
.A(n_77),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_122),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_83),
.A2(n_26),
.B1(n_24),
.B2(n_18),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_129),
.A2(n_138),
.B1(n_34),
.B2(n_38),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_71),
.B(n_24),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_130),
.B(n_137),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_70),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_87),
.A2(n_26),
.B1(n_11),
.B2(n_15),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_88),
.B(n_10),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_144),
.B(n_145),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_89),
.B(n_4),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_92),
.B(n_4),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_12),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_116),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_101),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_151),
.B(n_152),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_97),
.Y(n_153)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_100),
.B(n_74),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_154),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_108),
.B(n_1),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_170),
.Y(n_191)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_161),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_139),
.A2(n_96),
.B1(n_85),
.B2(n_34),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_157),
.Y(n_210)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_158),
.Y(n_193)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_102),
.B(n_2),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_163),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_160),
.A2(n_150),
.B1(n_154),
.B2(n_159),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_114),
.Y(n_161)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_3),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_164),
.B(n_165),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_3),
.Y(n_165)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_167),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_123),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_171),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_124),
.B(n_11),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_121),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_106),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_173),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_119),
.Y(n_173)
);

AO22x1_ASAP7_75t_L g174 ( 
.A1(n_116),
.A2(n_34),
.B1(n_38),
.B2(n_11),
.Y(n_174)
);

O2A1O1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_174),
.A2(n_179),
.B(n_141),
.C(n_139),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_12),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_183),
.Y(n_203)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_107),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_176),
.Y(n_189)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_177),
.Y(n_215)
);

AO22x1_ASAP7_75t_L g179 ( 
.A1(n_109),
.A2(n_34),
.B1(n_38),
.B2(n_117),
.Y(n_179)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_133),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_180),
.Y(n_214)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_107),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_182),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_132),
.B(n_120),
.Y(n_183)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_110),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_185),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_98),
.B(n_118),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_186),
.B(n_187),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_123),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_129),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_160),
.Y(n_206)
);

AO21x2_ASAP7_75t_L g197 ( 
.A1(n_155),
.A2(n_104),
.B(n_136),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_197),
.A2(n_201),
.B1(n_168),
.B2(n_170),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_183),
.A2(n_128),
.B1(n_136),
.B2(n_140),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_216),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_179),
.A2(n_99),
.B(n_135),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_204),
.A2(n_180),
.B(n_173),
.Y(n_234)
);

OAI21xp33_ASAP7_75t_SL g233 ( 
.A1(n_206),
.A2(n_99),
.B(n_153),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_154),
.B(n_119),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_212),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_119),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_162),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_159),
.B(n_140),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_181),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_223),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_174),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_220),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_221),
.A2(n_233),
.B1(n_242),
.B2(n_217),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_168),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_191),
.B(n_184),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_229),
.Y(n_253)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_226),
.Y(n_248)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_227),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_228),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_163),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_230),
.A2(n_234),
.B(n_236),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_204),
.A2(n_179),
.B(n_174),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_231),
.A2(n_198),
.B(n_207),
.Y(n_257)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_235),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_163),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_SL g236 ( 
.A(n_196),
.B(n_141),
.C(n_178),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_211),
.B(n_212),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_238),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_199),
.B(n_218),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_190),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_240),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_167),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_198),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_241),
.A2(n_211),
.B1(n_196),
.B2(n_216),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_197),
.A2(n_166),
.B1(n_131),
.B2(n_111),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_243),
.A2(n_256),
.B1(n_237),
.B2(n_230),
.Y(n_272)
);

XNOR2x1_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_208),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_225),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_220),
.A2(n_197),
.B1(n_206),
.B2(n_210),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_246),
.A2(n_247),
.B1(n_252),
.B2(n_258),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_220),
.A2(n_197),
.B1(n_213),
.B2(n_200),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_241),
.A2(n_196),
.B1(n_213),
.B2(n_197),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_251),
.A2(n_257),
.B(n_259),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_222),
.A2(n_197),
.B1(n_221),
.B2(n_223),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_222),
.A2(n_194),
.B1(n_192),
.B2(n_205),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_234),
.A2(n_194),
.B(n_202),
.Y(n_259)
);

BUFx24_ASAP7_75t_SL g263 ( 
.A(n_244),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_263),
.B(n_265),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_192),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_262),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_271),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_252),
.A2(n_247),
.B1(n_246),
.B2(n_249),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_268),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_230),
.B(n_231),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_232),
.Y(n_270)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_270),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_262),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_276),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_278),
.C(n_279),
.Y(n_296)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_274),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_249),
.A2(n_224),
.B1(n_235),
.B2(n_229),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_255),
.Y(n_277)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_236),
.C(n_239),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_245),
.B(n_227),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_249),
.A2(n_242),
.B1(n_215),
.B2(n_232),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_254),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_281),
.B(n_248),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_270),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_284),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_269),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_274),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_285),
.B(n_288),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_244),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_261),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_294),
.C(n_297),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_261),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_255),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_283),
.A2(n_275),
.B1(n_264),
.B2(n_267),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_298),
.A2(n_301),
.B1(n_305),
.B2(n_306),
.Y(n_320)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_287),
.Y(n_299)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_283),
.A2(n_275),
.B1(n_264),
.B2(n_259),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_304),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_295),
.A2(n_260),
.B1(n_280),
.B2(n_256),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_295),
.A2(n_257),
.B1(n_253),
.B2(n_268),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_289),
.A2(n_251),
.B(n_253),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_306),
.A2(n_289),
.B(n_281),
.Y(n_317)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_286),
.Y(n_307)
);

NAND4xp25_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_290),
.C(n_293),
.D(n_189),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_243),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_297),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_294),
.B(n_248),
.Y(n_309)
);

XNOR2x1_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_310),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_193),
.C(n_202),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_193),
.C(n_209),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_296),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_314),
.B(n_316),
.Y(n_335)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_317),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_318),
.B(n_321),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_303),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_323),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_320),
.A2(n_322),
.B1(n_301),
.B2(n_312),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_300),
.B(n_293),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_298),
.A2(n_292),
.B1(n_226),
.B2(n_205),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_309),
.C(n_310),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_308),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_324),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_329),
.B(n_332),
.Y(n_344)
);

OAI21x1_ASAP7_75t_L g337 ( 
.A1(n_330),
.A2(n_325),
.B(n_316),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_331),
.B(n_320),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_305),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_315),
.Y(n_333)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_333),
.Y(n_340)
);

INVxp33_ASAP7_75t_L g334 ( 
.A(n_322),
.Y(n_334)
);

AOI21xp33_ASAP7_75t_L g341 ( 
.A1(n_334),
.A2(n_313),
.B(n_226),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_314),
.B(n_209),
.Y(n_336)
);

NOR2xp67_ASAP7_75t_L g342 ( 
.A(n_336),
.B(n_313),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_337),
.B(n_338),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_323),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_339),
.B(n_341),
.Y(n_348)
);

AOI31xp67_ASAP7_75t_L g347 ( 
.A1(n_342),
.A2(n_326),
.A3(n_327),
.B(n_331),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_335),
.B(n_195),
.C(n_189),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_343),
.B(n_346),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_327),
.A2(n_195),
.B(n_185),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_345),
.B(n_153),
.Y(n_352)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_333),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_347),
.B(n_344),
.C(n_345),
.Y(n_354)
);

AOI322xp5_ASAP7_75t_L g349 ( 
.A1(n_338),
.A2(n_334),
.A3(n_335),
.B1(n_176),
.B2(n_182),
.C1(n_171),
.C2(n_112),
.Y(n_349)
);

AOI31xp67_ASAP7_75t_L g359 ( 
.A1(n_349),
.A2(n_353),
.A3(n_141),
.B(n_110),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_352),
.B(n_340),
.Y(n_355)
);

NOR2xp67_ASAP7_75t_L g353 ( 
.A(n_343),
.B(n_177),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_354),
.A2(n_356),
.B1(n_349),
.B2(n_146),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_355),
.B(n_356),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_351),
.B(n_143),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_350),
.B(n_158),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_357),
.B(n_105),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_348),
.A2(n_131),
.B1(n_111),
.B2(n_112),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_358),
.B(n_359),
.C(n_142),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_360),
.Y(n_365)
);

A2O1A1O1Ixp25_ASAP7_75t_L g364 ( 
.A1(n_361),
.A2(n_363),
.B(n_38),
.C(n_105),
.D(n_148),
.Y(n_364)
);

BUFx12f_ASAP7_75t_SL g366 ( 
.A(n_364),
.Y(n_366)
);

OAI21xp33_ASAP7_75t_L g367 ( 
.A1(n_366),
.A2(n_362),
.B(n_365),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_367),
.Y(n_368)
);


endmodule