module real_jpeg_24027_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_176;
wire n_288;
wire n_300;
wire n_166;
wire n_221;
wire n_286;
wire n_292;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_299;
wire n_173;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_200;
wire n_164;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_285;
wire n_304;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_58;
wire n_52;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_295;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_1),
.A2(n_19),
.B1(n_20),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_1),
.A2(n_35),
.B1(n_57),
.B2(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_1),
.A2(n_35),
.B1(n_45),
.B2(n_47),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_40),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_2),
.A2(n_40),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_2),
.A2(n_40),
.B1(n_45),
.B2(n_47),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_2),
.A2(n_19),
.B1(n_20),
.B2(n_40),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_2),
.A2(n_62),
.B(n_190),
.C(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_2),
.B(n_63),
.Y(n_204)
);

O2A1O1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_2),
.A2(n_20),
.B(n_25),
.C(n_215),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_2),
.B(n_44),
.C(n_45),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_2),
.B(n_23),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_2),
.B(n_120),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_2),
.B(n_42),
.Y(n_260)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_4),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_4),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_4),
.A2(n_22),
.B1(n_67),
.B2(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_4),
.A2(n_22),
.B1(n_45),
.B2(n_47),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_7),
.A2(n_58),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_7),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_7),
.A2(n_19),
.B1(n_20),
.B2(n_133),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_133),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_7),
.A2(n_45),
.B1(n_47),
.B2(n_133),
.Y(n_244)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_11),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_11),
.Y(n_121)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_11),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_111),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_110),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_93),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_15),
.B(n_93),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_15),
.B(n_303),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_15),
.B(n_303),
.Y(n_304)
);

FAx1_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_53),
.CI(n_78),
.CON(n_15),
.SN(n_15)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_16),
.A2(n_17),
.B(n_36),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_36),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_23),
.B(n_31),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_18),
.A2(n_71),
.B(n_72),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_19),
.A2(n_20),
.B1(n_25),
.B2(n_30),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_19),
.A2(n_20),
.B1(n_61),
.B2(n_62),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

OAI21xp33_ASAP7_75t_L g190 ( 
.A1(n_20),
.A2(n_40),
.B(n_61),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_23),
.B(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_24),
.B(n_34),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_24),
.B(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_24),
.A2(n_32),
.B(n_100),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_24)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_27),
.A2(n_28),
.B1(n_43),
.B2(n_44),
.Y(n_51)
);

OAI21xp33_ASAP7_75t_L g215 ( 
.A1(n_27),
.A2(n_30),
.B(n_40),
.Y(n_215)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_28),
.B(n_232),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_31),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_31),
.B(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_32),
.B(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_48),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_37),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_38),
.A2(n_41),
.B(n_75),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_39),
.B(n_50),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_41),
.A2(n_49),
.B(n_86),
.Y(n_125)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_42),
.B(n_52),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_42),
.B(n_219),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_45),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_45),
.B(n_256),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVxp33_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_49),
.B(n_229),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_52),
.Y(n_49)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_50),
.B(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_68),
.B1(n_76),
.B2(n_77),
.Y(n_53)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_54),
.A2(n_76),
.B1(n_95),
.B2(n_108),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_54),
.B(n_70),
.C(n_73),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_64),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_55),
.B(n_155),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_56),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_56),
.B(n_63),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_58),
.Y(n_132)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_59),
.B(n_65),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_59),
.B(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_65),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_63),
.A2(n_103),
.B(n_106),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_63),
.B(n_131),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_64),
.B(n_130),
.Y(n_185)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_68),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_73),
.B2(n_74),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_71),
.B(n_101),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_72),
.B(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_72),
.B(n_183),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_73),
.A2(n_74),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_73),
.B(n_172),
.C(n_174),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_73),
.A2(n_74),
.B1(n_174),
.B2(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_84),
.B(n_88),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_79),
.A2(n_85),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_79),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_79),
.A2(n_88),
.B1(n_89),
.B2(n_140),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_79),
.B(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_79),
.A2(n_140),
.B1(n_214),
.B2(n_272),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B(n_83),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_80),
.B(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_80),
.A2(n_145),
.B(n_146),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_80),
.B(n_83),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_80),
.B(n_243),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_81),
.Y(n_193)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_81),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_84),
.B(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_85),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_87),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_87),
.B(n_218),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B(n_92),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_109),
.Y(n_93)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_102),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_99),
.B(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_107),
.B(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_301),
.B(n_304),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_164),
.B(n_300),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_156),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_115),
.B(n_156),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_138),
.C(n_141),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_116),
.B(n_138),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_126),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_117),
.B(n_127),
.C(n_135),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_125),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_118),
.B(n_125),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_119),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_123),
.A2(n_145),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_123),
.B(n_249),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_134),
.B2(n_135),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_132),
.Y(n_191)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_137),
.B(n_176),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_141),
.B(n_298),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_153),
.C(n_154),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_142),
.A2(n_143),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_151),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_151),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_147),
.B(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_147),
.B(n_242),
.Y(n_261)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_152),
.B(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_153),
.A2(n_154),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_153),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_154),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_163),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_161),
.B2(n_162),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_158),
.B(n_162),
.C(n_163),
.Y(n_303)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_295),
.B(n_299),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_207),
.B(n_281),
.C(n_294),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_195),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_167),
.B(n_195),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_180),
.B2(n_194),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_178),
.B2(n_179),
.Y(n_169)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_170),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_170),
.B(n_179),
.C(n_194),
.Y(n_282)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_172),
.A2(n_173),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

INVxp67_ASAP7_75t_SL g184 ( 
.A(n_177),
.Y(n_184)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_180),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_188),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_181)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_182),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_182),
.B(n_187),
.C(n_188),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_185),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_192),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_201),
.C(n_202),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_196),
.A2(n_197),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_202),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.C(n_205),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_212),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_205),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_206),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_280),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_223),
.B(n_279),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_220),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_210),
.B(n_220),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.C(n_216),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_211),
.B(n_277),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_213),
.B(n_216),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_214),
.Y(n_272)
);

INVxp33_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_274),
.B(n_278),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_265),
.B(n_273),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_246),
.B(n_264),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_233),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_227),
.B(n_233),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_228),
.A2(n_230),
.B1(n_231),
.B2(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_228),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_240),
.B2(n_245),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_236),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_239),
.C(n_245),
.Y(n_266)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_237),
.Y(n_239)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_240),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_244),
.B(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_253),
.B(n_263),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_251),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_248),
.B(n_251),
.Y(n_263)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_249),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_259),
.B(n_262),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_260),
.B(n_261),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_266),
.B(n_267),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_271),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_270),
.C(n_271),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_275),
.B(n_276),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_282),
.B(n_283),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_293),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_291),
.B2(n_292),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_292),
.C(n_293),
.Y(n_296)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_296),
.B(n_297),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);


endmodule