module fake_jpeg_15445_n_234 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_234);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_234;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_29),
.Y(n_39)
);

INVxp33_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_46),
.Y(n_73)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_18),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_51),
.Y(n_81)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

NAND3xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_0),
.C(n_1),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_50),
.A2(n_36),
.B(n_27),
.C(n_16),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_18),
.B(n_0),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_55),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_16),
.B(n_1),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_56),
.B(n_20),
.Y(n_78)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_59),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_32),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_61),
.Y(n_94)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_29),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_39),
.A2(n_34),
.B1(n_33),
.B2(n_36),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_63),
.A2(n_86),
.B1(n_92),
.B2(n_98),
.Y(n_102)
);

OR2x2_ASAP7_75t_SL g64 ( 
.A(n_50),
.B(n_24),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_64),
.A2(n_67),
.B(n_76),
.C(n_97),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_27),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_65),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_66),
.B(n_78),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_55),
.A2(n_24),
.B1(n_35),
.B2(n_20),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_71),
.A2(n_96),
.B1(n_8),
.B2(n_10),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_79),
.Y(n_126)
);

A2O1A1O1Ixp25_ASAP7_75t_L g76 ( 
.A1(n_38),
.A2(n_30),
.B(n_28),
.C(n_37),
.D(n_26),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_32),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_37),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_84),
.B(n_85),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_40),
.B(n_35),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_40),
.A2(n_30),
.B1(n_19),
.B2(n_28),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_22),
.C(n_31),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_88),
.B(n_91),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_47),
.B(n_30),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_52),
.A2(n_19),
.B1(n_28),
.B2(n_26),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_52),
.A2(n_26),
.B1(n_25),
.B2(n_31),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_54),
.A2(n_22),
.B1(n_5),
.B2(n_7),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_2),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_58),
.A2(n_2),
.B1(n_5),
.B2(n_7),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_76),
.A2(n_58),
.B1(n_9),
.B2(n_10),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_99),
.A2(n_103),
.B1(n_98),
.B2(n_88),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_11),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_105),
.Y(n_133)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_14),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_8),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_114),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_77),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_115),
.Y(n_141)
);

NOR2x1_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_67),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_109),
.B(n_122),
.Y(n_150)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_113),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_84),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_77),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_86),
.B1(n_92),
.B2(n_66),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_116),
.A2(n_80),
.B1(n_74),
.B2(n_69),
.Y(n_135)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_117),
.Y(n_142)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_118),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_94),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_120),
.Y(n_149)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_122),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_65),
.B(n_97),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_127),
.Y(n_147)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_128),
.Y(n_156)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_129),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_111),
.A2(n_69),
.B1(n_74),
.B2(n_83),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_97),
.B(n_83),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_132),
.A2(n_151),
.B(n_117),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_134),
.A2(n_135),
.B1(n_145),
.B2(n_155),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_80),
.C(n_90),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_153),
.Y(n_161)
);

AND2x6_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_75),
.Y(n_139)
);

BUFx12_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_146),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_100),
.A2(n_103),
.B1(n_127),
.B2(n_118),
.Y(n_145)
);

AND2x6_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_126),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_150),
.B(n_106),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_108),
.B(n_126),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_114),
.C(n_126),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_157),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_102),
.A2(n_116),
.B1(n_123),
.B2(n_110),
.Y(n_155)
);

AND2x6_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_110),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_123),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_163),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_152),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_166),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_102),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_169),
.C(n_180),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_112),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_113),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_170),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_104),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_171),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_154),
.A2(n_121),
.B1(n_124),
.B2(n_129),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_173),
.A2(n_176),
.B1(n_177),
.B2(n_179),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_147),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_175),
.A2(n_178),
.B(n_158),
.Y(n_196)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_148),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_141),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_138),
.B(n_147),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_137),
.C(n_150),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_185),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_165),
.A2(n_162),
.B(n_178),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_184),
.A2(n_191),
.B(n_196),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_146),
.C(n_132),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_135),
.C(n_157),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_190),
.B(n_192),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_170),
.A2(n_140),
.B(n_156),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_143),
.C(n_139),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_160),
.A2(n_143),
.B1(n_140),
.B2(n_131),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_194),
.A2(n_195),
.B1(n_173),
.B2(n_164),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_169),
.A2(n_142),
.B1(n_131),
.B2(n_133),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_197),
.A2(n_175),
.B(n_163),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_199),
.Y(n_215)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_183),
.C(n_197),
.Y(n_211)
);

A2O1A1O1Ixp25_ASAP7_75t_L g204 ( 
.A1(n_196),
.A2(n_172),
.B(n_174),
.C(n_171),
.D(n_167),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_204),
.A2(n_208),
.B(n_191),
.Y(n_213)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_205),
.A2(n_206),
.B(n_207),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_186),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_187),
.B(n_188),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_188),
.B(n_172),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_194),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_212),
.C(n_213),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_185),
.C(n_190),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_217),
.Y(n_219)
);

MAJx2_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_184),
.C(n_193),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_216),
.A2(n_202),
.B(n_172),
.Y(n_223)
);

NOR2x1_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_189),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_215),
.A2(n_217),
.B1(n_192),
.B2(n_214),
.Y(n_218)
);

A2O1A1Ixp33_ASAP7_75t_SL g226 ( 
.A1(n_218),
.A2(n_174),
.B(n_199),
.C(n_209),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_210),
.B(n_200),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_220),
.B(n_222),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_205),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_212),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_202),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_224),
.B(n_226),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_225),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_221),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_227),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_228),
.C(n_226),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_232),
.B(n_233),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_231),
.B(n_230),
.Y(n_233)
);


endmodule