module real_jpeg_31849_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_572;
wire n_405;
wire n_412;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_22),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_1),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_1),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_1),
.Y(n_150)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_1),
.Y(n_332)
);

AND2x4_ASAP7_75t_L g35 ( 
.A(n_2),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_2),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_2),
.B(n_137),
.Y(n_136)
);

AND2x4_ASAP7_75t_L g184 ( 
.A(n_2),
.B(n_185),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_2),
.B(n_150),
.Y(n_210)
);

AND2x4_ASAP7_75t_L g225 ( 
.A(n_2),
.B(n_226),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_2),
.B(n_384),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_2),
.B(n_425),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_3),
.B(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_4),
.B(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_4),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_4),
.B(n_220),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_4),
.B(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_4),
.B(n_214),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_4),
.B(n_469),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_4),
.B(n_507),
.Y(n_506)
);

NAND2x1_ASAP7_75t_L g540 ( 
.A(n_4),
.B(n_541),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_5),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_5),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_5),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_6),
.Y(n_77)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_6),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_7),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_8),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_8),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_8),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_8),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_8),
.B(n_380),
.Y(n_379)
);

NAND2x1_ASAP7_75t_L g442 ( 
.A(n_8),
.B(n_443),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_8),
.B(n_54),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_8),
.B(n_511),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_9),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_9),
.B(n_127),
.Y(n_126)
);

NAND2x1_ASAP7_75t_L g169 ( 
.A(n_9),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_9),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_9),
.B(n_262),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_9),
.B(n_265),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_9),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_9),
.B(n_394),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_10),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_10),
.B(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_10),
.B(n_135),
.Y(n_134)
);

NAND2x1_ASAP7_75t_SL g167 ( 
.A(n_10),
.B(n_168),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_10),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_10),
.B(n_402),
.Y(n_401)
);

AND2x2_ASAP7_75t_SL g434 ( 
.A(n_10),
.B(n_194),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_10),
.B(n_481),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_11),
.Y(n_246)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_12),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_13),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_13),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_13),
.B(n_116),
.Y(n_115)
);

NAND2xp33_ASAP7_75t_SL g291 ( 
.A(n_13),
.B(n_292),
.Y(n_291)
);

NAND2x1_ASAP7_75t_L g304 ( 
.A(n_13),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_13),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_13),
.B(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_14),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_15),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_15),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_15),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_15),
.B(n_180),
.Y(n_179)
);

AND2x4_ASAP7_75t_SL g288 ( 
.A(n_15),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_15),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_15),
.B(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_15),
.B(n_329),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_16),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_16),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_16),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_17),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_17),
.B(n_86),
.Y(n_85)
);

NAND2xp33_ASAP7_75t_SL g193 ( 
.A(n_17),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_17),
.B(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_17),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_17),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_17),
.B(n_318),
.Y(n_317)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_528),
.B(n_568),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_458),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_449),
.Y(n_25)
);

NAND3xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_249),
.C(n_361),
.Y(n_26)
);

NOR2x1_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_199),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_151),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g451 ( 
.A(n_29),
.B(n_151),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_78),
.C(n_102),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_31),
.A2(n_78),
.B1(n_79),
.B2(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_31),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_50),
.Y(n_31)
);

OAI21x1_ASAP7_75t_L g196 ( 
.A1(n_32),
.A2(n_197),
.B(n_198),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_45),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_34),
.A2(n_35),
.B1(n_478),
.B2(n_482),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_34),
.A2(n_35),
.B1(n_183),
.B2(n_184),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_34),
.B(n_65),
.C(n_480),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_34),
.B(n_184),
.C(n_436),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

MAJx2_ASAP7_75t_L g155 ( 
.A(n_35),
.B(n_40),
.C(n_45),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_35),
.B(n_40),
.C(n_45),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_38),
.Y(n_168)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_44),
.Y(n_471)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_48),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_49),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_62),
.B2(n_63),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_51),
.B(n_62),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_51),
.B(n_62),
.Y(n_198)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_57),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_53),
.B(n_57),
.Y(n_101)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx5_ASAP7_75t_L g508 ( 
.A(n_55),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_57),
.A2(n_58),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJx2_ASAP7_75t_L g386 ( 
.A(n_58),
.B(n_210),
.C(n_213),
.Y(n_386)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_61),
.Y(n_163)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_69),
.C(n_74),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_65),
.B1(n_74),
.B2(n_83),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_64),
.B(n_422),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_64),
.A2(n_65),
.B1(n_479),
.B2(n_480),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_64),
.B(n_136),
.C(n_424),
.Y(n_484)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_67),
.Y(n_191)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_67),
.Y(n_220)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_67),
.Y(n_289)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_67),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_68),
.Y(n_269)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_72),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_77),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_77),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_77),
.Y(n_382)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_84),
.C(n_101),
.Y(n_79)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_80),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

MAJx2_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_89),
.C(n_95),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_85),
.B(n_89),
.C(n_95),
.Y(n_255)
);

XNOR2x1_ASAP7_75t_L g349 ( 
.A(n_85),
.B(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XNOR2x1_ASAP7_75t_L g350 ( 
.A(n_89),
.B(n_95),
.Y(n_350)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_94),
.Y(n_215)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_99),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_100),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_101),
.B(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_102),
.B(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_132),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_114),
.B1(n_130),
.B2(n_131),
.Y(n_103)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_109),
.B(n_112),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_109),
.Y(n_113)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_108),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_108),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_108),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_111),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_112),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_113),
.Y(n_237)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_130),
.C(n_132),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_121),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_115),
.B(n_122),
.C(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_117),
.Y(n_513)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_120),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_120),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_120),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XNOR2x2_ASAP7_75t_L g390 ( 
.A(n_123),
.B(n_391),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_123),
.B(n_210),
.C(n_393),
.Y(n_445)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_139),
.C(n_146),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_133),
.B(n_258),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_134),
.A2(n_178),
.B1(n_179),
.B2(n_182),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_134),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_134),
.B(n_179),
.C(n_184),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_134),
.A2(n_136),
.B1(n_182),
.B2(n_271),
.Y(n_270)
);

INVx4_ASAP7_75t_SL g287 ( 
.A(n_135),
.Y(n_287)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_136),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_136),
.A2(n_271),
.B1(n_423),
.B2(n_424),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_136),
.B(n_404),
.C(n_436),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_138),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_139),
.A2(n_140),
.B1(n_146),
.B2(n_147),
.Y(n_258)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_173),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_153),
.B(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_153),
.B(n_202),
.Y(n_203)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_157),
.B(n_159),
.C(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_165),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_160),
.B(n_169),
.C(n_229),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx4f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_163),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_169),
.B2(n_172),
.Y(n_165)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_166),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_166),
.A2(n_167),
.B1(n_432),
.B2(n_433),
.Y(n_431)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_169),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_171),
.Y(n_227)
);

AO21x1_ASAP7_75t_L g200 ( 
.A1(n_173),
.A2(n_201),
.B(n_203),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_196),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_187),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_187),
.C(n_196),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_183),
.B2(n_184),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVxp67_ASAP7_75t_SL g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_183),
.A2(n_184),
.B1(n_224),
.B2(n_225),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_183),
.B(n_225),
.C(n_434),
.Y(n_561)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_192),
.B1(n_193),
.B2(n_195),
.Y(n_188)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_189),
.Y(n_195)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_192),
.B(n_195),
.C(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OAI21x1_ASAP7_75t_L g450 ( 
.A1(n_199),
.A2(n_451),
.B(n_452),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_204),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g452 ( 
.A(n_200),
.B(n_204),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_205),
.B(n_364),
.C(n_365),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_232),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_207),
.Y(n_364)
);

XNOR2x1_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_216),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_208),
.B(n_217),
.C(n_231),
.Y(n_370)
);

XNOR2x1_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_210),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_210),
.B(n_261),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_210),
.A2(n_211),
.B1(n_392),
.B2(n_393),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_211),
.B(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_212),
.A2(n_213),
.B1(n_468),
.B2(n_472),
.Y(n_467)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_213),
.B(n_466),
.C(n_472),
.Y(n_498)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_228),
.B1(n_230),
.B2(n_231),
.Y(n_216)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

XNOR2x1_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_224),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_219),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_221),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_223),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_224),
.A2(n_225),
.B1(n_383),
.B2(n_385),
.Y(n_564)
);

AOI31xp33_ASAP7_75t_L g571 ( 
.A1(n_224),
.A2(n_385),
.A3(n_424),
.B(n_572),
.Y(n_571)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_225),
.B(n_397),
.C(n_398),
.Y(n_396)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_228),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_229),
.B(n_432),
.C(n_486),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_232),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_233),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_236),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_238),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_239),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_243),
.B1(n_247),
.B2(n_248),
.Y(n_240)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_241),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_243),
.Y(n_248)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_245),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

BUFx5_ASAP7_75t_L g406 ( 
.A(n_246),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_247),
.B(n_374),
.C(n_375),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_248),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_275),
.B(n_360),
.Y(n_249)
);

NOR2xp67_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_272),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_251),
.B(n_272),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_256),
.C(n_259),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_252),
.B(n_356),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_256),
.A2(n_257),
.B1(n_259),
.B2(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_259),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_264),
.C(n_270),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_260),
.B(n_264),
.Y(n_352)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_270),
.B(n_352),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_271),
.B(n_400),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_354),
.B(n_359),
.Y(n_275)
);

OAI21x1_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_342),
.B(n_353),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_310),
.B(n_341),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_294),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_279),
.B(n_294),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_288),
.C(n_290),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_280),
.A2(n_281),
.B1(n_337),
.B2(n_338),
.Y(n_336)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_285),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_285),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_288),
.A2(n_290),
.B1(n_291),
.B2(n_339),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_288),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_289),
.Y(n_309)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_300),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_296),
.B(n_299),
.C(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_300),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_301),
.B(n_304),
.C(n_348),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_308),
.Y(n_303)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_308),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_334),
.B(n_340),
.Y(n_310)
);

AOI21xp33_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_323),
.B(n_333),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_320),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_313),
.B(n_320),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_317),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_314),
.B(n_317),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_328),
.Y(n_323)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_336),
.Y(n_340)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_345),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g353 ( 
.A(n_343),
.B(n_345),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_351),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_349),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_347),
.B(n_349),
.C(n_351),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_355),
.B(n_358),
.Y(n_354)
);

NOR2xp67_ASAP7_75t_L g359 ( 
.A(n_355),
.B(n_358),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_361),
.A2(n_450),
.B(n_453),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_366),
.B1(n_412),
.B2(n_415),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_363),
.B(n_367),
.Y(n_456)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_387),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_368),
.B(n_407),
.C(n_414),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_369),
.A2(n_370),
.B1(n_371),
.B2(n_372),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_369),
.B(n_373),
.C(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

XNOR2x2_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_376),
.Y(n_372)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_376),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_386),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_379),
.B1(n_383),
.B2(n_385),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_378),
.B(n_385),
.C(n_386),
.Y(n_447)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_383),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_383),
.B(n_442),
.Y(n_441)
);

MAJx2_ASAP7_75t_L g464 ( 
.A(n_385),
.B(n_442),
.C(n_444),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_388),
.A2(n_389),
.B1(n_407),
.B2(n_411),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g414 ( 
.A(n_388),
.Y(n_414)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_395),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_390),
.B(n_396),
.C(n_399),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_399),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_404),
.Y(n_400)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_401),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_401),
.B(n_500),
.Y(n_499)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_407),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_409),
.C(n_410),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_413),
.Y(n_455)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

NOR2xp67_ASAP7_75t_L g454 ( 
.A(n_416),
.B(n_455),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_416),
.B(n_455),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_419),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_417),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_438),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_420),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_428),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_421),
.B(n_430),
.C(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_424),
.B(n_530),
.Y(n_529)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx6_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_430),
.B1(n_435),
.B2(n_437),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_430),
.Y(n_429)
);

XOR2x2_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_434),
.Y(n_430)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_432),
.Y(n_433)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_434),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_434),
.A2(n_486),
.B1(n_549),
.B2(n_550),
.Y(n_548)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_435),
.Y(n_437)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_437),
.Y(n_474)
);

INVxp33_ASAP7_75t_SL g524 ( 
.A(n_438),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_448),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_447),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_440),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_441),
.A2(n_444),
.B1(n_445),
.B2(n_446),
.Y(n_440)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_441),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_445),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_447),
.Y(n_489)
);

INVxp33_ASAP7_75t_L g488 ( 
.A(n_448),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_454),
.A2(n_456),
.B(n_457),
.Y(n_453)
);

NAND2x1_ASAP7_75t_SL g458 ( 
.A(n_459),
.B(n_520),
.Y(n_458)
);

AOI21x1_ASAP7_75t_L g553 ( 
.A1(n_459),
.A2(n_554),
.B(n_555),
.Y(n_553)
);

NAND2x1_ASAP7_75t_SL g459 ( 
.A(n_460),
.B(n_491),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_L g555 ( 
.A(n_460),
.B(n_491),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_475),
.C(n_487),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_462),
.B(n_476),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_473),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_465),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_464),
.B(n_465),
.C(n_493),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_467),
.Y(n_465)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_468),
.Y(n_472)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_471),
.Y(n_470)
);

INVxp67_ASAP7_75t_SL g493 ( 
.A(n_473),
.Y(n_493)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g476 ( 
.A(n_477),
.B(n_483),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_477),
.B(n_484),
.C(n_485),
.Y(n_516)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_478),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_479),
.A2(n_480),
.B1(n_563),
.B2(n_564),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_480),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_480),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_485),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_487),
.B(n_522),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_489),
.C(n_490),
.Y(n_487)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_492),
.A2(n_494),
.B(n_517),
.Y(n_491)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_492),
.Y(n_519)
);

NAND2x1p5_ASAP7_75t_L g517 ( 
.A(n_494),
.B(n_518),
.Y(n_517)
);

XOR2x2_ASAP7_75t_SL g494 ( 
.A(n_495),
.B(n_516),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_495),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_496),
.A2(n_497),
.B1(n_501),
.B2(n_502),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_499),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_498),
.B(n_501),
.C(n_552),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_499),
.Y(n_552)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

AO22x1_ASAP7_75t_L g502 ( 
.A1(n_503),
.A2(n_504),
.B1(n_514),
.B2(n_515),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_505),
.A2(n_506),
.B1(n_509),
.B2(n_510),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_506),
.B(n_509),
.C(n_514),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_516),
.Y(n_533)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_519),
.B(n_533),
.C(n_534),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_521),
.B(n_523),
.Y(n_520)
);

NOR2xp67_ASAP7_75t_SL g554 ( 
.A(n_521),
.B(n_523),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_525),
.C(n_527),
.Y(n_523)
);

INVxp67_ASAP7_75t_SL g525 ( 
.A(n_526),
.Y(n_525)
);

NAND3xp33_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_553),
.C(n_556),
.Y(n_528)
);

AOI31xp33_ASAP7_75t_L g568 ( 
.A1(n_529),
.A2(n_556),
.A3(n_569),
.B(n_571),
.Y(n_568)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_535),
.Y(n_531)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_532),
.B(n_535),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_536),
.B(n_551),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_537),
.B(n_538),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_537),
.B(n_538),
.C(n_551),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_548),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_540),
.A2(n_545),
.B1(n_546),
.B2(n_547),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_540),
.Y(n_546)
);

INVx3_ASAP7_75t_SL g541 ( 
.A(n_542),
.Y(n_541)
);

INVx4_ASAP7_75t_SL g542 ( 
.A(n_543),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_545),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_545),
.B(n_546),
.C(n_548),
.Y(n_566)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_549),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_SL g556 ( 
.A(n_557),
.B(n_560),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_558),
.B(n_567),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_559),
.B(n_566),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_560),
.A2(n_561),
.B1(n_562),
.B2(n_565),
.Y(n_559)
);

CKINVDCx16_ASAP7_75t_R g560 ( 
.A(n_561),
.Y(n_560)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_562),
.Y(n_565)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_573),
.Y(n_572)
);


endmodule