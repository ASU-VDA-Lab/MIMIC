module fake_jpeg_31162_n_411 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_411);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_411;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_16),
.B(n_14),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_44),
.B(n_48),
.Y(n_89)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_49),
.Y(n_88)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_16),
.B(n_12),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_53),
.B(n_57),
.Y(n_97)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_25),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_61),
.Y(n_104)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_63),
.Y(n_114)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_68),
.B(n_74),
.Y(n_117)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_31),
.B(n_12),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_70),
.B(n_79),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_71),
.A2(n_15),
.B1(n_18),
.B2(n_3),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_25),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_29),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_75),
.B(n_76),
.Y(n_128)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_18),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_78),
.B(n_82),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

BUFx8_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_80),
.Y(n_100)
);

BUFx16f_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_81),
.Y(n_134)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_18),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_83),
.A2(n_41),
.B1(n_20),
.B2(n_37),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

NAND2xp33_ASAP7_75t_SL g131 ( 
.A(n_84),
.B(n_42),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_31),
.B(n_12),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_22),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_71),
.A2(n_41),
.B(n_28),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_92),
.Y(n_164)
);

AO22x1_ASAP7_75t_SL g95 ( 
.A1(n_50),
.A2(n_35),
.B1(n_33),
.B2(n_30),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_95),
.A2(n_73),
.B1(n_65),
.B2(n_66),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_46),
.A2(n_29),
.B1(n_31),
.B2(n_36),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_99),
.A2(n_120),
.B1(n_133),
.B2(n_83),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_106),
.B(n_6),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_58),
.A2(n_20),
.B1(n_37),
.B2(n_19),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_107),
.A2(n_121),
.B1(n_123),
.B2(n_125),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_81),
.B(n_36),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_80),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_52),
.A2(n_22),
.B1(n_23),
.B2(n_32),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_110),
.A2(n_72),
.B1(n_63),
.B2(n_77),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_69),
.B(n_19),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_124),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_55),
.A2(n_23),
.B1(n_32),
.B2(n_19),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_81),
.A2(n_20),
.B1(n_37),
.B2(n_35),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_51),
.A2(n_35),
.B1(n_33),
.B2(n_30),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_62),
.B(n_33),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_67),
.A2(n_30),
.B1(n_27),
.B2(n_17),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_47),
.A2(n_27),
.B1(n_17),
.B2(n_15),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_127),
.A2(n_130),
.B1(n_42),
.B2(n_7),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_54),
.A2(n_27),
.B1(n_17),
.B2(n_15),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_79),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_135),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_136),
.B(n_137),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_118),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_56),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_138),
.B(n_141),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_80),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_140),
.B(n_105),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_118),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_142),
.A2(n_151),
.B(n_171),
.Y(n_193)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_143),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_97),
.B(n_84),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_144),
.B(n_147),
.Y(n_192)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_145),
.Y(n_201)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_146),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_104),
.B(n_42),
.Y(n_147)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_148),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_149),
.A2(n_153),
.B1(n_159),
.B2(n_165),
.Y(n_194)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_150),
.Y(n_212)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_132),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_154),
.B(n_155),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_42),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_86),
.Y(n_156)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

INVx6_ASAP7_75t_SL g188 ( 
.A(n_157),
.Y(n_188)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

INVx13_ASAP7_75t_L g202 ( 
.A(n_158),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_92),
.A2(n_49),
.B1(n_2),
.B2(n_4),
.Y(n_159)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_160),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_93),
.Y(n_162)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_162),
.Y(n_209)
);

BUFx24_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

INVx13_ASAP7_75t_L g200 ( 
.A(n_163),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_133),
.A2(n_49),
.B1(n_4),
.B2(n_5),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_89),
.B(n_106),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_166),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_119),
.A2(n_0),
.B1(n_5),
.B2(n_6),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_167),
.A2(n_176),
.B1(n_179),
.B2(n_88),
.Y(n_197)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_91),
.Y(n_169)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_169),
.Y(n_211)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_170),
.Y(n_213)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_102),
.Y(n_172)
);

INVx13_ASAP7_75t_L g216 ( 
.A(n_172),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_131),
.A2(n_42),
.B1(n_7),
.B2(n_8),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_173),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_174),
.B(n_175),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_119),
.B(n_7),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_95),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_108),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_177),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_116),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_178),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_124),
.A2(n_42),
.B1(n_8),
.B2(n_9),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_90),
.B(n_94),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_180),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_113),
.A2(n_9),
.B1(n_129),
.B2(n_101),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_181),
.A2(n_88),
.B1(n_122),
.B2(n_114),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_161),
.A2(n_91),
.B1(n_95),
.B2(n_105),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_182),
.A2(n_184),
.B(n_126),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_161),
.A2(n_164),
.B1(n_151),
.B2(n_143),
.Y(n_184)
);

CKINVDCx12_ASAP7_75t_R g189 ( 
.A(n_163),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_189),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_139),
.B(n_90),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_203),
.C(n_167),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_197),
.A2(n_160),
.B1(n_169),
.B2(n_157),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_139),
.B(n_94),
.C(n_101),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_164),
.B(n_96),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_205),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_180),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_210),
.B(n_221),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_140),
.B(n_102),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_152),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_168),
.A2(n_103),
.B1(n_114),
.B2(n_111),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_215),
.A2(n_222),
.B1(n_88),
.B2(n_170),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_163),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_201),
.Y(n_223)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_223),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_182),
.A2(n_149),
.B1(n_159),
.B2(n_165),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_224),
.A2(n_228),
.B1(n_234),
.B2(n_251),
.Y(n_279)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_225),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_226),
.B(n_200),
.Y(n_282)
);

O2A1O1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_210),
.A2(n_176),
.B(n_142),
.C(n_178),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_227),
.A2(n_122),
.B(n_219),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_184),
.A2(n_151),
.B1(n_179),
.B2(n_93),
.Y(n_228)
);

OA21x2_ASAP7_75t_L g229 ( 
.A1(n_204),
.A2(n_163),
.B(n_145),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_244),
.Y(n_264)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_230),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_232),
.A2(n_237),
.B1(n_248),
.B2(n_221),
.Y(n_258)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_233),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_198),
.A2(n_172),
.B1(n_111),
.B2(n_126),
.Y(n_234)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_191),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_236),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_194),
.A2(n_150),
.B1(n_146),
.B2(n_162),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_220),
.A2(n_158),
.B(n_177),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_238),
.A2(n_252),
.B(n_242),
.Y(n_268)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_239),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_185),
.B(n_154),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_240),
.B(n_243),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_191),
.Y(n_241)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_241),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_242),
.A2(n_205),
.B(n_192),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_185),
.B(n_158),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_213),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_257),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_249),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_194),
.A2(n_103),
.B1(n_156),
.B2(n_135),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_207),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_207),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_213),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_198),
.A2(n_220),
.B1(n_193),
.B2(n_203),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_218),
.A2(n_158),
.B(n_148),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_253),
.A2(n_208),
.B1(n_186),
.B2(n_209),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_189),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_254),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_190),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_255),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_218),
.A2(n_122),
.B1(n_193),
.B2(n_197),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_256),
.A2(n_200),
.B1(n_211),
.B2(n_202),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_199),
.B(n_122),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_258),
.A2(n_272),
.B1(n_234),
.B2(n_229),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_195),
.C(n_214),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_262),
.B(n_271),
.C(n_282),
.Y(n_294)
);

A2O1A1Ixp33_ASAP7_75t_SL g302 ( 
.A1(n_266),
.A2(n_281),
.B(n_284),
.C(n_254),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_248),
.A2(n_187),
.B1(n_217),
.B2(n_188),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_267),
.A2(n_232),
.B1(n_237),
.B2(n_236),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_268),
.A2(n_229),
.B(n_238),
.Y(n_295)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_269),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_217),
.C(n_196),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_227),
.A2(n_188),
.B1(n_209),
.B2(n_208),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_231),
.B(n_196),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_277),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_276),
.A2(n_288),
.B1(n_239),
.B2(n_244),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_231),
.B(n_183),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_183),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_223),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_243),
.B(n_202),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_202),
.Y(n_301)
);

AOI22x1_ASAP7_75t_L g281 ( 
.A1(n_224),
.A2(n_186),
.B1(n_219),
.B2(n_211),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_269),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_289),
.B(n_300),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_292),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_235),
.Y(n_293)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_293),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_295),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_296),
.A2(n_279),
.B1(n_264),
.B2(n_281),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_262),
.B(n_228),
.C(n_255),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_297),
.B(n_299),
.Y(n_320)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_263),
.Y(n_298)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_298),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_252),
.C(n_250),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_305),
.Y(n_317)
);

AO22x2_ASAP7_75t_L g333 ( 
.A1(n_302),
.A2(n_295),
.B1(n_314),
.B2(n_296),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_285),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_303),
.B(n_307),
.Y(n_319)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_263),
.Y(n_304)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_304),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_277),
.B(n_225),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_259),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_306),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_278),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_308),
.A2(n_313),
.B1(n_258),
.B2(n_286),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_283),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_309),
.B(n_287),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_264),
.B(n_249),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_290),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_271),
.B(n_246),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_266),
.Y(n_326)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_259),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_312),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_279),
.A2(n_284),
.B1(n_281),
.B2(n_288),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_268),
.A2(n_245),
.B(n_233),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_314),
.A2(n_264),
.B(n_265),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_315),
.A2(n_336),
.B(n_310),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_316),
.B(n_324),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_318),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_303),
.A2(n_274),
.B1(n_261),
.B2(n_260),
.Y(n_325)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_325),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_326),
.B(n_332),
.Y(n_346)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_329),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_313),
.A2(n_287),
.B1(n_286),
.B2(n_261),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_330),
.B(n_333),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_297),
.B(n_275),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_331),
.B(n_291),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_293),
.B(n_275),
.Y(n_332)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_332),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_302),
.A2(n_270),
.B(n_283),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_327),
.B(n_301),
.Y(n_340)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_340),
.Y(n_365)
);

NAND3xp33_ASAP7_75t_L g341 ( 
.A(n_319),
.B(n_298),
.C(n_304),
.Y(n_341)
);

NOR2xp67_ASAP7_75t_L g368 ( 
.A(n_341),
.B(n_334),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_342),
.A2(n_350),
.B(n_333),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_320),
.B(n_294),
.C(n_299),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_343),
.B(n_344),
.C(n_348),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_320),
.B(n_294),
.C(n_311),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_346),
.B(n_354),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_335),
.Y(n_347)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_347),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_326),
.B(n_291),
.C(n_289),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_349),
.B(n_317),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_323),
.A2(n_302),
.B(n_292),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_318),
.Y(n_352)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_352),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_315),
.B(n_290),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_317),
.B(n_305),
.Y(n_356)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_356),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_343),
.B(n_323),
.C(n_330),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_360),
.B(n_369),
.C(n_348),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_361),
.A2(n_367),
.B1(n_368),
.B2(n_353),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_346),
.B(n_336),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_363),
.B(n_342),
.Y(n_375)
);

AOI221xp5_ASAP7_75t_L g376 ( 
.A1(n_364),
.A2(n_345),
.B1(n_333),
.B2(n_302),
.C(n_338),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_340),
.A2(n_328),
.B1(n_335),
.B2(n_337),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_344),
.B(n_333),
.C(n_337),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_347),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_370),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_356),
.B(n_334),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_371),
.B(n_340),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_372),
.B(n_377),
.Y(n_384)
);

AOI22x1_ASAP7_75t_SL g373 ( 
.A1(n_364),
.A2(n_333),
.B1(n_350),
.B2(n_354),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_373),
.A2(n_363),
.B1(n_365),
.B2(n_369),
.Y(n_383)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_374),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_375),
.B(n_376),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_358),
.B(n_351),
.C(n_345),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_378),
.B(n_379),
.Y(n_391)
);

OAI221xp5_ASAP7_75t_L g379 ( 
.A1(n_359),
.A2(n_339),
.B1(n_355),
.B2(n_328),
.C(n_352),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_361),
.B(n_309),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_380),
.A2(n_382),
.B1(n_365),
.B2(n_307),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_357),
.A2(n_308),
.B1(n_322),
.B2(n_321),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_383),
.B(n_387),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_385),
.B(n_386),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_373),
.A2(n_338),
.B1(n_367),
.B2(n_324),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_376),
.A2(n_360),
.B(n_371),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_381),
.B(n_358),
.C(n_362),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_389),
.B(n_392),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_381),
.B(n_362),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_391),
.B(n_366),
.Y(n_393)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_393),
.Y(n_404)
);

AO221x1_ASAP7_75t_L g395 ( 
.A1(n_388),
.A2(n_366),
.B1(n_312),
.B2(n_306),
.C(n_270),
.Y(n_395)
);

NAND3xp33_ASAP7_75t_SL g402 ( 
.A(n_395),
.B(n_387),
.C(n_302),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_241),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_398),
.B(n_399),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_384),
.B(n_241),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_397),
.Y(n_400)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_400),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_402),
.A2(n_390),
.B1(n_302),
.B2(n_394),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_396),
.A2(n_392),
.B(n_390),
.Y(n_403)
);

NOR2xp67_ASAP7_75t_SL g406 ( 
.A(n_403),
.B(n_383),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_405),
.B(n_406),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_407),
.B(n_393),
.C(n_389),
.Y(n_408)
);

OAI321xp33_ASAP7_75t_L g410 ( 
.A1(n_408),
.A2(n_216),
.A3(n_230),
.B1(n_401),
.B2(n_404),
.C(n_409),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_410),
.B(n_216),
.Y(n_411)
);


endmodule