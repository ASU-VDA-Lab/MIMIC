module fake_jpeg_9750_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx8_ASAP7_75t_SL g27 ( 
.A(n_14),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_36),
.B(n_26),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_23),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_0),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_39),
.C(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_28),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_55),
.Y(n_86)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_58),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_16),
.B1(n_21),
.B2(n_31),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_48),
.A2(n_57),
.B1(n_65),
.B2(n_31),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_16),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_40),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_52),
.B(n_46),
.Y(n_76)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_60),
.C(n_32),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_34),
.A2(n_16),
.B1(n_31),
.B2(n_28),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_26),
.Y(n_59)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NAND2x1_ASAP7_75t_SL g60 ( 
.A(n_41),
.B(n_24),
.Y(n_60)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_37),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_34),
.A2(n_31),
.B1(n_28),
.B2(n_18),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_18),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_45),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_40),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_71),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_42),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_75),
.Y(n_115)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_76),
.B(n_52),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_42),
.B1(n_35),
.B2(n_34),
.Y(n_77)
);

AO22x1_ASAP7_75t_SL g95 ( 
.A1(n_77),
.A2(n_82),
.B1(n_60),
.B2(n_64),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_79),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_81),
.A2(n_18),
.B1(n_37),
.B2(n_26),
.Y(n_113)
);

CKINVDCx6p67_ASAP7_75t_R g82 ( 
.A(n_64),
.Y(n_82)
);

INVxp33_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_42),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_41),
.Y(n_110)
);

CKINVDCx12_ASAP7_75t_R g84 ( 
.A(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_87),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_18),
.B1(n_34),
.B2(n_35),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_65),
.B1(n_35),
.B2(n_62),
.Y(n_102)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_62),
.B1(n_53),
.B2(n_35),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_94),
.A2(n_95),
.B1(n_102),
.B2(n_107),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_77),
.Y(n_125)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_98),
.Y(n_129)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_99),
.B(n_98),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_110),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_106),
.B(n_17),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_71),
.A2(n_60),
.B1(n_61),
.B2(n_45),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_78),
.A2(n_58),
.B1(n_47),
.B2(n_61),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_74),
.B1(n_66),
.B2(n_90),
.Y(n_142)
);

NOR2x1_ASAP7_75t_R g111 ( 
.A(n_70),
.B(n_29),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_111),
.A2(n_114),
.B(n_104),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_113),
.A2(n_64),
.B1(n_37),
.B2(n_72),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_68),
.A2(n_86),
.B(n_77),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_79),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_89),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_69),
.B(n_51),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_77),
.Y(n_124)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_119),
.B(n_132),
.Y(n_161)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_121),
.A2(n_134),
.B1(n_135),
.B2(n_99),
.Y(n_158)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_128),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_124),
.B(n_140),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_125),
.A2(n_130),
.B(n_144),
.Y(n_159)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_127),
.B(n_134),
.Y(n_147)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

OR2x2_ASAP7_75t_SL g130 ( 
.A(n_111),
.B(n_32),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_87),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_131),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_117),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_95),
.A2(n_37),
.B1(n_56),
.B2(n_66),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_136),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_92),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_75),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_138),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_139),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_56),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_94),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_143),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_142),
.A2(n_145),
.B1(n_64),
.B2(n_116),
.Y(n_162)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_95),
.A2(n_56),
.B1(n_67),
.B2(n_29),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_112),
.A2(n_67),
.B1(n_37),
.B2(n_22),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_146),
.A2(n_100),
.B1(n_92),
.B2(n_112),
.Y(n_168)
);

OAI22x1_ASAP7_75t_SL g149 ( 
.A1(n_122),
.A2(n_102),
.B1(n_114),
.B2(n_96),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_SL g198 ( 
.A(n_149),
.B(n_160),
.C(n_163),
.Y(n_198)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_151),
.B(n_156),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_103),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_167),
.Y(n_180)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_157),
.B(n_164),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_158),
.A2(n_41),
.B(n_38),
.Y(n_204)
);

NAND2xp33_ASAP7_75t_SL g160 ( 
.A(n_125),
.B(n_96),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_162),
.A2(n_101),
.B1(n_119),
.B2(n_142),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_97),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_139),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_106),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_174),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_118),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_128),
.A2(n_100),
.B1(n_32),
.B2(n_19),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_169),
.A2(n_176),
.B1(n_25),
.B2(n_19),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_104),
.Y(n_173)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_133),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_121),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_125),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_143),
.A2(n_101),
.B1(n_17),
.B2(n_19),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_161),
.B(n_127),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_178),
.B(n_190),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_179),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_154),
.Y(n_183)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_183),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_184),
.A2(n_197),
.B1(n_158),
.B2(n_176),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_185),
.A2(n_192),
.B(n_193),
.Y(n_229)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_177),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_196),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_150),
.B(n_124),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_189),
.A2(n_200),
.B(n_202),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_132),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_171),
.A2(n_122),
.B1(n_144),
.B2(n_130),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_191),
.A2(n_162),
.B1(n_163),
.B2(n_172),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_161),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_147),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_166),
.Y(n_194)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_194),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_136),
.Y(n_195)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_153),
.A2(n_123),
.B1(n_17),
.B2(n_25),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_148),
.B(n_123),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_199),
.B(n_203),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_147),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_148),
.B(n_25),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_204),
.A2(n_205),
.B(n_164),
.Y(n_225)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_207),
.A2(n_30),
.B1(n_24),
.B2(n_33),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_198),
.B(n_155),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_213),
.C(n_224),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_216),
.Y(n_239)
);

A2O1A1O1Ixp25_ASAP7_75t_L g211 ( 
.A1(n_198),
.A2(n_149),
.B(n_159),
.C(n_160),
.D(n_165),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_204),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_167),
.C(n_205),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_181),
.A2(n_151),
.B1(n_150),
.B2(n_163),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_215),
.A2(n_202),
.B1(n_196),
.B2(n_182),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_192),
.B(n_165),
.Y(n_216)
);

XOR2x1_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_159),
.Y(n_220)
);

XOR2x2_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_189),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_222),
.A2(n_227),
.B(n_179),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_187),
.B(n_172),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_223),
.B(n_228),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_180),
.B(n_80),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_225),
.A2(n_230),
.B(n_201),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_41),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_184),
.C(n_195),
.Y(n_238)
);

OAI21xp33_ASAP7_75t_L g227 ( 
.A1(n_185),
.A2(n_152),
.B(n_13),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_193),
.B(n_152),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_181),
.A2(n_22),
.B(n_20),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_201),
.A2(n_139),
.B1(n_20),
.B2(n_73),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_231),
.A2(n_200),
.B1(n_186),
.B2(n_197),
.Y(n_233)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_232),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_233),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_235),
.B(n_251),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_225),
.Y(n_236)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_236),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_238),
.Y(n_254)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_241),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_182),
.C(n_194),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_243),
.C(n_248),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_213),
.B(n_29),
.C(n_33),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_215),
.A2(n_20),
.B1(n_29),
.B2(n_33),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_244),
.A2(n_245),
.B1(n_210),
.B2(n_206),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_206),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_247),
.B(n_249),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_208),
.B(n_33),
.C(n_30),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_221),
.Y(n_249)
);

NOR3xp33_ASAP7_75t_SL g250 ( 
.A(n_220),
.B(n_8),
.C(n_15),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_252),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_229),
.A2(n_8),
.B(n_15),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_214),
.B(n_7),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_253),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_235),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

AOI322xp5_ASAP7_75t_L g281 ( 
.A1(n_260),
.A2(n_247),
.A3(n_230),
.B1(n_209),
.B2(n_243),
.C1(n_30),
.C2(n_24),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_226),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_268),
.C(n_234),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_236),
.A2(n_219),
.B1(n_207),
.B2(n_229),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_267),
.A2(n_212),
.B1(n_248),
.B2(n_244),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_211),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_266),
.A2(n_241),
.B(n_212),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_270),
.A2(n_271),
.B(n_6),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_257),
.A2(n_239),
.B(n_219),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_268),
.B(n_222),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_279),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_256),
.A2(n_221),
.B(n_246),
.Y(n_274)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_274),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_275),
.Y(n_286)
);

OA21x2_ASAP7_75t_SL g276 ( 
.A1(n_262),
.A2(n_250),
.B(n_251),
.Y(n_276)
);

AOI21x1_ASAP7_75t_L g285 ( 
.A1(n_276),
.A2(n_263),
.B(n_264),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_261),
.A2(n_217),
.B1(n_231),
.B2(n_218),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_281),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_234),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_280),
.C(n_282),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_254),
.C(n_267),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_254),
.C(n_259),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_278),
.B(n_262),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_284),
.B(n_293),
.Y(n_302)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_285),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_30),
.C(n_24),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_290),
.C(n_292),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_0),
.C(n_1),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_291),
.B(n_6),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_0),
.C(n_1),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_271),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_272),
.C(n_270),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_297),
.C(n_299),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_269),
.C(n_7),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_269),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_303),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_7),
.C(n_13),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_6),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_290),
.C(n_289),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_302),
.B(n_292),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_304),
.A2(n_305),
.B(n_12),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_300),
.A2(n_283),
.B(n_286),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_307),
.A2(n_308),
.B1(n_2),
.B2(n_3),
.Y(n_312)
);

OAI221xp5_ASAP7_75t_L g308 ( 
.A1(n_295),
.A2(n_14),
.B1(n_10),
.B2(n_12),
.C(n_5),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_12),
.C(n_14),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_309),
.A2(n_2),
.B(n_3),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_311),
.Y(n_314)
);

A2O1A1Ixp33_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_310),
.B(n_312),
.C(n_306),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_313),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_2),
.C(n_3),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_2),
.C(n_4),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_4),
.C(n_5),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_4),
.Y(n_320)
);


endmodule