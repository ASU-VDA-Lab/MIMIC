module fake_jpeg_30448_n_247 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_107;
wire n_39;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_27),
.B(n_0),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_58),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_26),
.B(n_16),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_55),
.Y(n_72)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_26),
.B(n_16),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_31),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_63),
.Y(n_88)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_28),
.B(n_0),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_62),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_29),
.B(n_1),
.Y(n_62)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_20),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_43),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_64),
.A2(n_41),
.B1(n_20),
.B2(n_24),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_80),
.B1(n_89),
.B2(n_44),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_48),
.A2(n_20),
.B1(n_18),
.B2(n_33),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_84),
.B1(n_21),
.B2(n_22),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_60),
.A2(n_20),
.B1(n_35),
.B2(n_30),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_57),
.B(n_32),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_81),
.B(n_23),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_58),
.A2(n_18),
.B1(n_33),
.B2(n_21),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_61),
.A2(n_24),
.B1(n_35),
.B2(n_30),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_32),
.Y(n_90)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_87),
.A2(n_45),
.B1(n_47),
.B2(n_53),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_94),
.A2(n_102),
.B1(n_83),
.B2(n_77),
.Y(n_126)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

INVx4_ASAP7_75t_SL g127 ( 
.A(n_96),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_99),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_74),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_100),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_66),
.B(n_62),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_105),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_52),
.B1(n_51),
.B2(n_59),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_103),
.A2(n_104),
.B1(n_106),
.B2(n_111),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_75),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_19),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_66),
.B(n_43),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_108),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_66),
.B(n_39),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_87),
.A2(n_54),
.B1(n_46),
.B2(n_42),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_109),
.A2(n_110),
.B1(n_115),
.B2(n_82),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_70),
.A2(n_63),
.B1(n_39),
.B2(n_38),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_112),
.A2(n_114),
.B1(n_116),
.B2(n_85),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_38),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_19),
.C(n_23),
.Y(n_132)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_50),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_126),
.B1(n_133),
.B2(n_123),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_67),
.C(n_78),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_115),
.C(n_97),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_98),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_136),
.C(n_129),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_128),
.A2(n_99),
.B(n_115),
.C(n_100),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_135),
.B(n_118),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_102),
.C(n_91),
.Y(n_136)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_121),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_140),
.A2(n_150),
.B1(n_79),
.B2(n_75),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_104),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_144),
.Y(n_153)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_133),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_120),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_86),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_116),
.B1(n_114),
.B2(n_69),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_146),
.A2(n_148),
.B1(n_93),
.B2(n_69),
.Y(n_162)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_131),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_149),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_133),
.A2(n_109),
.B1(n_83),
.B2(n_77),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_151),
.A2(n_158),
.B(n_163),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_65),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_166),
.Y(n_172)
);

AO22x1_ASAP7_75t_SL g156 ( 
.A1(n_143),
.A2(n_126),
.B1(n_117),
.B2(n_119),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_140),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_119),
.B(n_111),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_132),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_161),
.B(n_134),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_144),
.A2(n_119),
.B(n_112),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_79),
.B1(n_82),
.B2(n_86),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_145),
.B1(n_103),
.B2(n_95),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_147),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_135),
.A2(n_121),
.B(n_88),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_167),
.A2(n_137),
.B1(n_168),
.B2(n_157),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_178),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_179),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_171),
.A2(n_173),
.B1(n_156),
.B2(n_165),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_167),
.A2(n_150),
.B1(n_142),
.B2(n_136),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_177),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_139),
.Y(n_178)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_165),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_182),
.Y(n_186)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

XNOR2x1_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_151),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_188),
.B(n_177),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_181),
.A2(n_158),
.B(n_168),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_190),
.A2(n_180),
.B(n_171),
.Y(n_200)
);

OAI31xp33_ASAP7_75t_L g192 ( 
.A1(n_170),
.A2(n_153),
.A3(n_163),
.B(n_157),
.Y(n_192)
);

OAI21xp33_ASAP7_75t_L g199 ( 
.A1(n_192),
.A2(n_189),
.B(n_176),
.Y(n_199)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_184),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_195),
.A2(n_180),
.B1(n_173),
.B2(n_181),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_197),
.A2(n_207),
.B1(n_187),
.B2(n_160),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_186),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_198),
.B(n_200),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_199),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_184),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_201),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_196),
.B(n_172),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_202),
.A2(n_185),
.B1(n_193),
.B2(n_194),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_179),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_205),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_193),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_204),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_191),
.A2(n_156),
.B1(n_152),
.B2(n_166),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_206),
.A2(n_138),
.B1(n_96),
.B2(n_65),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_191),
.A2(n_160),
.B1(n_148),
.B2(n_106),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_213),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_197),
.A2(n_187),
.B1(n_192),
.B2(n_190),
.Y(n_216)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_216),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_217),
.A2(n_148),
.B(n_138),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_214),
.A2(n_199),
.B(n_203),
.Y(n_221)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_221),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_209),
.B(n_206),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_225),
.Y(n_226)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_218),
.Y(n_223)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_223),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_207),
.Y(n_224)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_224),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_210),
.C(n_211),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_3),
.Y(n_236)
);

XNOR2x1_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_210),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_230),
.A2(n_213),
.B1(n_224),
.B2(n_204),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_227),
.A2(n_231),
.B1(n_229),
.B2(n_226),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_233),
.Y(n_238)
);

OAI21x1_ASAP7_75t_SL g234 ( 
.A1(n_230),
.A2(n_217),
.B(n_2),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_234),
.A2(n_235),
.B(n_4),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_227),
.A2(n_1),
.B(n_2),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_236),
.B(n_4),
.C(n_5),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_237),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_239),
.B(n_236),
.Y(n_240)
);

NAND3xp33_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_5),
.C(n_7),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_238),
.C(n_6),
.Y(n_242)
);

AOI321xp33_ASAP7_75t_L g244 ( 
.A1(n_242),
.A2(n_243),
.A3(n_5),
.B1(n_7),
.B2(n_9),
.C(n_10),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_244),
.B(n_11),
.Y(n_245)
);

OAI321xp33_ASAP7_75t_L g246 ( 
.A1(n_245),
.A2(n_11),
.A3(n_12),
.B1(n_13),
.B2(n_43),
.C(n_240),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_11),
.Y(n_247)
);


endmodule