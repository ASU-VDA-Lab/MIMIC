module fake_jpeg_5756_n_77 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_4),
.B(n_7),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_22),
.Y(n_28)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_12),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_27),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_24),
.B(n_26),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_11),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_25),
.A2(n_16),
.B(n_19),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_1),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_19),
.Y(n_29)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_33),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_26),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_32),
.A2(n_27),
.B1(n_21),
.B2(n_22),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_10),
.B1(n_14),
.B2(n_18),
.Y(n_55)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_13),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_15),
.B(n_11),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_26),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_41),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_25),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_34),
.A2(n_27),
.B1(n_21),
.B2(n_25),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_31),
.B1(n_22),
.B2(n_21),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

O2A1O1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_25),
.B(n_22),
.C(n_27),
.Y(n_47)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_48),
.A2(n_55),
.B1(n_45),
.B2(n_44),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_13),
.C(n_12),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_40),
.C(n_37),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_56),
.B(n_58),
.Y(n_64)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_46),
.B1(n_36),
.B2(n_45),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_59),
.A2(n_52),
.B1(n_51),
.B2(n_50),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_39),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_55),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_57),
.Y(n_67)
);

NAND4xp25_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_44),
.C(n_54),
.D(n_53),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_63),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_66),
.C(n_60),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_68),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_66),
.A2(n_14),
.B1(n_18),
.B2(n_2),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_64),
.C(n_69),
.Y(n_71)
);

MAJx2_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_7),
.C(n_8),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_62),
.B(n_65),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_73),
.B(n_72),
.Y(n_74)
);

OAI21x1_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_75),
.B(n_8),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_9),
.Y(n_77)
);


endmodule