module fake_netlist_1_2011_n_309 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_309, n_686);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_309;
output n_686;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_357;
wire n_90;
wire n_245;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_522;
wire n_264;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_SL g78 ( .A(n_27), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_10), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_73), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_0), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_33), .Y(n_82) );
INVxp67_ASAP7_75t_L g83 ( .A(n_15), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_48), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_12), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_19), .Y(n_86) );
CKINVDCx14_ASAP7_75t_R g87 ( .A(n_20), .Y(n_87) );
BUFx6f_ASAP7_75t_L g88 ( .A(n_17), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_16), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_28), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_45), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_24), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_66), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_43), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_11), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_44), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_35), .Y(n_97) );
CKINVDCx16_ASAP7_75t_R g98 ( .A(n_36), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_14), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_18), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_0), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_59), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_68), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_57), .Y(n_104) );
INVx2_ASAP7_75t_SL g105 ( .A(n_23), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_52), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_42), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_41), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_22), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_53), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_58), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_13), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_47), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_10), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_55), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_12), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_72), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_39), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_4), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_25), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_9), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_5), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_2), .Y(n_123) );
INVxp67_ASAP7_75t_SL g124 ( .A(n_31), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_95), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_101), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g127 ( .A(n_78), .B(n_1), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_87), .B(n_1), .Y(n_128) );
INVx3_ASAP7_75t_L g129 ( .A(n_101), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_82), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_105), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_88), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_95), .B(n_2), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_86), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_90), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_87), .B(n_3), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_91), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_88), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_88), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_92), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_88), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_93), .Y(n_142) );
INVx1_ASAP7_75t_SL g143 ( .A(n_122), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_96), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_97), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_103), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_104), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_107), .Y(n_148) );
BUFx3_ASAP7_75t_L g149 ( .A(n_108), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_109), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_113), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_115), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_118), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_120), .Y(n_154) );
OAI22xp5_ASAP7_75t_SL g155 ( .A1(n_122), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_79), .Y(n_156) );
OAI22xp5_ASAP7_75t_SL g157 ( .A1(n_106), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_81), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_98), .B(n_6), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_85), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_99), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_112), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_114), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_83), .B(n_7), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_116), .Y(n_165) );
AND2x4_ASAP7_75t_L g166 ( .A(n_119), .B(n_8), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_121), .Y(n_167) );
INVx1_ASAP7_75t_SL g168 ( .A(n_106), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_131), .B(n_102), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_150), .Y(n_170) );
INVxp67_ASAP7_75t_L g171 ( .A(n_125), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_138), .Y(n_172) );
NOR2xp67_ASAP7_75t_L g173 ( .A(n_146), .B(n_89), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_150), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_150), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_131), .B(n_102), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_130), .B(n_110), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_130), .B(n_110), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_134), .B(n_100), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_138), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_134), .B(n_100), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_150), .Y(n_182) );
INVx3_ASAP7_75t_L g183 ( .A(n_166), .Y(n_183) );
INVxp67_ASAP7_75t_L g184 ( .A(n_143), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_144), .B(n_94), .Y(n_185) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_156), .A2(n_123), .B(n_124), .C(n_111), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_150), .Y(n_187) );
OR2x2_ASAP7_75t_L g188 ( .A(n_168), .B(n_94), .Y(n_188) );
AND2x6_ASAP7_75t_SL g189 ( .A(n_166), .B(n_117), .Y(n_189) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_128), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_150), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_128), .B(n_84), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_144), .B(n_84), .Y(n_193) );
INVxp67_ASAP7_75t_SL g194 ( .A(n_136), .Y(n_194) );
BUFx3_ASAP7_75t_L g195 ( .A(n_151), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_138), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_145), .B(n_80), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_136), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_138), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_139), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_166), .A2(n_80), .B1(n_117), .B2(n_13), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_145), .B(n_54), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_147), .B(n_9), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_147), .B(n_56), .Y(n_204) );
BUFx6f_ASAP7_75t_SL g205 ( .A(n_166), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g206 ( .A1(n_157), .A2(n_11), .B1(n_14), .B2(n_21), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_158), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_151), .Y(n_208) );
INVx4_ASAP7_75t_L g209 ( .A(n_146), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_139), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_139), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_153), .B(n_26), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_153), .B(n_29), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_156), .A2(n_30), .B(n_32), .C(n_34), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_149), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_154), .B(n_37), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_154), .B(n_38), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_139), .Y(n_218) );
NOR3xp33_ASAP7_75t_L g219 ( .A(n_157), .B(n_40), .C(n_46), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_160), .A2(n_49), .B1(n_50), .B2(n_51), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_158), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_149), .B(n_60), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_149), .B(n_61), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_158), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_158), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_219), .A2(n_155), .B1(n_163), .B2(n_162), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_209), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_177), .B(n_163), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_209), .Y(n_229) );
BUFx2_ASAP7_75t_L g230 ( .A(n_184), .Y(n_230) );
INVx3_ASAP7_75t_L g231 ( .A(n_209), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_205), .A2(n_146), .B1(n_152), .B2(n_137), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_194), .A2(n_155), .B1(n_162), .B2(n_161), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_215), .B(n_146), .Y(n_234) );
BUFx2_ASAP7_75t_L g235 ( .A(n_188), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_178), .B(n_160), .Y(n_236) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_188), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_179), .B(n_161), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_171), .B(n_167), .Y(n_239) );
AND2x4_ASAP7_75t_L g240 ( .A(n_192), .B(n_159), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_185), .B(n_167), .Y(n_241) );
BUFx2_ASAP7_75t_L g242 ( .A(n_190), .Y(n_242) );
OAI22xp5_ASAP7_75t_SL g243 ( .A1(n_206), .A2(n_133), .B1(n_165), .B2(n_126), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_203), .Y(n_244) );
INVx5_ASAP7_75t_L g245 ( .A(n_207), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_193), .B(n_140), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_215), .Y(n_247) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_195), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_195), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_197), .B(n_140), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_183), .Y(n_251) );
BUFx12f_ASAP7_75t_L g252 ( .A(n_189), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_183), .B(n_152), .Y(n_253) );
INVx5_ASAP7_75t_L g254 ( .A(n_207), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g255 ( .A1(n_205), .A2(n_198), .B1(n_190), .B2(n_183), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_205), .A2(n_198), .B1(n_181), .B2(n_201), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_207), .Y(n_257) );
AND2x4_ASAP7_75t_L g258 ( .A(n_186), .B(n_165), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_169), .Y(n_259) );
BUFx10_ASAP7_75t_L g260 ( .A(n_202), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_173), .B(n_127), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_221), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_176), .B(n_135), .Y(n_263) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_221), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_173), .B(n_148), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_204), .A2(n_142), .B1(n_137), .B2(n_135), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_217), .B(n_148), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_224), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_224), .Y(n_269) );
OR2x6_ASAP7_75t_L g270 ( .A(n_206), .B(n_164), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_216), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_170), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_225), .Y(n_273) );
AOI22x1_ASAP7_75t_L g274 ( .A1(n_225), .A2(n_142), .B1(n_151), .B2(n_158), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_220), .B(n_151), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_212), .B(n_129), .Y(n_276) );
AOI22xp5_ASAP7_75t_L g277 ( .A1(n_213), .A2(n_151), .B1(n_126), .B2(n_158), .Y(n_277) );
BUFx6f_ASAP7_75t_L g278 ( .A(n_222), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g279 ( .A1(n_223), .A2(n_151), .B1(n_129), .B2(n_132), .Y(n_279) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_170), .Y(n_280) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_174), .Y(n_281) );
BUFx3_ASAP7_75t_L g282 ( .A(n_174), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_175), .Y(n_283) );
BUFx2_ASAP7_75t_L g284 ( .A(n_214), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_172), .B(n_129), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_172), .B(n_129), .Y(n_286) );
OR2x2_ASAP7_75t_L g287 ( .A(n_175), .B(n_141), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_182), .A2(n_141), .B1(n_132), .B2(n_64), .Y(n_288) );
BUFx2_ASAP7_75t_L g289 ( .A(n_180), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_251), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_228), .A2(n_182), .B(n_187), .Y(n_291) );
OAI22xp5_ASAP7_75t_L g292 ( .A1(n_256), .A2(n_187), .B1(n_191), .B2(n_208), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_236), .A2(n_191), .B(n_208), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_238), .A2(n_218), .B(n_211), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_230), .B(n_218), .Y(n_295) );
BUFx12f_ASAP7_75t_L g296 ( .A(n_252), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_235), .B(n_211), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_253), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_237), .B(n_210), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_234), .A2(n_210), .B(n_200), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_287), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_253), .Y(n_302) );
INVx3_ASAP7_75t_L g303 ( .A(n_231), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_231), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_234), .A2(n_200), .B(n_199), .Y(n_305) );
BUFx2_ASAP7_75t_L g306 ( .A(n_242), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_286), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_259), .B(n_199), .Y(n_308) );
UNKNOWN g309 ( );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_239), .B(n_196), .Y(n_310) );
NAND2x1p5_ASAP7_75t_L g311 ( .A(n_227), .B(n_196), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_240), .B(n_180), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_248), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_263), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_229), .Y(n_315) );
INVxp67_ASAP7_75t_SL g316 ( .A(n_247), .Y(n_316) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_247), .Y(n_317) );
CKINVDCx11_ASAP7_75t_R g318 ( .A(n_270), .Y(n_318) );
INVx3_ASAP7_75t_L g319 ( .A(n_248), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_244), .B(n_141), .Y(n_320) );
AOI21x1_ASAP7_75t_SL g321 ( .A1(n_246), .A2(n_62), .B(n_63), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_250), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_285), .Y(n_323) );
A2O1A1Ixp33_ASAP7_75t_SL g324 ( .A1(n_241), .A2(n_267), .B(n_271), .C(n_232), .Y(n_324) );
NAND2xp5_ASAP7_75t_SL g325 ( .A(n_247), .B(n_141), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_258), .B(n_132), .Y(n_326) );
AND2x4_ASAP7_75t_L g327 ( .A(n_240), .B(n_65), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_270), .B(n_141), .Y(n_328) );
INVxp67_ASAP7_75t_SL g329 ( .A(n_255), .Y(n_329) );
INVx3_ASAP7_75t_L g330 ( .A(n_248), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_275), .A2(n_141), .B(n_132), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_289), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_278), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_270), .B(n_132), .Y(n_334) );
AOI21xp5_ASAP7_75t_SL g335 ( .A1(n_255), .A2(n_132), .B(n_69), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_272), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_284), .A2(n_67), .B(n_70), .Y(n_337) );
NAND2x1p5_ASAP7_75t_L g338 ( .A(n_265), .B(n_71), .Y(n_338) );
OAI22xp5_ASAP7_75t_SL g339 ( .A1(n_243), .A2(n_233), .B1(n_226), .B2(n_258), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_261), .B(n_74), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_283), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_336), .Y(n_342) );
AOI22xp5_ASAP7_75t_L g343 ( .A1(n_339), .A2(n_243), .B1(n_226), .B2(n_266), .Y(n_343) );
OAI21x1_ASAP7_75t_L g344 ( .A1(n_321), .A2(n_288), .B(n_279), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_318), .B(n_260), .Y(n_345) );
OAI21xp5_ASAP7_75t_L g346 ( .A1(n_298), .A2(n_277), .B(n_279), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_336), .Y(n_347) );
AND2x4_ASAP7_75t_L g348 ( .A(n_322), .B(n_276), .Y(n_348) );
OAI22xp33_ASAP7_75t_L g349 ( .A1(n_306), .A2(n_278), .B1(n_277), .B2(n_288), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_302), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_314), .Y(n_351) );
OAI21x1_ASAP7_75t_L g352 ( .A1(n_331), .A2(n_274), .B(n_249), .Y(n_352) );
BUFx12f_ASAP7_75t_L g353 ( .A(n_296), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_290), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_306), .Y(n_355) );
AND2x4_ASAP7_75t_L g356 ( .A(n_327), .B(n_278), .Y(n_356) );
OA21x2_ASAP7_75t_L g357 ( .A1(n_326), .A2(n_262), .B(n_268), .Y(n_357) );
INVx2_ASAP7_75t_SL g358 ( .A(n_313), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_341), .Y(n_359) );
INVx3_ASAP7_75t_L g360 ( .A(n_313), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_341), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_309), .B(n_260), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_290), .Y(n_363) );
BUFx2_ASAP7_75t_L g364 ( .A(n_295), .Y(n_364) );
AND2x4_ASAP7_75t_L g365 ( .A(n_327), .B(n_254), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_320), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_329), .B(n_308), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_315), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_320), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_315), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_308), .B(n_254), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_328), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_328), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_313), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_367), .B(n_299), .Y(n_375) );
INVx2_ASAP7_75t_SL g376 ( .A(n_355), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_342), .Y(n_377) );
AND2x4_ASAP7_75t_L g378 ( .A(n_350), .B(n_327), .Y(n_378) );
AND2x4_ASAP7_75t_L g379 ( .A(n_350), .B(n_334), .Y(n_379) );
NOR3xp33_ASAP7_75t_L g380 ( .A(n_362), .B(n_318), .C(n_334), .Y(n_380) );
NAND2x1p5_ASAP7_75t_SL g381 ( .A(n_367), .B(n_325), .Y(n_381) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_358), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_364), .B(n_297), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_351), .B(n_299), .Y(n_384) );
INVx2_ASAP7_75t_SL g385 ( .A(n_342), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_342), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_351), .B(n_295), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_347), .B(n_301), .Y(n_388) );
BUFx2_ASAP7_75t_L g389 ( .A(n_364), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_347), .B(n_301), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_347), .Y(n_391) );
NOR2x1_ASAP7_75t_SL g392 ( .A(n_359), .B(n_313), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_359), .B(n_307), .Y(n_393) );
NAND3xp33_ASAP7_75t_L g394 ( .A(n_343), .B(n_335), .C(n_337), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_343), .B(n_332), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_359), .B(n_297), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_361), .B(n_317), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_361), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_361), .B(n_323), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_354), .B(n_312), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_362), .B(n_324), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_370), .Y(n_402) );
AOI221xp5_ASAP7_75t_L g403 ( .A1(n_395), .A2(n_373), .B1(n_372), .B2(n_345), .C(n_348), .Y(n_403) );
OA21x2_ASAP7_75t_L g404 ( .A1(n_401), .A2(n_344), .B(n_346), .Y(n_404) );
INVxp67_ASAP7_75t_SL g405 ( .A(n_385), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_399), .B(n_373), .Y(n_406) );
AO21x2_ASAP7_75t_L g407 ( .A1(n_394), .A2(n_349), .B(n_344), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_377), .Y(n_408) );
BUFx2_ASAP7_75t_L g409 ( .A(n_385), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_386), .Y(n_410) );
OAI33xp33_ASAP7_75t_L g411 ( .A1(n_397), .A2(n_372), .A3(n_383), .B1(n_396), .B2(n_354), .B3(n_363), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_386), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_377), .B(n_370), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_391), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_386), .Y(n_415) );
AOI31xp33_ASAP7_75t_SL g416 ( .A1(n_380), .A2(n_370), .A3(n_353), .B(n_369), .Y(n_416) );
INVx2_ASAP7_75t_SL g417 ( .A(n_402), .Y(n_417) );
INVx3_ASAP7_75t_L g418 ( .A(n_382), .Y(n_418) );
INVx3_ASAP7_75t_L g419 ( .A(n_382), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_402), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_402), .Y(n_421) );
OAI21xp33_ASAP7_75t_L g422 ( .A1(n_394), .A2(n_335), .B(n_363), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_391), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_398), .B(n_368), .Y(n_424) );
AO21x2_ASAP7_75t_L g425 ( .A1(n_392), .A2(n_344), .B(n_381), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g426 ( .A1(n_387), .A2(n_348), .B1(n_369), .B2(n_366), .C(n_368), .Y(n_426) );
OAI22xp33_ASAP7_75t_L g427 ( .A1(n_389), .A2(n_353), .B1(n_366), .B2(n_369), .Y(n_427) );
OAI21x1_ASAP7_75t_L g428 ( .A1(n_398), .A2(n_374), .B(n_360), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_389), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_399), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_388), .Y(n_431) );
BUFx2_ASAP7_75t_L g432 ( .A(n_378), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_388), .Y(n_433) );
AO21x2_ASAP7_75t_L g434 ( .A1(n_392), .A2(n_346), .B(n_374), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_390), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_390), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_435), .B(n_375), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_424), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_430), .B(n_396), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_430), .B(n_375), .Y(n_440) );
INVxp67_ASAP7_75t_L g441 ( .A(n_411), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_403), .A2(n_378), .B1(n_379), .B2(n_384), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_424), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_424), .Y(n_444) );
INVxp67_ASAP7_75t_SL g445 ( .A(n_410), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_413), .B(n_376), .Y(n_446) );
NAND3xp33_ASAP7_75t_L g447 ( .A(n_403), .B(n_376), .C(n_340), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_408), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_435), .B(n_393), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_408), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_431), .B(n_383), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_435), .B(n_393), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_414), .Y(n_453) );
NOR2x1_ASAP7_75t_L g454 ( .A(n_416), .B(n_378), .Y(n_454) );
BUFx2_ASAP7_75t_L g455 ( .A(n_409), .Y(n_455) );
INVx1_ASAP7_75t_SL g456 ( .A(n_413), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_414), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_423), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_412), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_423), .Y(n_460) );
AND2x4_ASAP7_75t_L g461 ( .A(n_423), .B(n_379), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_413), .B(n_387), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_431), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_433), .B(n_384), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_433), .B(n_397), .Y(n_465) );
AND2x4_ASAP7_75t_L g466 ( .A(n_417), .B(n_379), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_412), .Y(n_467) );
OAI22xp33_ASAP7_75t_SL g468 ( .A1(n_429), .A2(n_378), .B1(n_379), .B2(n_338), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_436), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_436), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_406), .B(n_400), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_412), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_406), .B(n_400), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_410), .Y(n_474) );
INVxp67_ASAP7_75t_L g475 ( .A(n_411), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_429), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_426), .A2(n_356), .B1(n_348), .B2(n_365), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_415), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_426), .B(n_366), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_415), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_415), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_420), .B(n_381), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_420), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_420), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_448), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_442), .A2(n_432), .B1(n_427), .B2(n_422), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_450), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_462), .B(n_409), .Y(n_488) );
INVx1_ASAP7_75t_SL g489 ( .A(n_456), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_438), .B(n_417), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_453), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_457), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_446), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_443), .B(n_417), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_437), .B(n_405), .Y(n_495) );
BUFx3_ASAP7_75t_L g496 ( .A(n_455), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_463), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_469), .Y(n_498) );
OAI33xp33_ASAP7_75t_L g499 ( .A1(n_441), .A2(n_422), .A3(n_292), .B1(n_416), .B2(n_421), .B3(n_381), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_470), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_476), .Y(n_501) );
NOR2x1_ASAP7_75t_L g502 ( .A(n_454), .B(n_421), .Y(n_502) );
AND2x4_ASAP7_75t_SL g503 ( .A(n_437), .B(n_371), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_444), .B(n_421), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_449), .B(n_405), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_458), .Y(n_506) );
INVx1_ASAP7_75t_SL g507 ( .A(n_449), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_460), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_445), .B(n_432), .Y(n_509) );
NOR2xp67_ASAP7_75t_SL g510 ( .A(n_447), .B(n_353), .Y(n_510) );
INVxp67_ASAP7_75t_L g511 ( .A(n_445), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_452), .B(n_418), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_452), .B(n_418), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_474), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_471), .B(n_418), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_473), .B(n_418), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_468), .B(n_419), .Y(n_517) );
NAND3xp33_ASAP7_75t_L g518 ( .A(n_441), .B(n_404), .C(n_356), .Y(n_518) );
NAND2xp33_ASAP7_75t_L g519 ( .A(n_442), .B(n_382), .Y(n_519) );
OAI221xp5_ASAP7_75t_L g520 ( .A1(n_475), .A2(n_338), .B1(n_404), .B2(n_316), .C(n_371), .Y(n_520) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_459), .Y(n_521) );
INVx1_ASAP7_75t_SL g522 ( .A(n_439), .Y(n_522) );
INVxp67_ASAP7_75t_L g523 ( .A(n_478), .Y(n_523) );
INVxp67_ASAP7_75t_L g524 ( .A(n_480), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_451), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_477), .A2(n_356), .B1(n_365), .B2(n_419), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_461), .B(n_419), .Y(n_527) );
INVxp67_ASAP7_75t_L g528 ( .A(n_483), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_465), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_440), .B(n_419), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_475), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_459), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_467), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_461), .B(n_466), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_464), .Y(n_535) );
NAND2x1_ASAP7_75t_L g536 ( .A(n_466), .B(n_382), .Y(n_536) );
INVxp67_ASAP7_75t_L g537 ( .A(n_484), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_461), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_467), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_472), .Y(n_540) );
NOR3xp33_ASAP7_75t_L g541 ( .A(n_479), .B(n_356), .C(n_365), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_522), .B(n_482), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_501), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_507), .B(n_481), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_531), .B(n_466), .Y(n_545) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_521), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_535), .B(n_481), .Y(n_547) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_521), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_525), .B(n_472), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_489), .B(n_404), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_493), .B(n_404), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_529), .B(n_404), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_514), .B(n_434), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_485), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_534), .B(n_425), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_488), .B(n_434), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_512), .B(n_513), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_502), .B(n_428), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_497), .B(n_498), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_500), .B(n_434), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_487), .Y(n_561) );
A2O1A1Ixp33_ASAP7_75t_R g562 ( .A1(n_517), .A2(n_296), .B(n_365), .C(n_338), .Y(n_562) );
OAI21xp5_ASAP7_75t_L g563 ( .A1(n_510), .A2(n_428), .B(n_348), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_491), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_492), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_506), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_508), .Y(n_567) );
INVxp67_ASAP7_75t_L g568 ( .A(n_496), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_495), .B(n_434), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_505), .B(n_428), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_523), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_523), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_499), .B(n_425), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_524), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_524), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_532), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_533), .Y(n_577) );
NAND4xp25_ASAP7_75t_L g578 ( .A(n_486), .B(n_310), .C(n_294), .D(n_291), .Y(n_578) );
NAND2xp33_ASAP7_75t_L g579 ( .A(n_541), .B(n_382), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_527), .B(n_538), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_511), .B(n_382), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_503), .B(n_425), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_515), .B(n_425), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_528), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_516), .B(n_407), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_539), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_509), .B(n_407), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_528), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_537), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_537), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_511), .Y(n_591) );
OAI21xp5_ASAP7_75t_SL g592 ( .A1(n_541), .A2(n_360), .B(n_358), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_490), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_571), .B(n_494), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_559), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_572), .B(n_530), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_579), .A2(n_499), .B1(n_519), .B2(n_486), .Y(n_597) );
NOR4xp25_ASAP7_75t_L g598 ( .A(n_568), .B(n_520), .C(n_517), .D(n_518), .Y(n_598) );
NOR3x1_ASAP7_75t_L g599 ( .A(n_592), .B(n_520), .C(n_526), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_557), .B(n_509), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_580), .B(n_540), .Y(n_601) );
NAND4xp75_ASAP7_75t_L g602 ( .A(n_562), .B(n_504), .C(n_519), .D(n_357), .Y(n_602) );
OAI211xp5_ASAP7_75t_L g603 ( .A1(n_568), .A2(n_536), .B(n_357), .C(n_360), .Y(n_603) );
A2O1A1Ixp33_ASAP7_75t_SL g604 ( .A1(n_573), .A2(n_360), .B(n_330), .C(n_319), .Y(n_604) );
AOI211xp5_ASAP7_75t_SL g605 ( .A1(n_579), .A2(n_374), .B(n_330), .C(n_319), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_543), .B(n_407), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_580), .B(n_407), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_546), .B(n_358), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_574), .B(n_357), .Y(n_609) );
NOR3xp33_ASAP7_75t_L g610 ( .A(n_578), .B(n_330), .C(n_319), .Y(n_610) );
NOR2xp67_ASAP7_75t_L g611 ( .A(n_546), .B(n_75), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_545), .A2(n_593), .B1(n_582), .B2(n_556), .Y(n_612) );
OR2x2_ASAP7_75t_L g613 ( .A(n_542), .B(n_357), .Y(n_613) );
OAI211xp5_ASAP7_75t_L g614 ( .A1(n_563), .A2(n_293), .B(n_333), .C(n_300), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_555), .B(n_76), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_554), .B(n_561), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_564), .B(n_77), .Y(n_617) );
OAI211xp5_ASAP7_75t_L g618 ( .A1(n_585), .A2(n_333), .B(n_305), .C(n_304), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_565), .Y(n_619) );
AOI21xp33_ASAP7_75t_L g620 ( .A1(n_573), .A2(n_333), .B(n_313), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_566), .B(n_333), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_575), .B(n_333), .Y(n_622) );
AOI211xp5_ASAP7_75t_L g623 ( .A1(n_587), .A2(n_352), .B(n_304), .C(n_303), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_567), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_584), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_588), .Y(n_626) );
NOR3xp33_ASAP7_75t_L g627 ( .A(n_589), .B(n_303), .C(n_352), .Y(n_627) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_590), .A2(n_303), .B1(n_311), .B2(n_269), .C(n_273), .Y(n_628) );
OAI221xp5_ASAP7_75t_L g629 ( .A1(n_552), .A2(n_311), .B1(n_254), .B2(n_245), .C(n_257), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_591), .Y(n_630) );
NAND4xp25_ASAP7_75t_SL g631 ( .A(n_597), .B(n_570), .C(n_544), .D(n_550), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_619), .Y(n_632) );
O2A1O1Ixp33_ASAP7_75t_L g633 ( .A1(n_598), .A2(n_581), .B(n_548), .C(n_558), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_595), .B(n_549), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_624), .Y(n_635) );
AND2x4_ASAP7_75t_L g636 ( .A(n_600), .B(n_548), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_616), .A2(n_583), .B1(n_547), .B2(n_569), .C(n_553), .Y(n_637) );
NOR2xp67_ASAP7_75t_L g638 ( .A(n_603), .B(n_581), .Y(n_638) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_611), .B(n_558), .Y(n_639) );
AOI21xp5_ASAP7_75t_L g640 ( .A1(n_604), .A2(n_560), .B(n_551), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_596), .B(n_586), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_612), .B(n_586), .Y(n_642) );
AND2x4_ASAP7_75t_L g643 ( .A(n_625), .B(n_577), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_597), .B(n_576), .Y(n_644) );
NOR2x1p5_ASAP7_75t_L g645 ( .A(n_602), .B(n_576), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_626), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_616), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_630), .B(n_577), .Y(n_648) );
NOR3xp33_ASAP7_75t_L g649 ( .A(n_610), .B(n_352), .C(n_311), .Y(n_649) );
NOR2x1_ASAP7_75t_L g650 ( .A(n_608), .B(n_282), .Y(n_650) );
INVx1_ASAP7_75t_SL g651 ( .A(n_601), .Y(n_651) );
INVxp33_ASAP7_75t_SL g652 ( .A(n_599), .Y(n_652) );
NOR3xp33_ASAP7_75t_L g653 ( .A(n_610), .B(n_245), .C(n_264), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_641), .Y(n_654) );
BUFx2_ASAP7_75t_L g655 ( .A(n_636), .Y(n_655) );
NOR3x1_ASAP7_75t_L g656 ( .A(n_652), .B(n_594), .C(n_614), .Y(n_656) );
AOI32xp33_ASAP7_75t_L g657 ( .A1(n_651), .A2(n_605), .A3(n_607), .B1(n_615), .B2(n_617), .Y(n_657) );
OAI211xp5_ASAP7_75t_L g658 ( .A1(n_633), .A2(n_606), .B(n_623), .C(n_618), .Y(n_658) );
INVxp33_ASAP7_75t_L g659 ( .A(n_650), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_637), .B(n_606), .Y(n_660) );
OAI211xp5_ASAP7_75t_SL g661 ( .A1(n_644), .A2(n_620), .B(n_629), .C(n_613), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_631), .A2(n_627), .B1(n_621), .B2(n_609), .Y(n_662) );
NAND3xp33_ASAP7_75t_L g663 ( .A(n_640), .B(n_627), .C(n_622), .Y(n_663) );
OR2x2_ASAP7_75t_L g664 ( .A(n_642), .B(n_628), .Y(n_664) );
NOR3xp33_ASAP7_75t_L g665 ( .A(n_639), .B(n_245), .C(n_264), .Y(n_665) );
NAND4xp75_ASAP7_75t_L g666 ( .A(n_638), .B(n_264), .C(n_280), .D(n_281), .Y(n_666) );
AND2x4_ASAP7_75t_L g667 ( .A(n_645), .B(n_280), .Y(n_667) );
XNOR2x1_ASAP7_75t_L g668 ( .A(n_664), .B(n_636), .Y(n_668) );
XOR2xp5_ASAP7_75t_L g669 ( .A(n_659), .B(n_647), .Y(n_669) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_654), .Y(n_670) );
BUFx2_ASAP7_75t_L g671 ( .A(n_655), .Y(n_671) );
INVx4_ASAP7_75t_L g672 ( .A(n_667), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_660), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_656), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_667), .Y(n_675) );
NAND3xp33_ASAP7_75t_SL g676 ( .A(n_674), .B(n_657), .C(n_662), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_670), .Y(n_677) );
OAI221xp5_ASAP7_75t_L g678 ( .A1(n_671), .A2(n_658), .B1(n_663), .B2(n_665), .C(n_661), .Y(n_678) );
NAND3xp33_ASAP7_75t_SL g679 ( .A(n_673), .B(n_653), .C(n_649), .Y(n_679) );
OAI322xp33_ASAP7_75t_L g680 ( .A1(n_678), .A2(n_669), .A3(n_668), .B1(n_670), .B2(n_672), .C1(n_675), .C2(n_634), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g681 ( .A1(n_676), .A2(n_675), .B(n_672), .Y(n_681) );
OAI211xp5_ASAP7_75t_SL g682 ( .A1(n_677), .A2(n_632), .B(n_635), .C(n_646), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_681), .B(n_679), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_680), .A2(n_648), .B(n_643), .Y(n_684) );
OAI222xp33_ASAP7_75t_L g685 ( .A1(n_683), .A2(n_682), .B1(n_643), .B2(n_666), .C1(n_281), .C2(n_280), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_685), .A2(n_684), .B(n_281), .Y(n_686) );
endmodule