module real_jpeg_5872_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_0),
.A2(n_90),
.B1(n_92),
.B2(n_94),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_0),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_0),
.A2(n_94),
.B1(n_127),
.B2(n_131),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_0),
.A2(n_94),
.B1(n_145),
.B2(n_147),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_0),
.A2(n_94),
.B1(n_399),
.B2(n_400),
.Y(n_398)
);

BUFx5_ASAP7_75t_L g197 ( 
.A(n_1),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_1),
.Y(n_204)
);

INVx8_ASAP7_75t_L g233 ( 
.A(n_1),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_1),
.Y(n_243)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_1),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_1),
.Y(n_432)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_2),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_2),
.Y(n_146)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_2),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_2),
.Y(n_438)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_3),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_3),
.A2(n_54),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

OAI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_3),
.A2(n_54),
.B1(n_403),
.B2(n_404),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_SL g412 ( 
.A1(n_3),
.A2(n_54),
.B1(n_92),
.B2(n_413),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_4),
.A2(n_207),
.B1(n_285),
.B2(n_287),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_4),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_4),
.A2(n_287),
.B1(n_382),
.B2(n_384),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_4),
.A2(n_274),
.B1(n_287),
.B2(n_411),
.Y(n_410)
);

OAI22xp33_ASAP7_75t_L g465 ( 
.A1(n_4),
.A2(n_287),
.B1(n_345),
.B2(n_466),
.Y(n_465)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_6),
.A2(n_161),
.B1(n_164),
.B2(n_168),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_6),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_6),
.B(n_178),
.C(n_180),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_6),
.B(n_74),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_6),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_6),
.B(n_125),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_6),
.B(n_274),
.Y(n_273)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_7),
.Y(n_542)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_8),
.Y(n_105)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_8),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_8),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_9),
.A2(n_83),
.B1(n_84),
.B2(n_87),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_9),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_9),
.A2(n_87),
.B1(n_134),
.B2(n_139),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_9),
.A2(n_87),
.B1(n_395),
.B2(n_396),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_9),
.A2(n_87),
.B1(n_403),
.B2(n_420),
.Y(n_419)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_11),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_11),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_11),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_12),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_12),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_12),
.A2(n_191),
.B1(n_216),
.B2(n_238),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_12),
.A2(n_216),
.B1(n_315),
.B2(n_317),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_12),
.A2(n_51),
.B1(n_216),
.B2(n_436),
.Y(n_435)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_13),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_14),
.Y(n_546)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_16),
.A2(n_185),
.B1(n_189),
.B2(n_190),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_16),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_16),
.A2(n_176),
.B1(n_189),
.B2(n_264),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g379 ( 
.A1(n_16),
.A2(n_91),
.B1(n_189),
.B2(n_279),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_16),
.A2(n_51),
.B1(n_53),
.B2(n_189),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_17),
.A2(n_58),
.B1(n_60),
.B2(n_62),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_17),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g363 ( 
.A1(n_17),
.A2(n_62),
.B1(n_187),
.B2(n_326),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_17),
.A2(n_62),
.B1(n_131),
.B2(n_407),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_17),
.A2(n_62),
.B1(n_450),
.B2(n_452),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_18),
.A2(n_110),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_18),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_18),
.A2(n_171),
.B1(n_206),
.B2(n_208),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_18),
.A2(n_85),
.B1(n_171),
.B2(n_278),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_18),
.A2(n_171),
.B1(n_371),
.B2(n_376),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_540),
.B(n_543),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_150),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_148),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_143),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_23),
.B(n_143),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_132),
.C(n_140),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_24),
.A2(n_25),
.B1(n_536),
.B2(n_537),
.Y(n_535)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_63),
.C(n_95),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g527 ( 
.A(n_26),
.B(n_528),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_50),
.B1(n_55),
.B2(n_57),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_27),
.A2(n_55),
.B1(n_57),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_27),
.A2(n_55),
.B1(n_133),
.B2(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_27),
.A2(n_374),
.B(n_415),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_27),
.A2(n_55),
.B1(n_415),
.B2(n_435),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_27),
.A2(n_50),
.B1(n_55),
.B2(n_513),
.Y(n_512)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_28),
.A2(n_370),
.B(n_373),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_28),
.B(n_375),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_36),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_SL g347 ( 
.A(n_32),
.Y(n_347)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_40),
.B1(n_44),
.B2(n_48),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_39),
.Y(n_349)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx5_ASAP7_75t_L g453 ( 
.A(n_42),
.Y(n_453)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_43),
.Y(n_271)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_43),
.Y(n_280)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_43),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_43),
.Y(n_451)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_47),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_47),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_53),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_55),
.B(n_168),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_55),
.A2(n_435),
.B(n_467),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_56),
.B(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_56),
.B(n_465),
.Y(n_464)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_59),
.Y(n_356)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_59),
.Y(n_466)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_63),
.A2(n_95),
.B1(n_96),
.B2(n_529),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_63),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_82),
.B1(n_88),
.B2(n_89),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_64),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_64),
.A2(n_88),
.B1(n_314),
.B2(n_379),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_64),
.A2(n_88),
.B1(n_410),
.B2(n_412),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_64),
.A2(n_82),
.B1(n_88),
.B2(n_517),
.Y(n_516)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_74),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_70),
.Y(n_296)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_70),
.Y(n_303)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_74),
.A2(n_141),
.B(n_142),
.Y(n_140)
);

AOI22x1_ASAP7_75t_L g439 ( 
.A1(n_74),
.A2(n_141),
.B1(n_321),
.B2(n_440),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_74),
.A2(n_141),
.B1(n_448),
.B2(n_449),
.Y(n_447)
);

AO22x2_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_78),
.B2(n_80),
.Y(n_74)
);

INVx5_ASAP7_75t_L g383 ( 
.A(n_76),
.Y(n_383)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_77),
.Y(n_215)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_77),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_77),
.Y(n_264)
);

INVx11_ASAP7_75t_L g172 ( 
.A(n_78),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_79),
.Y(n_163)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_79),
.Y(n_167)
);

INVx6_ASAP7_75t_L g422 ( 
.A(n_79),
.Y(n_422)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_88),
.B(n_277),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_88),
.A2(n_314),
.B(n_320),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI32xp33_ASAP7_75t_L g290 ( 
.A1(n_91),
.A2(n_273),
.A3(n_291),
.B1(n_293),
.B2(n_297),
.Y(n_290)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_93),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_95),
.A2(n_96),
.B1(n_515),
.B2(n_516),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_95),
.B(n_512),
.C(n_515),
.Y(n_523)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_124),
.B(n_126),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_97),
.A2(n_160),
.B(n_169),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_97),
.A2(n_124),
.B1(n_214),
.B2(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_97),
.A2(n_169),
.B(n_263),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_97),
.A2(n_124),
.B1(n_381),
.B2(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_98),
.B(n_170),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_98),
.A2(n_125),
.B1(n_402),
.B2(n_406),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_98),
.A2(n_125),
.B1(n_406),
.B2(n_419),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_98),
.A2(n_125),
.B1(n_419),
.B2(n_456),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_113),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_103),
.B1(n_106),
.B2(n_110),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_107),
.A2(n_114),
.B1(n_118),
.B2(n_121),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_SL g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_112),
.Y(n_385)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_113),
.A2(n_214),
.B(n_220),
.Y(n_213)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_116),
.Y(n_181)
);

INVx8_ASAP7_75t_L g327 ( 
.A(n_116),
.Y(n_327)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_116),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_117),
.Y(n_194)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_120),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_120),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_120),
.Y(n_286)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_123),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_124),
.A2(n_220),
.B(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_125),
.B(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_126),
.Y(n_456)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_132),
.B(n_140),
.Y(n_537)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_138),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_141),
.A2(n_267),
.B(n_276),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_141),
.B(n_321),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_141),
.A2(n_276),
.B(n_480),
.Y(n_479)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_534),
.B(n_539),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_506),
.B(n_531),
.Y(n_151)
);

OAI311xp33_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_388),
.A3(n_482),
.B1(n_500),
.C1(n_505),
.Y(n_152)
);

AOI21x1_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_333),
.B(n_387),
.Y(n_153)
);

AO21x1_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_305),
.B(n_332),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_257),
.B(n_304),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_223),
.B(n_256),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_182),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_158),
.B(n_182),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_173),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_159),
.A2(n_173),
.B1(n_174),
.B2(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_159),
.Y(n_254)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_163),
.Y(n_407)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_167),
.Y(n_292)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_167),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_168),
.A2(n_195),
.B(n_202),
.Y(n_234)
);

OAI21xp33_ASAP7_75t_SL g267 ( 
.A1(n_168),
.A2(n_268),
.B(n_272),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_168),
.B(n_354),
.Y(n_353)
);

OAI21xp33_ASAP7_75t_SL g370 ( 
.A1(n_168),
.A2(n_353),
.B(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_172),
.Y(n_403)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_211),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_183),
.B(n_212),
.C(n_222),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_195),
.B(n_202),
.Y(n_183)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_184),
.Y(n_250)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_187),
.Y(n_396)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx4_ASAP7_75t_SL g191 ( 
.A(n_192),
.Y(n_191)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_194),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_194),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_195),
.A2(n_359),
.B1(n_360),
.B2(n_362),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_195),
.A2(n_394),
.B1(n_397),
.B2(n_398),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_195),
.A2(n_329),
.B(n_398),
.Y(n_423)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_196),
.B(n_205),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_196),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_196),
.A2(n_284),
.B1(n_325),
.B2(n_328),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_196),
.A2(n_363),
.B1(n_430),
.B2(n_431),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_201),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx3_ASAP7_75t_SL g209 ( 
.A(n_210),
.Y(n_209)
);

INVx5_ASAP7_75t_L g326 ( 
.A(n_210),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_221),
.B2(n_222),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_215),
.Y(n_405)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_247),
.B(n_255),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_235),
.B(n_246),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_234),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_231),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_228),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_233),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_245),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_245),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_241),
.B(n_244),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_237),
.Y(n_249)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx3_ASAP7_75t_SL g241 ( 
.A(n_242),
.Y(n_241)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_243),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_244),
.A2(n_283),
.B(n_288),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_253),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_253),
.Y(n_255)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_258),
.B(n_259),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_281),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_265),
.B2(n_266),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_262),
.B(n_265),
.C(n_281),
.Y(n_306)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_271),
.Y(n_316)
);

INVxp33_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_277),
.Y(n_321)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_280),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_290),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_282),
.B(n_290),
.Y(n_311)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp33_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_301),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_306),
.B(n_307),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_312),
.B2(n_331),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_310),
.B(n_311),
.C(n_331),
.Y(n_334)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_312),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_322),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_313),
.B(n_323),
.C(n_324),
.Y(n_364)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_325),
.Y(n_359)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_326),
.Y(n_399)
);

INVx4_ASAP7_75t_L g400 ( 
.A(n_327),
.Y(n_400)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_328),
.Y(n_397)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx8_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_334),
.B(n_335),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_367),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_364),
.B1(n_365),
.B2(n_366),
.Y(n_336)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_337),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_339),
.B1(n_357),
.B2(n_358),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_339),
.B(n_357),
.Y(n_478)
);

OAI32xp33_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_343),
.A3(n_346),
.B1(n_348),
.B2(n_353),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_342),
.Y(n_411)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx8_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_364),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_364),
.B(n_365),
.C(n_367),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_369),
.B1(n_377),
.B2(n_386),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_368),
.B(n_378),
.C(n_380),
.Y(n_491)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx6_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_377),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_378),
.B(n_380),
.Y(n_377)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_379),
.Y(n_480)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx5_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

NAND2xp33_ASAP7_75t_SL g388 ( 
.A(n_389),
.B(n_468),
.Y(n_388)
);

A2O1A1Ixp33_ASAP7_75t_SL g500 ( 
.A1(n_389),
.A2(n_468),
.B(n_501),
.C(n_504),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_441),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_390),
.B(n_441),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_416),
.C(n_425),
.Y(n_390)
);

FAx1_ASAP7_75t_SL g481 ( 
.A(n_391),
.B(n_416),
.CI(n_425),
.CON(n_481),
.SN(n_481)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_408),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_392),
.B(n_409),
.C(n_414),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_401),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_393),
.B(n_401),
.Y(n_474)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_394),
.Y(n_430)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_402),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g404 ( 
.A(n_405),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_414),
.Y(n_408)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_410),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_412),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_417),
.A2(n_418),
.B1(n_423),
.B2(n_424),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_418),
.B(n_423),
.Y(n_460)
);

INVx3_ASAP7_75t_SL g420 ( 
.A(n_421),
.Y(n_420)
);

INVx8_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_423),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_423),
.A2(n_424),
.B1(n_462),
.B2(n_463),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_423),
.A2(n_460),
.B(n_463),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_433),
.C(n_439),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_426),
.B(n_472),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_427),
.B(n_429),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_427),
.B(n_429),
.Y(n_490)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_433),
.A2(n_434),
.B1(n_439),
.B2(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx8_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g473 ( 
.A(n_439),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_443),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_442),
.B(n_445),
.C(n_458),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_444),
.A2(n_445),
.B1(n_458),
.B2(n_459),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_446),
.A2(n_454),
.B(n_457),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_447),
.B(n_455),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_449),
.Y(n_517)
);

INVx6_ASAP7_75t_SL g450 ( 
.A(n_451),
.Y(n_450)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

FAx1_ASAP7_75t_SL g508 ( 
.A(n_457),
.B(n_509),
.CI(n_510),
.CON(n_508),
.SN(n_508)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_457),
.B(n_509),
.C(n_510),
.Y(n_530)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_461),
.Y(n_459)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_467),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_465),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_481),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_469),
.B(n_481),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_474),
.C(n_475),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_470),
.A2(n_471),
.B1(n_474),
.B2(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_474),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_475),
.B(n_493),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_478),
.C(n_479),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_476),
.A2(n_477),
.B1(n_479),
.B2(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_478),
.B(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_479),
.Y(n_488)
);

BUFx24_ASAP7_75t_SL g549 ( 
.A(n_481),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_483),
.B(n_495),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_484),
.A2(n_502),
.B(n_503),
.Y(n_501)
);

NOR2x1_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_492),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_485),
.B(n_492),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_489),
.C(n_491),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_486),
.B(n_498),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_489),
.A2(n_490),
.B1(n_491),
.B2(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_491),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_497),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_496),
.B(n_497),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_520),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_508),
.B(n_519),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_508),
.B(n_519),
.Y(n_532)
);

BUFx24_ASAP7_75t_SL g548 ( 
.A(n_508),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_511),
.A2(n_512),
.B1(n_514),
.B2(n_518),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_511),
.A2(n_512),
.B1(n_526),
.B2(n_527),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_511),
.B(n_522),
.C(n_526),
.Y(n_538)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_514),
.Y(n_518)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_520),
.A2(n_532),
.B(n_533),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_521),
.B(n_530),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_521),
.B(n_530),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_522),
.A2(n_523),
.B1(n_524),
.B2(n_525),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_535),
.B(n_538),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_535),
.B(n_538),
.Y(n_539)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx5_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx13_ASAP7_75t_L g545 ( 
.A(n_542),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_544),
.B(n_546),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);


endmodule