module real_aes_9079_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g509 ( .A1(n_0), .A2(n_173), .B(n_510), .C(n_513), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_1), .B(n_505), .Y(n_514) );
INVx1_ASAP7_75t_L g114 ( .A(n_2), .Y(n_114) );
INVx1_ASAP7_75t_L g171 ( .A(n_3), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_4), .B(n_174), .Y(n_578) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_5), .A2(n_127), .B1(n_130), .B2(n_131), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_5), .Y(n_131) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_6), .A2(n_473), .B(n_549), .Y(n_548) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_7), .A2(n_181), .B(n_528), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_8), .A2(n_38), .B1(n_161), .B2(n_209), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_9), .B(n_181), .Y(n_189) );
AND2x6_ASAP7_75t_L g176 ( .A(n_10), .B(n_177), .Y(n_176) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_11), .A2(n_176), .B(n_478), .C(n_522), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g127 ( .A1(n_12), .A2(n_42), .B1(n_128), .B2(n_129), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_12), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_13), .B(n_39), .Y(n_115) );
INVx1_ASAP7_75t_L g155 ( .A(n_14), .Y(n_155) );
INVx1_ASAP7_75t_L g152 ( .A(n_15), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_16), .B(n_157), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_17), .B(n_174), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_18), .B(n_148), .Y(n_255) );
AO32x2_ASAP7_75t_L g225 ( .A1(n_19), .A2(n_147), .A3(n_181), .B1(n_200), .B2(n_226), .Y(n_225) );
AOI222xp33_ASAP7_75t_SL g125 ( .A1(n_20), .A2(n_126), .B1(n_132), .B2(n_751), .C1(n_752), .C2(n_754), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_21), .B(n_161), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_22), .B(n_148), .Y(n_178) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_23), .A2(n_57), .B1(n_161), .B2(n_209), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_24), .Y(n_124) );
AOI22xp33_ASAP7_75t_SL g211 ( .A1(n_25), .A2(n_84), .B1(n_157), .B2(n_161), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_26), .B(n_161), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_27), .A2(n_200), .B(n_478), .C(n_496), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_28), .A2(n_200), .B(n_478), .C(n_531), .Y(n_530) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_29), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_30), .B(n_202), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_31), .A2(n_473), .B(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_32), .B(n_202), .Y(n_243) );
INVx2_ASAP7_75t_L g159 ( .A(n_33), .Y(n_159) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_34), .A2(n_476), .B(n_480), .C(n_486), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_35), .B(n_161), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_36), .B(n_202), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_37), .B(n_220), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_40), .B(n_494), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_41), .Y(n_526) );
INVx1_ASAP7_75t_L g129 ( .A(n_42), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_43), .B(n_174), .Y(n_543) );
OAI22xp5_ASAP7_75t_SL g764 ( .A1(n_44), .A2(n_765), .B1(n_767), .B2(n_768), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_44), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_45), .B(n_473), .Y(n_529) );
OAI22xp5_ASAP7_75t_SL g134 ( .A1(n_46), .A2(n_135), .B1(n_136), .B2(n_457), .Y(n_134) );
INVx1_ASAP7_75t_L g457 ( .A(n_46), .Y(n_457) );
OAI22xp5_ASAP7_75t_SL g765 ( .A1(n_46), .A2(n_48), .B1(n_457), .B2(n_766), .Y(n_765) );
A2O1A1Ixp33_ASAP7_75t_L g540 ( .A1(n_47), .A2(n_476), .B(n_486), .C(n_541), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_48), .Y(n_766) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_49), .B(n_161), .Y(n_184) );
INVx1_ASAP7_75t_L g511 ( .A(n_50), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g208 ( .A1(n_51), .A2(n_93), .B1(n_209), .B2(n_210), .Y(n_208) );
INVx1_ASAP7_75t_L g542 ( .A(n_52), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_53), .B(n_161), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_54), .B(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_55), .B(n_473), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_56), .B(n_169), .Y(n_188) );
AOI22xp33_ASAP7_75t_SL g253 ( .A1(n_58), .A2(n_62), .B1(n_157), .B2(n_161), .Y(n_253) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_59), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_60), .B(n_161), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_61), .B(n_161), .Y(n_217) );
INVx1_ASAP7_75t_L g177 ( .A(n_63), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_64), .B(n_473), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_65), .B(n_505), .Y(n_554) );
A2O1A1Ixp33_ASAP7_75t_L g551 ( .A1(n_66), .A2(n_163), .B(n_169), .C(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_67), .B(n_161), .Y(n_172) );
INVx1_ASAP7_75t_L g151 ( .A(n_68), .Y(n_151) );
OAI22xp33_ASAP7_75t_SL g761 ( .A1(n_69), .A2(n_762), .B1(n_769), .B2(n_770), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_69), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_70), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_71), .B(n_174), .Y(n_484) );
AO32x2_ASAP7_75t_L g206 ( .A1(n_72), .A2(n_181), .A3(n_200), .B1(n_207), .B2(n_212), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_73), .B(n_175), .Y(n_523) );
INVx1_ASAP7_75t_L g196 ( .A(n_74), .Y(n_196) );
INVx1_ASAP7_75t_L g238 ( .A(n_75), .Y(n_238) );
CKINVDCx16_ASAP7_75t_R g508 ( .A(n_76), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_77), .A2(n_105), .B1(n_116), .B2(n_772), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_78), .B(n_483), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g575 ( .A1(n_79), .A2(n_478), .B(n_486), .C(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_80), .B(n_157), .Y(n_239) );
CKINVDCx16_ASAP7_75t_R g550 ( .A(n_81), .Y(n_550) );
INVx1_ASAP7_75t_L g109 ( .A(n_82), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_83), .B(n_482), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_85), .B(n_209), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_86), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_87), .B(n_157), .Y(n_242) );
INVx2_ASAP7_75t_L g149 ( .A(n_88), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g582 ( .A(n_89), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_90), .B(n_199), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_91), .B(n_157), .Y(n_185) );
OR2x2_ASAP7_75t_L g111 ( .A(n_92), .B(n_112), .Y(n_111) );
OR2x2_ASAP7_75t_L g460 ( .A(n_92), .B(n_113), .Y(n_460) );
INVx2_ASAP7_75t_L g464 ( .A(n_92), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_94), .A2(n_103), .B1(n_157), .B2(n_158), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_95), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g481 ( .A(n_96), .Y(n_481) );
INVxp67_ASAP7_75t_L g553 ( .A(n_97), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_98), .B(n_157), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_99), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g519 ( .A(n_100), .Y(n_519) );
INVx1_ASAP7_75t_L g577 ( .A(n_101), .Y(n_577) );
AND2x2_ASAP7_75t_L g544 ( .A(n_102), .B(n_202), .Y(n_544) );
CKINVDCx6p67_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g773 ( .A(n_106), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .Y(n_106) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_111), .Y(n_123) );
HB1xp67_ASAP7_75t_L g771 ( .A(n_111), .Y(n_771) );
NOR2x2_ASAP7_75t_L g756 ( .A(n_112), .B(n_464), .Y(n_756) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
OR2x2_ASAP7_75t_L g463 ( .A(n_113), .B(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
BUFx3_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI22xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_125), .B1(n_757), .B2(n_760), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g118 ( .A(n_119), .B(n_122), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g759 ( .A(n_121), .Y(n_759) );
AOI21xp5_ASAP7_75t_L g760 ( .A1(n_122), .A2(n_761), .B(n_771), .Y(n_760) );
NOR2xp33_ASAP7_75t_SL g122 ( .A(n_123), .B(n_124), .Y(n_122) );
INVx1_ASAP7_75t_L g751 ( .A(n_126), .Y(n_751) );
CKINVDCx14_ASAP7_75t_R g130 ( .A(n_127), .Y(n_130) );
OAI22x1_ASAP7_75t_SL g132 ( .A1(n_133), .A2(n_458), .B1(n_461), .B2(n_465), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OAI22xp5_ASAP7_75t_SL g752 ( .A1(n_134), .A2(n_458), .B1(n_463), .B2(n_753), .Y(n_752) );
OAI22xp5_ASAP7_75t_SL g762 ( .A1(n_135), .A2(n_136), .B1(n_763), .B2(n_764), .Y(n_762) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_SL g136 ( .A(n_137), .B(n_423), .Y(n_136) );
NOR3xp33_ASAP7_75t_L g137 ( .A(n_138), .B(n_327), .C(n_411), .Y(n_137) );
NAND4xp25_ASAP7_75t_L g138 ( .A(n_139), .B(n_270), .C(n_292), .D(n_308), .Y(n_138) );
AOI221xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_203), .B1(n_229), .B2(n_248), .C(n_256), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_179), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_142), .B(n_248), .Y(n_282) );
NAND4xp25_ASAP7_75t_L g322 ( .A(n_142), .B(n_310), .C(n_323), .D(n_325), .Y(n_322) );
INVxp67_ASAP7_75t_L g439 ( .A(n_142), .Y(n_439) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
OR2x2_ASAP7_75t_L g321 ( .A(n_143), .B(n_259), .Y(n_321) );
AND2x2_ASAP7_75t_L g345 ( .A(n_143), .B(n_179), .Y(n_345) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g312 ( .A(n_144), .B(n_247), .Y(n_312) );
AND2x2_ASAP7_75t_L g352 ( .A(n_144), .B(n_333), .Y(n_352) );
AND2x2_ASAP7_75t_L g369 ( .A(n_144), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_144), .B(n_180), .Y(n_393) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g246 ( .A(n_145), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g264 ( .A(n_145), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g276 ( .A(n_145), .B(n_180), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_145), .B(n_190), .Y(n_298) );
OA21x2_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_153), .B(n_178), .Y(n_145) );
OA21x2_ASAP7_75t_L g190 ( .A1(n_146), .A2(n_191), .B(n_201), .Y(n_190) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_147), .B(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_148), .Y(n_181) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
AND2x2_ASAP7_75t_SL g202 ( .A(n_149), .B(n_150), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
OAI21xp5_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_167), .B(n_176), .Y(n_153) );
O2A1O1Ixp33_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_160), .C(n_163), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_156), .A2(n_523), .B(n_524), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_156), .A2(n_532), .B(n_533), .Y(n_531) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g162 ( .A(n_159), .Y(n_162) );
INVx1_ASAP7_75t_L g170 ( .A(n_159), .Y(n_170) );
INVx3_ASAP7_75t_L g237 ( .A(n_161), .Y(n_237) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_161), .Y(n_579) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g209 ( .A(n_162), .Y(n_209) );
BUFx3_ASAP7_75t_L g210 ( .A(n_162), .Y(n_210) );
AND2x6_ASAP7_75t_L g478 ( .A(n_162), .B(n_479), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g576 ( .A1(n_163), .A2(n_577), .B(n_578), .C(n_579), .Y(n_576) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_164), .A2(n_241), .B(n_242), .Y(n_240) );
INVx4_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g483 ( .A(n_165), .Y(n_483) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx3_ASAP7_75t_L g175 ( .A(n_166), .Y(n_175) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_166), .Y(n_199) );
INVx1_ASAP7_75t_L g220 ( .A(n_166), .Y(n_220) );
AND2x2_ASAP7_75t_L g474 ( .A(n_166), .B(n_170), .Y(n_474) );
INVx1_ASAP7_75t_L g479 ( .A(n_166), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_171), .B(n_172), .C(n_173), .Y(n_167) );
O2A1O1Ixp5_ASAP7_75t_L g195 ( .A1(n_168), .A2(n_196), .B(n_197), .C(n_198), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_168), .A2(n_497), .B(n_498), .Y(n_496) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_173), .A2(n_187), .B(n_188), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_173), .A2(n_199), .B1(n_227), .B2(n_228), .Y(n_226) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_173), .A2(n_199), .B1(n_252), .B2(n_253), .Y(n_251) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_174), .A2(n_184), .B(n_185), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_174), .A2(n_193), .B(n_194), .Y(n_192) );
O2A1O1Ixp5_ASAP7_75t_SL g236 ( .A1(n_174), .A2(n_237), .B(n_238), .C(n_239), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_174), .B(n_553), .Y(n_552) );
INVx5_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
OAI22xp5_ASAP7_75t_SL g207 ( .A1(n_175), .A2(n_199), .B1(n_208), .B2(n_211), .Y(n_207) );
OAI21xp5_ASAP7_75t_L g182 ( .A1(n_176), .A2(n_183), .B(n_186), .Y(n_182) );
BUFx3_ASAP7_75t_L g200 ( .A(n_176), .Y(n_200) );
OAI21xp5_ASAP7_75t_L g215 ( .A1(n_176), .A2(n_216), .B(n_221), .Y(n_215) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_176), .A2(n_236), .B(n_240), .Y(n_235) );
AND2x4_ASAP7_75t_L g473 ( .A(n_176), .B(n_474), .Y(n_473) );
INVx4_ASAP7_75t_SL g487 ( .A(n_176), .Y(n_487) );
NAND2x1p5_ASAP7_75t_L g520 ( .A(n_176), .B(n_474), .Y(n_520) );
AND2x2_ASAP7_75t_L g279 ( .A(n_179), .B(n_280), .Y(n_279) );
AOI221xp5_ASAP7_75t_L g328 ( .A1(n_179), .A2(n_329), .B1(n_332), .B2(n_334), .C(n_338), .Y(n_328) );
AND2x2_ASAP7_75t_L g387 ( .A(n_179), .B(n_352), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_179), .B(n_369), .Y(n_421) );
AND2x2_ASAP7_75t_L g179 ( .A(n_180), .B(n_190), .Y(n_179) );
INVx3_ASAP7_75t_L g247 ( .A(n_180), .Y(n_247) );
AND2x2_ASAP7_75t_L g296 ( .A(n_180), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g350 ( .A(n_180), .B(n_265), .Y(n_350) );
AND2x2_ASAP7_75t_L g408 ( .A(n_180), .B(n_409), .Y(n_408) );
OA21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_189), .Y(n_180) );
INVx4_ASAP7_75t_L g250 ( .A(n_181), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_181), .A2(n_529), .B(n_530), .Y(n_528) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_181), .Y(n_547) );
AND2x2_ASAP7_75t_L g248 ( .A(n_190), .B(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g265 ( .A(n_190), .Y(n_265) );
INVx1_ASAP7_75t_L g320 ( .A(n_190), .Y(n_320) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_190), .Y(n_326) );
AND2x2_ASAP7_75t_L g371 ( .A(n_190), .B(n_247), .Y(n_371) );
OR2x2_ASAP7_75t_L g410 ( .A(n_190), .B(n_249), .Y(n_410) );
OAI21xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_195), .B(n_200), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_198), .A2(n_222), .B(n_223), .Y(n_221) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx4_ASAP7_75t_L g512 ( .A(n_199), .Y(n_512) );
NAND3xp33_ASAP7_75t_L g269 ( .A(n_200), .B(n_250), .C(n_251), .Y(n_269) );
INVx2_ASAP7_75t_L g212 ( .A(n_202), .Y(n_212) );
OA21x2_ASAP7_75t_L g214 ( .A1(n_202), .A2(n_215), .B(n_224), .Y(n_214) );
OA21x2_ASAP7_75t_L g234 ( .A1(n_202), .A2(n_235), .B(n_243), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_202), .A2(n_472), .B(n_475), .Y(n_471) );
INVx1_ASAP7_75t_L g502 ( .A(n_202), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_202), .A2(n_539), .B(n_540), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_203), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_213), .Y(n_203) );
AND2x2_ASAP7_75t_L g406 ( .A(n_204), .B(n_403), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_204), .B(n_388), .Y(n_438) );
BUFx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g337 ( .A(n_205), .B(n_261), .Y(n_337) );
AND2x2_ASAP7_75t_L g386 ( .A(n_205), .B(n_232), .Y(n_386) );
INVx1_ASAP7_75t_L g432 ( .A(n_205), .Y(n_432) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_206), .Y(n_245) );
AND2x2_ASAP7_75t_L g287 ( .A(n_206), .B(n_261), .Y(n_287) );
INVx1_ASAP7_75t_L g304 ( .A(n_206), .Y(n_304) );
AND2x2_ASAP7_75t_L g310 ( .A(n_206), .B(n_225), .Y(n_310) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_210), .Y(n_485) );
INVx2_ASAP7_75t_L g513 ( .A(n_210), .Y(n_513) );
INVx1_ASAP7_75t_L g499 ( .A(n_212), .Y(n_499) );
AND2x2_ASAP7_75t_L g378 ( .A(n_213), .B(n_286), .Y(n_378) );
INVx2_ASAP7_75t_L g443 ( .A(n_213), .Y(n_443) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_225), .Y(n_213) );
AND2x2_ASAP7_75t_L g260 ( .A(n_214), .B(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g273 ( .A(n_214), .B(n_233), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_214), .B(n_232), .Y(n_301) );
INVx1_ASAP7_75t_L g307 ( .A(n_214), .Y(n_307) );
INVx1_ASAP7_75t_L g324 ( .A(n_214), .Y(n_324) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_214), .Y(n_336) );
INVx2_ASAP7_75t_L g404 ( .A(n_214), .Y(n_404) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B(n_219), .Y(n_216) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g261 ( .A(n_225), .Y(n_261) );
BUFx2_ASAP7_75t_L g358 ( .A(n_225), .Y(n_358) );
AND2x2_ASAP7_75t_L g403 ( .A(n_225), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_244), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_231), .B(n_340), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g426 ( .A1(n_231), .A2(n_402), .B(n_416), .Y(n_426) );
AND2x2_ASAP7_75t_L g451 ( .A(n_231), .B(n_337), .Y(n_451) );
BUFx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g373 ( .A(n_233), .Y(n_373) );
AND2x2_ASAP7_75t_L g402 ( .A(n_233), .B(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_234), .Y(n_286) );
INVx2_ASAP7_75t_L g305 ( .A(n_234), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_234), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
INVx2_ASAP7_75t_L g259 ( .A(n_245), .Y(n_259) );
OR2x2_ASAP7_75t_L g272 ( .A(n_245), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g340 ( .A(n_245), .B(n_336), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_245), .B(n_436), .Y(n_435) );
OR2x2_ASAP7_75t_L g441 ( .A(n_245), .B(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_245), .B(n_378), .Y(n_453) );
AND2x2_ASAP7_75t_L g332 ( .A(n_246), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g355 ( .A(n_246), .B(n_248), .Y(n_355) );
INVx2_ASAP7_75t_L g267 ( .A(n_247), .Y(n_267) );
AND2x2_ASAP7_75t_L g295 ( .A(n_247), .B(n_268), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_247), .B(n_320), .Y(n_376) );
AND2x2_ASAP7_75t_L g290 ( .A(n_248), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g437 ( .A(n_248), .Y(n_437) );
AND2x2_ASAP7_75t_L g449 ( .A(n_248), .B(n_312), .Y(n_449) );
AND2x2_ASAP7_75t_L g275 ( .A(n_249), .B(n_265), .Y(n_275) );
INVx1_ASAP7_75t_L g370 ( .A(n_249), .Y(n_370) );
AO21x1_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_251), .B(n_254), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_250), .B(n_489), .Y(n_488) );
INVx3_ASAP7_75t_L g505 ( .A(n_250), .Y(n_505) );
AO21x2_ASAP7_75t_L g517 ( .A1(n_250), .A2(n_518), .B(n_525), .Y(n_517) );
AO21x2_ASAP7_75t_L g573 ( .A1(n_250), .A2(n_574), .B(n_581), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_250), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x4_ASAP7_75t_L g268 ( .A(n_255), .B(n_269), .Y(n_268) );
INVxp67_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_262), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_259), .B(n_306), .Y(n_315) );
OR2x2_ASAP7_75t_L g447 ( .A(n_259), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g364 ( .A(n_260), .B(n_305), .Y(n_364) );
AND2x2_ASAP7_75t_L g372 ( .A(n_260), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g431 ( .A(n_260), .B(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g455 ( .A(n_260), .B(n_302), .Y(n_455) );
NOR2xp67_ASAP7_75t_L g413 ( .A(n_261), .B(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g442 ( .A(n_261), .B(n_305), .Y(n_442) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2x1p5_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
AND2x2_ASAP7_75t_L g294 ( .A(n_264), .B(n_295), .Y(n_294) );
INVxp67_ASAP7_75t_L g456 ( .A(n_264), .Y(n_456) );
NOR2x1_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVx1_ASAP7_75t_L g291 ( .A(n_267), .Y(n_291) );
AND2x2_ASAP7_75t_L g342 ( .A(n_267), .B(n_275), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_267), .B(n_410), .Y(n_436) );
INVx2_ASAP7_75t_L g281 ( .A(n_268), .Y(n_281) );
INVx3_ASAP7_75t_L g333 ( .A(n_268), .Y(n_333) );
OR2x2_ASAP7_75t_L g361 ( .A(n_268), .B(n_362), .Y(n_361) );
AOI311xp33_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_274), .A3(n_276), .B(n_277), .C(n_288), .Y(n_270) );
O2A1O1Ixp33_ASAP7_75t_L g308 ( .A1(n_271), .A2(n_309), .B(n_311), .C(n_313), .Y(n_308) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_SL g293 ( .A(n_273), .Y(n_293) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g311 ( .A(n_275), .B(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_275), .B(n_291), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_275), .B(n_276), .Y(n_444) );
AND2x2_ASAP7_75t_L g366 ( .A(n_276), .B(n_280), .Y(n_366) );
AOI21xp33_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_282), .B(n_283), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g424 ( .A(n_280), .B(n_312), .Y(n_424) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_281), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g318 ( .A(n_281), .Y(n_318) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
AND2x2_ASAP7_75t_L g309 ( .A(n_285), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g354 ( .A(n_287), .Y(n_354) );
AND2x4_ASAP7_75t_L g416 ( .A(n_287), .B(n_385), .Y(n_416) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AOI222xp33_ASAP7_75t_L g367 ( .A1(n_290), .A2(n_356), .B1(n_368), .B2(n_372), .C1(n_374), .C2(n_378), .Y(n_367) );
A2O1A1Ixp33_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_294), .B(n_296), .C(n_299), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_293), .B(n_337), .Y(n_360) );
INVx1_ASAP7_75t_L g382 ( .A(n_295), .Y(n_382) );
INVx1_ASAP7_75t_L g316 ( .A(n_297), .Y(n_316) );
OR2x2_ASAP7_75t_L g381 ( .A(n_298), .B(n_382), .Y(n_381) );
OAI21xp33_ASAP7_75t_SL g299 ( .A1(n_300), .A2(n_302), .B(n_306), .Y(n_299) );
NAND3xp33_ASAP7_75t_L g317 ( .A(n_300), .B(n_318), .C(n_319), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_300), .A2(n_337), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_304), .Y(n_357) );
AND2x2_ASAP7_75t_SL g323 ( .A(n_305), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g414 ( .A(n_305), .Y(n_414) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_305), .Y(n_430) );
INVx2_ASAP7_75t_L g388 ( .A(n_306), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_310), .B(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g362 ( .A(n_312), .Y(n_362) );
OAI221xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_316), .B1(n_317), .B2(n_321), .C(n_322), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_316), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_SL g450 ( .A(n_316), .Y(n_450) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g331 ( .A(n_323), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_323), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g389 ( .A(n_323), .B(n_337), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_323), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g422 ( .A(n_323), .B(n_357), .Y(n_422) );
BUFx3_ASAP7_75t_L g385 ( .A(n_324), .Y(n_385) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND5xp2_ASAP7_75t_L g327 ( .A(n_328), .B(n_346), .C(n_367), .D(n_379), .E(n_394), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AOI32xp33_ASAP7_75t_L g419 ( .A1(n_331), .A2(n_358), .A3(n_374), .B1(n_420), .B2(n_422), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_333), .B(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g343 ( .A(n_337), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_341), .B1(n_343), .B2(n_344), .Y(n_338) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
AOI221xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_353), .B1(n_355), .B2(n_356), .C(n_359), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g418 ( .A(n_350), .B(n_369), .Y(n_418) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AOI221xp5_ASAP7_75t_L g433 ( .A1(n_355), .A2(n_416), .B1(n_434), .B2(n_439), .C(n_440), .Y(n_433) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
INVx2_ASAP7_75t_L g399 ( .A(n_358), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_361), .B1(n_363), .B2(n_365), .Y(n_359) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
INVx1_ASAP7_75t_L g377 ( .A(n_369), .Y(n_377) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
AOI222xp33_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_383), .B1(n_387), .B2(n_388), .C1(n_389), .C2(n_390), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_386), .Y(n_383) );
INVxp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OAI22xp33_ASAP7_75t_L g434 ( .A1(n_388), .A2(n_435), .B1(n_437), .B2(n_438), .Y(n_434) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
AOI21xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_397), .B(n_400), .Y(n_394) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AOI21xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_405), .B(n_407), .Y(n_400) );
INVx2_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g448 ( .A(n_403), .Y(n_448) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
A2O1A1Ixp33_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_415), .B(n_417), .C(n_419), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AOI211xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_425), .B(n_427), .C(n_452), .Y(n_423) );
CKINVDCx16_ASAP7_75t_R g428 ( .A(n_424), .Y(n_428) );
INVxp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OAI211xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_429), .B(n_433), .C(n_445), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
AOI21xp33_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_443), .B(n_444), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_449), .B1(n_450), .B2(n_451), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AOI21xp33_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_454), .B(n_456), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g753 ( .A(n_465), .Y(n_753) );
OR3x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_665), .C(n_708), .Y(n_465) );
NAND5xp2_ASAP7_75t_L g466 ( .A(n_467), .B(n_592), .C(n_622), .D(n_639), .E(n_654), .Y(n_466) );
AOI221xp5_ASAP7_75t_SL g467 ( .A1(n_468), .A2(n_515), .B1(n_555), .B2(n_561), .C(n_565), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_490), .Y(n_468) );
OR2x2_ASAP7_75t_L g570 ( .A(n_469), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g609 ( .A(n_469), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g627 ( .A(n_469), .B(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_469), .B(n_563), .Y(n_644) );
OR2x2_ASAP7_75t_L g656 ( .A(n_469), .B(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_469), .B(n_615), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_469), .B(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_469), .B(n_593), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_469), .B(n_601), .Y(n_707) );
AND2x2_ASAP7_75t_L g739 ( .A(n_469), .B(n_503), .Y(n_739) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_469), .Y(n_747) );
INVx5_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_470), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g567 ( .A(n_470), .B(n_545), .Y(n_567) );
BUFx2_ASAP7_75t_L g589 ( .A(n_470), .Y(n_589) );
AND2x2_ASAP7_75t_L g618 ( .A(n_470), .B(n_491), .Y(n_618) );
AND2x2_ASAP7_75t_L g673 ( .A(n_470), .B(n_571), .Y(n_673) );
OR2x6_ASAP7_75t_L g470 ( .A(n_471), .B(n_488), .Y(n_470) );
BUFx2_ASAP7_75t_L g494 ( .A(n_473), .Y(n_494) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_SL g507 ( .A1(n_477), .A2(n_487), .B(n_508), .C(n_509), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_L g549 ( .A1(n_477), .A2(n_487), .B(n_550), .C(n_551), .Y(n_549) );
INVx5_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_482), .B(n_484), .C(n_485), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_L g541 ( .A1(n_482), .A2(n_485), .B(n_542), .C(n_543), .Y(n_541) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_490), .B(n_627), .Y(n_636) );
OAI32xp33_ASAP7_75t_L g650 ( .A1(n_490), .A2(n_586), .A3(n_651), .B1(n_652), .B2(n_653), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_490), .B(n_652), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_490), .B(n_570), .Y(n_693) );
INVx1_ASAP7_75t_SL g722 ( .A(n_490), .Y(n_722) );
NAND4xp25_ASAP7_75t_L g731 ( .A(n_490), .B(n_517), .C(n_673), .D(n_732), .Y(n_731) );
AND2x4_ASAP7_75t_L g490 ( .A(n_491), .B(n_503), .Y(n_490) );
INVx5_ASAP7_75t_L g564 ( .A(n_491), .Y(n_564) );
AND2x2_ASAP7_75t_L g593 ( .A(n_491), .B(n_504), .Y(n_593) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_491), .Y(n_672) );
AND2x2_ASAP7_75t_L g742 ( .A(n_491), .B(n_689), .Y(n_742) );
OR2x6_ASAP7_75t_L g491 ( .A(n_492), .B(n_500), .Y(n_491) );
AOI21xp5_ASAP7_75t_SL g492 ( .A1(n_493), .A2(n_495), .B(n_499), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
AND2x4_ASAP7_75t_L g615 ( .A(n_503), .B(n_564), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_503), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g649 ( .A(n_503), .B(n_571), .Y(n_649) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g563 ( .A(n_504), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g601 ( .A(n_504), .B(n_573), .Y(n_601) );
AND2x2_ASAP7_75t_L g610 ( .A(n_504), .B(n_572), .Y(n_610) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_506), .B(n_514), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
AOI222xp33_ASAP7_75t_L g678 ( .A1(n_515), .A2(n_679), .B1(n_681), .B2(n_683), .C1(n_686), .C2(n_687), .Y(n_678) );
AND2x4_ASAP7_75t_L g515 ( .A(n_516), .B(n_534), .Y(n_515) );
AND2x2_ASAP7_75t_L g611 ( .A(n_516), .B(n_612), .Y(n_611) );
NAND3xp33_ASAP7_75t_L g728 ( .A(n_516), .B(n_589), .C(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_527), .Y(n_516) );
INVx5_ASAP7_75t_SL g560 ( .A(n_517), .Y(n_560) );
OAI322xp33_ASAP7_75t_L g565 ( .A1(n_517), .A2(n_566), .A3(n_568), .B1(n_569), .B2(n_583), .C1(n_586), .C2(n_588), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_517), .B(n_558), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_517), .B(n_546), .Y(n_737) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_520), .B(n_521), .Y(n_518) );
INVx2_ASAP7_75t_L g558 ( .A(n_527), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_527), .B(n_536), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_534), .B(n_596), .Y(n_651) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OR2x2_ASAP7_75t_L g630 ( .A(n_535), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_545), .Y(n_535) );
OR2x2_ASAP7_75t_L g559 ( .A(n_536), .B(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_536), .B(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g598 ( .A(n_536), .B(n_546), .Y(n_598) );
AND2x2_ASAP7_75t_L g621 ( .A(n_536), .B(n_558), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_536), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g637 ( .A(n_536), .B(n_596), .Y(n_637) );
AND2x2_ASAP7_75t_L g645 ( .A(n_536), .B(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_536), .B(n_605), .Y(n_695) );
INVx5_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g585 ( .A(n_537), .B(n_560), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_537), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g612 ( .A(n_537), .B(n_546), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_537), .B(n_659), .Y(n_700) );
OR2x2_ASAP7_75t_L g716 ( .A(n_537), .B(n_660), .Y(n_716) );
AND2x2_ASAP7_75t_SL g723 ( .A(n_537), .B(n_677), .Y(n_723) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_537), .Y(n_730) );
OR2x6_ASAP7_75t_L g537 ( .A(n_538), .B(n_544), .Y(n_537) );
AND2x2_ASAP7_75t_L g584 ( .A(n_545), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g634 ( .A(n_545), .B(n_558), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_545), .B(n_560), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_545), .B(n_596), .Y(n_718) );
INVx3_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_546), .B(n_560), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_546), .B(n_558), .Y(n_606) );
OR2x2_ASAP7_75t_L g660 ( .A(n_546), .B(n_558), .Y(n_660) );
AND2x2_ASAP7_75t_L g677 ( .A(n_546), .B(n_557), .Y(n_677) );
INVxp67_ASAP7_75t_L g699 ( .A(n_546), .Y(n_699) );
AND2x2_ASAP7_75t_L g726 ( .A(n_546), .B(n_596), .Y(n_726) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_546), .Y(n_733) );
OA21x2_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B(n_554), .Y(n_546) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_559), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_557), .B(n_607), .Y(n_680) );
INVx1_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g596 ( .A(n_558), .B(n_560), .Y(n_596) );
OR2x2_ASAP7_75t_L g663 ( .A(n_558), .B(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g607 ( .A(n_559), .Y(n_607) );
OR2x2_ASAP7_75t_L g668 ( .A(n_559), .B(n_660), .Y(n_668) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g568 ( .A(n_563), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_563), .B(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_L g569 ( .A(n_564), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_564), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_564), .B(n_571), .Y(n_603) );
INVx2_ASAP7_75t_L g648 ( .A(n_564), .Y(n_648) );
AND2x2_ASAP7_75t_L g661 ( .A(n_564), .B(n_601), .Y(n_661) );
AND2x2_ASAP7_75t_L g686 ( .A(n_564), .B(n_610), .Y(n_686) );
INVx1_ASAP7_75t_L g638 ( .A(n_569), .Y(n_638) );
INVx2_ASAP7_75t_SL g625 ( .A(n_570), .Y(n_625) );
INVx1_ASAP7_75t_L g628 ( .A(n_571), .Y(n_628) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_572), .Y(n_591) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
BUFx2_ASAP7_75t_L g689 ( .A(n_573), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_580), .Y(n_574) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g658 ( .A(n_585), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g664 ( .A(n_585), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_585), .A2(n_667), .B1(n_669), .B2(n_674), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_585), .B(n_677), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_586), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_SL g620 ( .A(n_587), .Y(n_620) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
OR2x2_ASAP7_75t_L g602 ( .A(n_589), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_589), .B(n_593), .Y(n_653) );
AND2x2_ASAP7_75t_L g676 ( .A(n_589), .B(n_677), .Y(n_676) );
BUFx2_ASAP7_75t_L g652 ( .A(n_591), .Y(n_652) );
AOI211xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .B(n_599), .C(n_613), .Y(n_592) );
INVx1_ASAP7_75t_L g616 ( .A(n_593), .Y(n_616) );
OAI221xp5_ASAP7_75t_SL g724 ( .A1(n_593), .A2(n_725), .B1(n_727), .B2(n_728), .C(n_731), .Y(n_724) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
INVx1_ASAP7_75t_L g743 ( .A(n_596), .Y(n_743) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g692 ( .A(n_598), .B(n_631), .Y(n_692) );
A2O1A1Ixp33_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_602), .B(n_604), .C(n_608), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
OAI32xp33_ASAP7_75t_L g717 ( .A1(n_606), .A2(n_607), .A3(n_670), .B1(n_707), .B2(n_718), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .Y(n_608) );
AND2x2_ASAP7_75t_L g749 ( .A(n_609), .B(n_648), .Y(n_749) );
AND2x2_ASAP7_75t_L g696 ( .A(n_610), .B(n_648), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_610), .B(n_618), .Y(n_714) );
AOI31xp33_ASAP7_75t_SL g613 ( .A1(n_614), .A2(n_616), .A3(n_617), .B(n_619), .Y(n_613) );
INVxp67_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_615), .B(n_627), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_615), .B(n_625), .Y(n_712) );
AOI221xp5_ASAP7_75t_L g734 ( .A1(n_615), .A2(n_645), .B1(n_735), .B2(n_738), .C(n_740), .Y(n_734) );
CKINVDCx16_ASAP7_75t_R g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
AND2x2_ASAP7_75t_L g640 ( .A(n_620), .B(n_641), .Y(n_640) );
AOI222xp33_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_629), .B1(n_632), .B2(n_635), .C1(n_637), .C2(n_638), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_624), .B(n_626), .Y(n_623) );
INVx1_ASAP7_75t_L g705 ( .A(n_624), .Y(n_705) );
INVx1_ASAP7_75t_L g727 ( .A(n_627), .Y(n_727) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_630), .A2(n_741), .B1(n_743), .B2(n_744), .Y(n_740) );
INVx1_ASAP7_75t_L g646 ( .A(n_631), .Y(n_646) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_643), .B1(n_645), .B2(n_647), .C(n_650), .Y(n_639) );
INVx1_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g684 ( .A(n_642), .B(n_685), .Y(n_684) );
OR2x2_ASAP7_75t_L g736 ( .A(n_642), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g711 ( .A(n_647), .Y(n_711) );
AND2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
INVx1_ASAP7_75t_L g675 ( .A(n_648), .Y(n_675) );
INVx1_ASAP7_75t_L g657 ( .A(n_649), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_652), .B(n_739), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_658), .B1(n_661), .B2(n_662), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g748 ( .A(n_661), .Y(n_748) );
INVxp33_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_663), .B(n_707), .Y(n_706) );
OAI32xp33_ASAP7_75t_L g697 ( .A1(n_664), .A2(n_698), .A3(n_699), .B1(n_700), .B2(n_701), .Y(n_697) );
NAND4xp25_ASAP7_75t_L g665 ( .A(n_666), .B(n_678), .C(n_690), .D(n_702), .Y(n_665) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
NAND2xp33_ASAP7_75t_SL g669 ( .A(n_670), .B(n_671), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_673), .B(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
CKINVDCx16_ASAP7_75t_R g683 ( .A(n_684), .Y(n_683) );
AOI221xp5_ASAP7_75t_L g719 ( .A1(n_687), .A2(n_703), .B1(n_720), .B2(n_723), .C(n_724), .Y(n_719) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g738 ( .A(n_689), .B(n_739), .Y(n_738) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_693), .B1(n_694), .B2(n_696), .C(n_697), .Y(n_690) );
INVx1_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_699), .B(n_730), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_705), .B(n_706), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NAND4xp25_ASAP7_75t_L g708 ( .A(n_709), .B(n_719), .C(n_734), .D(n_745), .Y(n_708) );
O2A1O1Ixp33_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_713), .B(n_715), .C(n_717), .Y(n_709) );
NAND2xp5_ASAP7_75t_SL g710 ( .A(n_711), .B(n_712), .Y(n_710) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVxp67_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g750 ( .A(n_737), .Y(n_750) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
OAI21xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_749), .B(n_750), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
BUFx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g770 ( .A(n_762), .Y(n_770) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_765), .Y(n_768) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
endmodule