module fake_jpeg_789_n_501 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_501);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_501;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_16),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_47),
.B(n_50),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_13),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_51),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_52),
.Y(n_131)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_54),
.Y(n_136)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_23),
.B(n_13),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_56),
.B(n_60),
.Y(n_116)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_58),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_23),
.B(n_0),
.Y(n_60)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_62),
.Y(n_114)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_17),
.B(n_0),
.Y(n_64)
);

NAND2xp33_ASAP7_75t_SL g154 ( 
.A(n_64),
.B(n_3),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_24),
.B(n_1),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_67),
.B(n_74),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_24),
.B(n_1),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_79),
.Y(n_142)
);

BUFx4f_ASAP7_75t_SL g80 ( 
.A(n_42),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_86),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_82),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_83),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_35),
.B(n_1),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_85),
.B(n_89),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_44),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_44),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_88),
.B(n_92),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_35),
.B(n_1),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_38),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_30),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_18),
.Y(n_94)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

BUFx4f_ASAP7_75t_SL g96 ( 
.A(n_41),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_96),
.B(n_39),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_58),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_99),
.B(n_143),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_46),
.A2(n_43),
.B1(n_41),
.B2(n_44),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_103),
.A2(n_109),
.B1(n_115),
.B2(n_121),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_21),
.B1(n_29),
.B2(n_41),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_45),
.A2(n_21),
.B1(n_44),
.B2(n_43),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_65),
.A2(n_43),
.B1(n_34),
.B2(n_36),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_68),
.A2(n_43),
.B1(n_37),
.B2(n_34),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_123),
.A2(n_147),
.B1(n_91),
.B2(n_87),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_50),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_134),
.A2(n_62),
.B1(n_79),
.B2(n_81),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_77),
.A2(n_69),
.B1(n_71),
.B2(n_37),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_141),
.A2(n_70),
.B1(n_95),
.B2(n_93),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_64),
.B(n_48),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_49),
.A2(n_36),
.B1(n_33),
.B2(n_32),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_58),
.B(n_31),
.C(n_22),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_154),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_SL g150 ( 
.A1(n_61),
.A2(n_22),
.B(n_39),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_150),
.B(n_39),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_48),
.B(n_2),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_80),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_155),
.Y(n_163)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_156),
.Y(n_220)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_157),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_140),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_159),
.B(n_161),
.Y(n_235)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_160),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_119),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_162),
.B(n_167),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_164),
.B(n_175),
.Y(n_237)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_165),
.Y(n_228)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_100),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_166),
.Y(n_236)
);

AND2x2_ASAP7_75t_SL g167 ( 
.A(n_107),
.B(n_120),
.Y(n_167)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_132),
.Y(n_168)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_168),
.Y(n_231)
);

BUFx2_ASAP7_75t_SL g169 ( 
.A(n_137),
.Y(n_169)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_169),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_113),
.B(n_61),
.Y(n_171)
);

AND2x2_ASAP7_75t_SL g203 ( 
.A(n_171),
.B(n_200),
.Y(n_203)
);

AND2x4_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_80),
.Y(n_172)
);

NAND2xp33_ASAP7_75t_SL g209 ( 
.A(n_172),
.B(n_197),
.Y(n_209)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_111),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_173),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_112),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_174),
.Y(n_229)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_132),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_177),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_104),
.B(n_96),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_178),
.B(n_182),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_144),
.B(n_22),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_180),
.Y(n_214)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_112),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_181),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_110),
.B(n_96),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_146),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_190),
.Y(n_226)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_117),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_185),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_101),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_186),
.Y(n_219)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_135),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_187),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_103),
.A2(n_51),
.B1(n_54),
.B2(n_52),
.Y(n_188)
);

A2O1A1Ixp33_ASAP7_75t_SL g204 ( 
.A1(n_188),
.A2(n_194),
.B(n_201),
.C(n_109),
.Y(n_204)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_101),
.Y(n_189)
);

INVx8_ASAP7_75t_L g233 ( 
.A(n_189),
.Y(n_233)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

BUFx8_ASAP7_75t_L g191 ( 
.A(n_105),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_193),
.Y(n_230)
);

NAND3xp33_ASAP7_75t_SL g193 ( 
.A(n_116),
.B(n_22),
.C(n_83),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_195),
.A2(n_202),
.B1(n_115),
.B2(n_121),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_98),
.B(n_65),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_105),
.Y(n_222)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_125),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_126),
.A2(n_84),
.B1(n_82),
.B2(n_76),
.Y(n_198)
);

NAND2xp33_ASAP7_75t_SL g221 ( 
.A(n_198),
.B(n_199),
.Y(n_221)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_149),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_108),
.B(n_73),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_124),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_123),
.A2(n_72),
.B1(n_22),
.B2(n_39),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_204),
.B(n_216),
.Y(n_244)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_207),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_194),
.A2(n_102),
.B(n_153),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_212),
.A2(n_191),
.B(n_164),
.Y(n_264)
);

FAx1_ASAP7_75t_SL g213 ( 
.A(n_179),
.B(n_153),
.CI(n_22),
.CON(n_213),
.SN(n_213)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_213),
.B(n_230),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_195),
.A2(n_125),
.B1(n_145),
.B2(n_127),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_158),
.A2(n_151),
.B1(n_145),
.B2(n_127),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_218),
.B(n_114),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_222),
.B(n_180),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_204),
.A2(n_170),
.B1(n_158),
.B2(n_163),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_238),
.A2(n_255),
.B1(n_256),
.B2(n_261),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_203),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_240),
.Y(n_268)
);

AND2x6_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_161),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_237),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_241),
.B(n_245),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_158),
.C(n_171),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_248),
.C(n_250),
.Y(n_270)
);

NAND3xp33_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_171),
.C(n_182),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_159),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_246),
.B(n_265),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_203),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_253),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_212),
.B(n_178),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_209),
.A2(n_172),
.B(n_157),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_249),
.A2(n_264),
.B(n_206),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_166),
.C(n_165),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_227),
.Y(n_251)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

AOI21xp33_ASAP7_75t_L g252 ( 
.A1(n_210),
.A2(n_192),
.B(n_172),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_252),
.A2(n_230),
.B(n_204),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_215),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_205),
.A2(n_188),
.B1(n_167),
.B2(n_177),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_205),
.A2(n_167),
.B1(n_200),
.B2(n_186),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_258),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_209),
.A2(n_191),
.B(n_172),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_259),
.A2(n_230),
.B(n_206),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_232),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_236),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_204),
.A2(n_200),
.B1(n_189),
.B2(n_124),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_262),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_263),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_225),
.B(n_160),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_203),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_273),
.A2(n_276),
.B(n_286),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_274),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_246),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_275),
.B(n_280),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_203),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_277),
.B(n_295),
.C(n_248),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_265),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_251),
.Y(n_282)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_282),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_250),
.B(n_219),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_287),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_258),
.A2(n_235),
.B(n_204),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_245),
.B(n_219),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_254),
.Y(n_288)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_288),
.Y(n_300)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_289),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_243),
.A2(n_205),
.B1(n_226),
.B2(n_213),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_290),
.A2(n_248),
.B1(n_266),
.B2(n_264),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_238),
.A2(n_221),
.B(n_217),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_291),
.B(n_293),
.Y(n_311)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_262),
.Y(n_292)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_292),
.Y(n_313)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_262),
.Y(n_294)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_294),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_242),
.B(n_223),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_279),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_297),
.B(n_301),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_289),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_269),
.A2(n_243),
.B1(n_244),
.B2(n_240),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_302),
.A2(n_310),
.B1(n_312),
.B2(n_319),
.Y(n_329)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_281),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_304),
.B(n_306),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_305),
.B(n_307),
.C(n_318),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_275),
.B(n_253),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_270),
.B(n_247),
.C(n_239),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_309),
.B(n_277),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_269),
.A2(n_244),
.B1(n_261),
.B2(n_255),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_274),
.A2(n_286),
.B1(n_290),
.B2(n_279),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_283),
.B(n_260),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_314),
.B(n_315),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_287),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_278),
.Y(n_316)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_316),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_278),
.Y(n_317)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_317),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_270),
.B(n_249),
.C(n_259),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_272),
.A2(n_226),
.B1(n_263),
.B2(n_240),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_268),
.A2(n_256),
.B1(n_207),
.B2(n_226),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_320),
.A2(n_322),
.B1(n_293),
.B2(n_280),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_272),
.A2(n_252),
.B1(n_221),
.B2(n_217),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_284),
.B(n_273),
.Y(n_323)
);

INVxp33_ASAP7_75t_L g338 ( 
.A(n_323),
.Y(n_338)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_267),
.Y(n_324)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_324),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_305),
.B(n_295),
.Y(n_327)
);

MAJx2_ASAP7_75t_L g356 ( 
.A(n_327),
.B(n_349),
.C(n_350),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_328),
.B(n_341),
.Y(n_360)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_324),
.Y(n_333)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_333),
.Y(n_361)
);

OAI21x1_ASAP7_75t_L g335 ( 
.A1(n_298),
.A2(n_284),
.B(n_268),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_335),
.B(n_339),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_336),
.A2(n_348),
.B1(n_227),
.B2(n_223),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_315),
.A2(n_276),
.B(n_291),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_299),
.Y(n_340)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_340),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_307),
.B(n_298),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_318),
.B(n_277),
.C(n_285),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_343),
.C(n_303),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_311),
.B(n_283),
.C(n_267),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_299),
.Y(n_344)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_344),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_296),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_345),
.B(n_347),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_309),
.B(n_271),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_346),
.B(n_351),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_323),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_302),
.A2(n_310),
.B1(n_297),
.B2(n_319),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_322),
.B(n_288),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_312),
.B(n_282),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_323),
.B(n_271),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_300),
.Y(n_352)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_352),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_308),
.B(n_303),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_353),
.B(n_346),
.Y(n_379)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_300),
.Y(n_354)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_354),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_357),
.B(n_379),
.Y(n_404)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_332),
.Y(n_359)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_359),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_338),
.A2(n_321),
.B(n_320),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_363),
.A2(n_371),
.B(n_378),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_348),
.A2(n_329),
.B1(n_336),
.B2(n_338),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_365),
.A2(n_370),
.B1(n_337),
.B2(n_216),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_328),
.B(n_321),
.Y(n_368)
);

OAI322xp33_ASAP7_75t_L g387 ( 
.A1(n_368),
.A2(n_358),
.A3(n_356),
.B1(n_379),
.B2(n_367),
.C1(n_374),
.C2(n_377),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_343),
.B(n_296),
.Y(n_369)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_369),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_329),
.A2(n_355),
.B1(n_308),
.B2(n_330),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_351),
.A2(n_325),
.B(n_313),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_334),
.B(n_304),
.Y(n_372)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_372),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_353),
.Y(n_374)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_374),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_327),
.B(n_325),
.C(n_313),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_375),
.B(n_383),
.C(n_368),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_326),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_L g401 ( 
.A1(n_376),
.A2(n_380),
.B1(n_211),
.B2(n_176),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_349),
.A2(n_294),
.B(n_292),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_331),
.B(n_281),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_341),
.B(n_218),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_381),
.B(n_185),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_382),
.A2(n_224),
.B1(n_228),
.B2(n_211),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_342),
.B(n_224),
.C(n_228),
.Y(n_383)
);

FAx1_ASAP7_75t_SL g384 ( 
.A(n_356),
.B(n_350),
.CI(n_337),
.CON(n_384),
.SN(n_384)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_384),
.B(n_387),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_388),
.A2(n_391),
.B1(n_408),
.B2(n_136),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_389),
.B(n_407),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_375),
.B(n_229),
.C(n_214),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_390),
.B(n_399),
.Y(n_417)
);

BUFx12f_ASAP7_75t_SL g393 ( 
.A(n_370),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_393),
.A2(n_394),
.B(n_395),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_363),
.A2(n_365),
.B(n_371),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_378),
.A2(n_229),
.B(n_208),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_380),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_396),
.B(n_403),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_367),
.A2(n_229),
.B(n_236),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_398),
.A2(n_183),
.B(n_173),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_357),
.B(n_220),
.C(n_208),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_360),
.B(n_220),
.C(n_234),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_400),
.B(n_407),
.Y(n_421)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_401),
.Y(n_416)
);

INVx13_ASAP7_75t_L g402 ( 
.A(n_361),
.Y(n_402)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_402),
.Y(n_426)
);

AOI322xp5_ASAP7_75t_SL g403 ( 
.A1(n_372),
.A2(n_201),
.A3(n_181),
.B1(n_174),
.B2(n_231),
.C1(n_233),
.C2(n_137),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_359),
.A2(n_231),
.B1(n_233),
.B2(n_168),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_405),
.A2(n_114),
.B1(n_128),
.B2(n_131),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_360),
.B(n_197),
.C(n_190),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_381),
.A2(n_383),
.B1(n_373),
.B2(n_366),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_409),
.Y(n_427)
);

CKINVDCx14_ASAP7_75t_R g410 ( 
.A(n_408),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_410),
.B(n_411),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_389),
.B(n_364),
.C(n_362),
.Y(n_411)
);

NOR2xp67_ASAP7_75t_SL g440 ( 
.A(n_412),
.B(n_423),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_413),
.B(n_395),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_156),
.C(n_199),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_415),
.B(n_419),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_406),
.B(n_187),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_388),
.Y(n_420)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_420),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_394),
.B(n_106),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_422),
.B(n_424),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_390),
.B(n_142),
.C(n_151),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_404),
.B(n_136),
.Y(n_424)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_385),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_428),
.B(n_385),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_429),
.B(n_431),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_400),
.B(n_128),
.C(n_97),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_430),
.B(n_398),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_412),
.B(n_386),
.C(n_397),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_432),
.B(n_439),
.Y(n_451)
);

OA21x2_ASAP7_75t_L g434 ( 
.A1(n_425),
.A2(n_386),
.B(n_393),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_434),
.Y(n_460)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_437),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_438),
.B(n_3),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_411),
.B(n_397),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_441),
.B(n_442),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_414),
.B(n_392),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_421),
.B(n_392),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_444),
.B(n_446),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_418),
.A2(n_384),
.B(n_402),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_445),
.A2(n_413),
.B(n_415),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_426),
.B(n_405),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_427),
.B(n_384),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_447),
.B(n_449),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_427),
.B(n_131),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_440),
.B(n_417),
.C(n_422),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_454),
.B(n_455),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_444),
.B(n_416),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_443),
.B(n_425),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_457),
.B(n_461),
.Y(n_473)
);

AO21x1_ASAP7_75t_L g471 ( 
.A1(n_458),
.A2(n_464),
.B(n_4),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_435),
.A2(n_429),
.B(n_423),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_459),
.A2(n_460),
.B(n_463),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_432),
.B(n_430),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_434),
.B(n_97),
.C(n_106),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_462),
.B(n_463),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_434),
.B(n_39),
.C(n_59),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_448),
.B(n_3),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_465),
.B(n_6),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_450),
.B(n_433),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g482 ( 
.A(n_466),
.B(n_468),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_453),
.B(n_436),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_451),
.B(n_436),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_469),
.B(n_472),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_452),
.A2(n_441),
.B(n_38),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_470),
.A2(n_477),
.B(n_7),
.Y(n_481)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_471),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_460),
.B(n_4),
.C(n_5),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_12),
.Y(n_474)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_474),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_476),
.B(n_478),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_454),
.B(n_7),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_473),
.B(n_464),
.C(n_8),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_479),
.B(n_9),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_481),
.B(n_487),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_466),
.B(n_7),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_484),
.A2(n_486),
.B(n_12),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_467),
.A2(n_7),
.B(n_8),
.Y(n_486)
);

O2A1O1Ixp33_ASAP7_75t_SL g488 ( 
.A1(n_482),
.A2(n_474),
.B(n_475),
.C(n_10),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_488),
.A2(n_483),
.B(n_480),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_484),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_489),
.B(n_490),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_491),
.B(n_492),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_485),
.B(n_8),
.C(n_9),
.Y(n_492)
);

OAI32xp33_ASAP7_75t_L g497 ( 
.A1(n_493),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_489),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_495),
.B(n_497),
.Y(n_498)
);

BUFx24_ASAP7_75t_SL g499 ( 
.A(n_494),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_499),
.Y(n_500)
);

A2O1A1Ixp33_ASAP7_75t_L g501 ( 
.A1(n_500),
.A2(n_498),
.B(n_496),
.C(n_10),
.Y(n_501)
);


endmodule