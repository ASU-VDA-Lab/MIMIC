module fake_jpeg_10892_n_641 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_641);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_641;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_544;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_5),
.B(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_17),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_59),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_60),
.B(n_66),
.Y(n_134)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_61),
.Y(n_148)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_63),
.Y(n_142)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_64),
.Y(n_136)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_65),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_9),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_67),
.Y(n_194)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_68),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_69),
.Y(n_144)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_71),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_72),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_73),
.Y(n_145)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_74),
.Y(n_163)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_75),
.Y(n_156)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_78),
.Y(n_164)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_79),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_81),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_82),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_83),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_20),
.B(n_18),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_84),
.B(n_88),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_86),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_87),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_25),
.B(n_9),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_90),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_91),
.Y(n_202)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_92),
.Y(n_157)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_93),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_31),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_94),
.B(n_106),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_95),
.Y(n_185)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_96),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g174 ( 
.A(n_98),
.Y(n_174)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_99),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_35),
.Y(n_100)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_100),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_29),
.Y(n_101)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_101),
.Y(n_171)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_39),
.Y(n_102)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_102),
.Y(n_195)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_103),
.Y(n_176)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_104),
.Y(n_178)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_27),
.Y(n_105)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_105),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_20),
.B(n_18),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_49),
.B(n_9),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_107),
.B(n_112),
.Y(n_188)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_31),
.Y(n_108)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_108),
.Y(n_173)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_109),
.Y(n_180)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_31),
.Y(n_110)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_110),
.Y(n_179)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_111),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_58),
.B(n_10),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_43),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_114),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_44),
.Y(n_115)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_115),
.Y(n_193)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_29),
.Y(n_116)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_116),
.Y(n_197)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_117),
.Y(n_186)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_27),
.Y(n_118)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_118),
.Y(n_212)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_119),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_44),
.Y(n_120)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_44),
.Y(n_121)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_121),
.Y(n_177)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_56),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_122),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_51),
.A2(n_18),
.B1(n_17),
.B2(n_16),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_123),
.A2(n_107),
.B(n_88),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_58),
.B(n_15),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_124),
.B(n_28),
.Y(n_214)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_43),
.Y(n_125)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_125),
.Y(n_199)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_44),
.Y(n_126)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_126),
.Y(n_203)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_43),
.Y(n_127)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_127),
.Y(n_217)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_46),
.Y(n_128)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_128),
.Y(n_218)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_45),
.Y(n_129)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_129),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_91),
.A2(n_72),
.B1(n_73),
.B2(n_51),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_133),
.A2(n_138),
.B1(n_154),
.B2(n_182),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_137),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_91),
.A2(n_29),
.B1(n_48),
.B2(n_54),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_60),
.B(n_56),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_139),
.Y(n_233)
);

OA22x2_ASAP7_75t_L g281 ( 
.A1(n_140),
.A2(n_146),
.B1(n_154),
.B2(n_138),
.Y(n_281)
);

O2A1O1Ixp33_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_56),
.B(n_23),
.C(n_36),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_66),
.B(n_40),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_153),
.B(n_162),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_79),
.A2(n_54),
.B1(n_48),
.B2(n_46),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_112),
.B(n_40),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_124),
.B(n_21),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_175),
.B(n_196),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_98),
.A2(n_46),
.B1(n_47),
.B2(n_30),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_111),
.A2(n_46),
.B1(n_47),
.B2(n_30),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_184),
.A2(n_208),
.B1(n_210),
.B2(n_213),
.Y(n_241)
);

AND2x2_ASAP7_75t_SL g190 ( 
.A(n_125),
.B(n_56),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_190),
.B(n_121),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_114),
.B(n_37),
.Y(n_196)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_127),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_198),
.Y(n_252)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_128),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_207),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_101),
.A2(n_54),
.B1(n_48),
.B2(n_47),
.Y(n_208)
);

HAxp5_ASAP7_75t_SL g209 ( 
.A(n_69),
.B(n_21),
.CON(n_209),
.SN(n_209)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_209),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_71),
.A2(n_54),
.B1(n_48),
.B2(n_47),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_78),
.Y(n_211)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_211),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_82),
.A2(n_55),
.B1(n_45),
.B2(n_50),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_134),
.Y(n_234)
);

BUFx12_ASAP7_75t_L g215 ( 
.A(n_83),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_215),
.Y(n_269)
);

BUFx2_ASAP7_75t_SL g216 ( 
.A(n_86),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_216),
.Y(n_254)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_87),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_219),
.Y(n_286)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_97),
.Y(n_220)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_220),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_115),
.A2(n_23),
.B1(n_32),
.B2(n_36),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_37),
.B1(n_52),
.B2(n_2),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_137),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_222),
.B(n_225),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_144),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_223),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_215),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_130),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_226),
.B(n_243),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_146),
.A2(n_50),
.B1(n_55),
.B2(n_28),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_227),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_231),
.Y(n_320)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_159),
.Y(n_232)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_232),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_234),
.B(n_235),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_172),
.B(n_52),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_188),
.B(n_32),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_236),
.B(n_239),
.Y(n_302)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_206),
.Y(n_237)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_237),
.Y(n_300)
);

INVx11_ASAP7_75t_L g238 ( 
.A(n_168),
.Y(n_238)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_238),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_188),
.B(n_41),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_204),
.Y(n_240)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_240),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_139),
.B(n_120),
.C(n_41),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_242),
.B(n_260),
.C(n_276),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_136),
.Y(n_243)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_202),
.Y(n_244)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_244),
.Y(n_301)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_205),
.Y(n_245)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_245),
.Y(n_305)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_247),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_248),
.A2(n_266),
.B1(n_272),
.B2(n_278),
.Y(n_341)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_161),
.Y(n_249)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_249),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_134),
.B(n_0),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_250),
.B(n_271),
.Y(n_323)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_166),
.Y(n_251)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_251),
.Y(n_344)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_212),
.Y(n_253)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_253),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_194),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_255),
.B(n_259),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_133),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_256),
.B(n_170),
.Y(n_337)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_176),
.Y(n_257)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_257),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_144),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_258),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_195),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_150),
.B(n_17),
.C(n_15),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_172),
.B(n_15),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_261),
.B(n_284),
.Y(n_312)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_218),
.Y(n_262)
);

INVx5_ASAP7_75t_L g314 ( 
.A(n_262),
.Y(n_314)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_178),
.Y(n_263)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_263),
.Y(n_350)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_199),
.Y(n_264)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_264),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_160),
.Y(n_265)
);

INVx6_ASAP7_75t_L g304 ( 
.A(n_265),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_208),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_266)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_160),
.Y(n_267)
);

INVx5_ASAP7_75t_L g319 ( 
.A(n_267),
.Y(n_319)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_145),
.Y(n_270)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_270),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_150),
.B(n_151),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_221),
.A2(n_14),
.B1(n_11),
.B2(n_2),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_203),
.Y(n_274)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_274),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_190),
.B(n_0),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_132),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_277),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_210),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_142),
.B(n_3),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_279),
.B(n_174),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_164),
.Y(n_280)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_280),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_281),
.Y(n_335)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_171),
.Y(n_282)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_282),
.Y(n_348)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_180),
.Y(n_283)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_283),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_158),
.B(n_3),
.Y(n_284)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_185),
.Y(n_285)
);

BUFx24_ASAP7_75t_L g331 ( 
.A(n_285),
.Y(n_331)
);

O2A1O1Ixp33_ASAP7_75t_L g287 ( 
.A1(n_168),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_287)
);

A2O1A1Ixp33_ASAP7_75t_L g329 ( 
.A1(n_287),
.A2(n_187),
.B(n_200),
.C(n_156),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_213),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_288),
.A2(n_295),
.B1(n_297),
.B2(n_287),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_216),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_289),
.A2(n_291),
.B1(n_296),
.B2(n_298),
.Y(n_306)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_135),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_290),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_169),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_143),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_292),
.B(n_240),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_181),
.B(n_8),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_293),
.B(n_231),
.C(n_260),
.Y(n_352)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_186),
.Y(n_294)
);

INVx13_ASAP7_75t_L g330 ( 
.A(n_294),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_155),
.A2(n_8),
.B1(n_193),
.B2(n_141),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_177),
.A2(n_201),
.B1(n_189),
.B2(n_192),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_201),
.A2(n_189),
.B1(n_164),
.B2(n_192),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_191),
.A2(n_165),
.B1(n_163),
.B2(n_200),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_197),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_299),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_246),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_303),
.B(n_342),
.Y(n_387)
);

AOI32xp33_ASAP7_75t_L g310 ( 
.A1(n_271),
.A2(n_131),
.A3(n_147),
.B1(n_157),
.B2(n_149),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_310),
.A2(n_286),
.B(n_269),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_276),
.A2(n_148),
.B(n_152),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_317),
.A2(n_349),
.B(n_338),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_L g324 ( 
.A1(n_288),
.A2(n_241),
.B1(n_281),
.B2(n_230),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_324),
.A2(n_269),
.B1(n_262),
.B2(n_286),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_325),
.B(n_340),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_329),
.B(n_254),
.Y(n_366)
);

AO22x2_ASAP7_75t_L g333 ( 
.A1(n_281),
.A2(n_174),
.B1(n_183),
.B2(n_167),
.Y(n_333)
);

AO21x2_ASAP7_75t_SL g377 ( 
.A1(n_333),
.A2(n_254),
.B(n_268),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_337),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_250),
.B(n_173),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_338),
.B(n_349),
.C(n_313),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_281),
.A2(n_179),
.B1(n_191),
.B2(n_163),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_339),
.Y(n_369)
);

OR2x2_ASAP7_75t_L g340 ( 
.A(n_236),
.B(n_165),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_275),
.B(n_224),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_343),
.B(n_267),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_238),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_346),
.B(n_358),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_276),
.A2(n_231),
.B(n_242),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_351),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_352),
.B(n_237),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_224),
.B(n_239),
.Y(n_358)
);

OAI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_273),
.A2(n_233),
.B1(n_253),
.B2(n_247),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_359),
.A2(n_252),
.B1(n_268),
.B2(n_299),
.Y(n_391)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_304),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_360),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_361),
.A2(n_362),
.B(n_366),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_335),
.A2(n_290),
.B(n_285),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_335),
.A2(n_293),
.B1(n_279),
.B2(n_283),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_364),
.A2(n_365),
.B1(n_377),
.B2(n_356),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_320),
.A2(n_293),
.B1(n_274),
.B2(n_286),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_367),
.A2(n_373),
.B1(n_376),
.B2(n_390),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_328),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_368),
.B(n_384),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_353),
.Y(n_370)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_370),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_371),
.B(n_403),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_325),
.B(n_323),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_372),
.B(n_380),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_374),
.B(n_396),
.Y(n_416)
);

INVx3_ASAP7_75t_SL g375 ( 
.A(n_304),
.Y(n_375)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_375),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_341),
.A2(n_294),
.B1(n_264),
.B2(n_229),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_313),
.B(n_352),
.C(n_323),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_378),
.B(n_379),
.C(n_388),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_340),
.B(n_257),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_327),
.A2(n_322),
.B1(n_306),
.B2(n_333),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_382),
.A2(n_404),
.B1(n_345),
.B2(n_305),
.Y(n_419)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_309),
.Y(n_383)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_383),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_334),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_322),
.A2(n_244),
.B(n_245),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_385),
.A2(n_391),
.B(n_395),
.Y(n_439)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_309),
.Y(n_386)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_386),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_302),
.B(n_251),
.C(n_232),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_302),
.B(n_263),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_389),
.B(n_394),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_343),
.A2(n_223),
.B1(n_280),
.B2(n_265),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_341),
.A2(n_258),
.B1(n_229),
.B2(n_228),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_392),
.A2(n_399),
.B1(n_402),
.B2(n_376),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_318),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_393),
.B(n_406),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_311),
.B(n_249),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_327),
.A2(n_252),
.B(n_270),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_307),
.B(n_282),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_321),
.B(n_228),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_397),
.B(n_400),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_333),
.A2(n_317),
.B1(n_329),
.B2(n_312),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_321),
.B(n_303),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_333),
.A2(n_306),
.B1(n_346),
.B2(n_336),
.Y(n_402)
);

NAND2x1p5_ASAP7_75t_L g403 ( 
.A(n_333),
.B(n_308),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_SL g404 ( 
.A1(n_305),
.A2(n_319),
.B1(n_301),
.B2(n_314),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_332),
.B(n_356),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_405),
.B(n_393),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_331),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_374),
.B(n_332),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_409),
.B(n_415),
.C(n_432),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_410),
.A2(n_441),
.B1(n_367),
.B2(n_373),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_379),
.B(n_300),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_419),
.A2(n_422),
.B(n_391),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_368),
.B(n_355),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_420),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_384),
.B(n_301),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_421),
.Y(n_473)
);

AOI32xp33_ASAP7_75t_L g422 ( 
.A1(n_381),
.A2(n_331),
.A3(n_326),
.B1(n_300),
.B2(n_348),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_378),
.B(n_326),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_SL g474 ( 
.A(n_423),
.B(n_364),
.Y(n_474)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_400),
.Y(n_424)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_424),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_405),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_425),
.B(n_442),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_427),
.A2(n_444),
.B1(n_377),
.B2(n_369),
.Y(n_453)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_383),
.Y(n_428)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_428),
.Y(n_460)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_386),
.Y(n_429)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_429),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_372),
.B(n_348),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_361),
.B(n_331),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_434),
.B(n_381),
.C(n_371),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_436),
.B(n_438),
.Y(n_459)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_397),
.Y(n_437)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_437),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_389),
.B(n_344),
.Y(n_438)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_392),
.Y(n_440)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_440),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_382),
.A2(n_336),
.B1(n_319),
.B2(n_354),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_360),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_401),
.B(n_347),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_443),
.B(n_401),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_402),
.A2(n_354),
.B1(n_353),
.B2(n_314),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_412),
.B(n_396),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_446),
.B(n_452),
.C(n_471),
.Y(n_493)
);

BUFx24_ASAP7_75t_SL g449 ( 
.A(n_445),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_449),
.B(n_465),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_445),
.B(n_406),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_451),
.B(n_456),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_412),
.B(n_396),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_453),
.A2(n_413),
.B1(n_429),
.B2(n_428),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_454),
.A2(n_458),
.B1(n_461),
.B2(n_464),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_436),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_418),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_457),
.B(n_462),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_410),
.A2(n_367),
.B1(n_399),
.B2(n_390),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_441),
.A2(n_367),
.B1(n_366),
.B2(n_403),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_433),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_424),
.A2(n_403),
.B1(n_377),
.B2(n_380),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_425),
.B(n_394),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_435),
.A2(n_362),
.B(n_385),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_467),
.A2(n_468),
.B(n_451),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_435),
.A2(n_430),
.B(n_439),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_469),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_443),
.B(n_387),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_470),
.B(n_438),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_416),
.B(n_388),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_409),
.B(n_388),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_472),
.B(n_476),
.C(n_437),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_SL g485 ( 
.A(n_474),
.B(n_415),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_433),
.B(n_387),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_475),
.Y(n_510)
);

OR2x6_ASAP7_75t_L g513 ( 
.A(n_477),
.B(n_479),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_440),
.A2(n_403),
.B1(n_377),
.B2(n_398),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_478),
.A2(n_377),
.B1(n_427),
.B2(n_426),
.Y(n_486)
);

CKINVDCx14_ASAP7_75t_R g479 ( 
.A(n_431),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_430),
.A2(n_363),
.B(n_395),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_480),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_471),
.B(n_416),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_482),
.B(n_487),
.Y(n_528)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_484),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_SL g517 ( 
.A(n_485),
.B(n_489),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_486),
.A2(n_511),
.B1(n_450),
.B2(n_466),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_447),
.B(n_423),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_447),
.B(n_434),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_488),
.B(n_491),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_SL g489 ( 
.A(n_446),
.B(n_432),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_472),
.B(n_407),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_452),
.B(n_407),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_492),
.B(n_494),
.C(n_500),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_478),
.Y(n_496)
);

INVx1_ASAP7_75t_SL g543 ( 
.A(n_496),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_468),
.A2(n_419),
.B(n_431),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_497),
.Y(n_524)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_498),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_474),
.B(n_476),
.C(n_475),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_458),
.A2(n_426),
.B1(n_444),
.B2(n_439),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_501),
.A2(n_507),
.B1(n_509),
.B2(n_481),
.Y(n_519)
);

NAND2x1_ASAP7_75t_L g502 ( 
.A(n_467),
.B(n_422),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_502),
.B(n_512),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_505),
.A2(n_508),
.B1(n_464),
.B2(n_481),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_474),
.B(n_365),
.C(n_417),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_506),
.B(n_514),
.C(n_515),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_454),
.A2(n_417),
.B1(n_414),
.B2(n_413),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_453),
.A2(n_414),
.B1(n_442),
.B2(n_408),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_461),
.A2(n_404),
.B1(n_408),
.B2(n_411),
.Y(n_509)
);

AOI211xp5_ASAP7_75t_SL g511 ( 
.A1(n_477),
.A2(n_375),
.B(n_360),
.C(n_330),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_448),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_469),
.B(n_330),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_470),
.B(n_315),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_510),
.B(n_457),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_518),
.B(n_531),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_519),
.A2(n_535),
.B1(n_539),
.B2(n_513),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_487),
.B(n_480),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_520),
.B(n_527),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_508),
.Y(n_521)
);

INVx1_ASAP7_75t_SL g552 ( 
.A(n_521),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_490),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_522),
.B(n_542),
.Y(n_548)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_499),
.Y(n_523)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_523),
.Y(n_550)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_512),
.Y(n_525)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_525),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_500),
.B(n_459),
.Y(n_527)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_511),
.Y(n_530)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_530),
.Y(n_556)
);

CKINVDCx16_ASAP7_75t_R g531 ( 
.A(n_505),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_483),
.B(n_462),
.Y(n_532)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_532),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_534),
.A2(n_544),
.B1(n_479),
.B2(n_507),
.Y(n_545)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_514),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_537),
.B(n_541),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_495),
.A2(n_501),
.B1(n_486),
.B2(n_496),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_493),
.B(n_450),
.C(n_466),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_540),
.B(n_506),
.C(n_494),
.Y(n_546)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_515),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_491),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_513),
.A2(n_456),
.B1(n_459),
.B2(n_448),
.Y(n_544)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_545),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_546),
.B(n_562),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_540),
.Y(n_549)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_549),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_529),
.B(n_493),
.C(n_482),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_553),
.B(n_560),
.C(n_566),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_543),
.A2(n_509),
.B1(n_504),
.B2(n_503),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g577 ( 
.A1(n_555),
.A2(n_535),
.B1(n_519),
.B2(n_530),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_516),
.A2(n_455),
.B1(n_513),
.B2(n_473),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_558),
.B(n_559),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_539),
.A2(n_513),
.B1(n_465),
.B2(n_504),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_529),
.B(n_488),
.C(n_492),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_528),
.B(n_489),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_561),
.B(n_563),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_533),
.B(n_484),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_SL g563 ( 
.A(n_520),
.B(n_485),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_564),
.A2(n_521),
.B1(n_513),
.B2(n_502),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_538),
.B(n_527),
.C(n_528),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_538),
.B(n_533),
.C(n_526),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_567),
.B(n_517),
.C(n_524),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_565),
.B(n_522),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_572),
.B(n_573),
.Y(n_590)
);

AO221x1_ASAP7_75t_L g573 ( 
.A1(n_550),
.A2(n_526),
.B1(n_463),
.B2(n_460),
.C(n_543),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_561),
.B(n_517),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_574),
.B(n_582),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_554),
.B(n_544),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_575),
.B(n_586),
.Y(n_588)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_577),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_SL g578 ( 
.A1(n_556),
.A2(n_536),
.B(n_530),
.Y(n_578)
);

OAI21xp5_ASAP7_75t_L g587 ( 
.A1(n_578),
.A2(n_556),
.B(n_564),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_579),
.B(n_567),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_560),
.B(n_546),
.C(n_566),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_581),
.B(n_547),
.C(n_553),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g582 ( 
.A(n_547),
.B(n_534),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_583),
.A2(n_584),
.B1(n_585),
.B2(n_545),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_552),
.A2(n_502),
.B1(n_463),
.B2(n_460),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_552),
.A2(n_375),
.B1(n_370),
.B2(n_344),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_548),
.Y(n_586)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_587),
.Y(n_603)
);

OAI21xp5_ASAP7_75t_L g589 ( 
.A1(n_568),
.A2(n_548),
.B(n_551),
.Y(n_589)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_589),
.A2(n_593),
.B(n_578),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_592),
.B(n_602),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_L g593 ( 
.A1(n_568),
.A2(n_557),
.B(n_555),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g604 ( 
.A(n_594),
.B(n_577),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_596),
.B(n_598),
.Y(n_610)
);

XOR2xp5_ASAP7_75t_L g597 ( 
.A(n_582),
.B(n_562),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_597),
.B(n_583),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_581),
.B(n_563),
.C(n_370),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_576),
.B(n_570),
.C(n_569),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_599),
.B(n_601),
.Y(n_611)
);

INVx6_ASAP7_75t_L g600 ( 
.A(n_576),
.Y(n_600)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_600),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_570),
.B(n_315),
.C(n_316),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g602 ( 
.A(n_579),
.B(n_316),
.Y(n_602)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_604),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_599),
.B(n_600),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_605),
.B(n_609),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_607),
.B(n_591),
.Y(n_616)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_608),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_SL g609 ( 
.A1(n_595),
.A2(n_580),
.B1(n_575),
.B2(n_584),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_602),
.B(n_580),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_612),
.B(n_615),
.Y(n_624)
);

XOR2xp5_ASAP7_75t_L g613 ( 
.A(n_591),
.B(n_571),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_613),
.B(n_598),
.C(n_597),
.Y(n_625)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_590),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_616),
.B(n_617),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_606),
.B(n_596),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_610),
.B(n_601),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_619),
.B(n_621),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_611),
.B(n_589),
.Y(n_621)
);

A2O1A1Ixp33_ASAP7_75t_SL g622 ( 
.A1(n_608),
.A2(n_587),
.B(n_595),
.C(n_588),
.Y(n_622)
);

AOI21x1_ASAP7_75t_L g626 ( 
.A1(n_622),
.A2(n_588),
.B(n_593),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_625),
.B(n_607),
.Y(n_629)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_626),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_629),
.A2(n_630),
.B(n_631),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_623),
.A2(n_603),
.B(n_614),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_624),
.B(n_604),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_SL g632 ( 
.A1(n_628),
.A2(n_618),
.B(n_620),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_SL g636 ( 
.A1(n_632),
.A2(n_634),
.B(n_622),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_SL g634 ( 
.A1(n_627),
.A2(n_622),
.B(n_613),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_636),
.A2(n_637),
.B(n_633),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_635),
.B(n_609),
.C(n_612),
.Y(n_637)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_638),
.Y(n_639)
);

OAI321xp33_ASAP7_75t_L g640 ( 
.A1(n_639),
.A2(n_585),
.A3(n_571),
.B1(n_574),
.B2(n_350),
.C(n_347),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_640),
.A2(n_350),
.B1(n_357),
.B2(n_346),
.Y(n_641)
);


endmodule