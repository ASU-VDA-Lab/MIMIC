module fake_jpeg_18357_n_90 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_90);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_90;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx4f_ASAP7_75t_SL g38 ( 
.A(n_10),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_20),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_48),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_49),
.A2(n_38),
.B1(n_41),
.B2(n_13),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_51),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_47),
.A2(n_39),
.B(n_36),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_4),
.B(n_5),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_50),
.A2(n_37),
.B1(n_40),
.B2(n_43),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_5),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_42),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_61),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_39),
.B1(n_17),
.B2(n_18),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_54),
.B(n_1),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_53),
.B(n_2),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_64),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_60),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_52),
.B(n_3),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_67),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_68),
.A2(n_70),
.B(n_7),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_59),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_6),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_73),
.B(n_19),
.Y(n_80)
);

NOR4xp25_ASAP7_75t_SL g73 ( 
.A(n_67),
.B(n_8),
.C(n_9),
.D(n_11),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_74),
.A2(n_69),
.B1(n_23),
.B2(n_24),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_65),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_81),
.C(n_76),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_80),
.A2(n_78),
.B(n_25),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_83),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_21),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_29),
.C(n_32),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_77),
.Y(n_90)
);


endmodule