module fake_ibex_952_n_1260 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_116, n_61, n_201, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_166, n_195, n_163, n_26, n_188, n_200, n_114, n_199, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_202, n_158, n_132, n_174, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_207, n_54, n_19, n_1260);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_116;
input n_61;
input n_201;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_166;
input n_195;
input n_163;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_207;
input n_54;
input n_19;

output n_1260;

wire n_1084;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_273;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1134;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_280;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_875;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_242;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_279;
wire n_374;
wire n_235;
wire n_538;
wire n_1155;
wire n_459;
wire n_518;
wire n_852;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_715;
wire n_530;
wire n_1214;
wire n_420;
wire n_769;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_230;
wire n_917;
wire n_968;
wire n_1253;
wire n_352;
wire n_558;
wire n_666;
wire n_219;
wire n_1071;
wire n_793;
wire n_937;
wire n_234;
wire n_973;
wire n_1038;
wire n_618;
wire n_662;
wire n_979;
wire n_209;
wire n_1215;
wire n_629;
wire n_573;
wire n_359;
wire n_262;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_369;
wire n_257;
wire n_869;
wire n_718;
wire n_553;
wire n_554;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_564;
wire n_562;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_397;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_499;
wire n_702;
wire n_971;
wire n_451;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_744;
wire n_314;
wire n_563;
wire n_881;
wire n_734;
wire n_1073;
wire n_1108;
wire n_382;
wire n_1239;
wire n_1209;
wire n_288;
wire n_379;
wire n_551;
wire n_729;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_695;
wire n_639;
wire n_482;
wire n_282;
wire n_870;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_462;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_252;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_241;
wire n_231;
wire n_657;
wire n_1156;
wire n_749;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1031;
wire n_372;
wire n_256;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1015;
wire n_663;
wire n_1152;
wire n_371;
wire n_1036;
wire n_974;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_258;
wire n_1129;
wire n_1244;
wire n_449;
wire n_421;
wire n_738;
wire n_1217;
wire n_236;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_840;
wire n_1203;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_944;
wire n_623;
wire n_585;
wire n_483;
wire n_1137;
wire n_222;
wire n_660;
wire n_524;
wire n_1200;
wire n_295;
wire n_1120;
wire n_576;
wire n_388;
wire n_290;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1028;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_267;
wire n_1009;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_413;
wire n_1069;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_998;
wire n_1115;
wire n_801;
wire n_1046;
wire n_882;
wire n_942;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_444;
wire n_986;
wire n_495;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_227;
wire n_1087;
wire n_757;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_517;
wire n_211;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_272;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_863;
wire n_597;
wire n_285;
wire n_1128;
wire n_291;
wire n_318;
wire n_268;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_997;
wire n_891;
wire n_303;
wire n_717;
wire n_668;
wire n_871;
wire n_266;
wire n_485;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_460;
wire n_461;
wire n_903;
wire n_1095;
wire n_1048;
wire n_774;
wire n_588;
wire n_1251;
wire n_1247;
wire n_528;
wire n_260;
wire n_836;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1163;
wire n_677;
wire n_213;
wire n_964;
wire n_916;
wire n_503;
wire n_292;
wire n_895;
wire n_687;
wire n_1035;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_281;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_529;
wire n_626;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_920;
wire n_664;
wire n_1067;
wire n_255;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_578;
wire n_432;
wire n_403;
wire n_423;
wire n_357;
wire n_226;
wire n_216;
wire n_996;
wire n_915;
wire n_1174;
wire n_542;
wire n_900;
wire n_377;
wire n_647;
wire n_317;
wire n_326;
wire n_270;
wire n_259;
wire n_339;
wire n_276;
wire n_348;
wire n_220;
wire n_674;
wire n_287;
wire n_552;
wire n_251;
wire n_1112;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_224;
wire n_508;
wire n_453;
wire n_400;
wire n_1055;
wire n_673;
wire n_798;
wire n_278;
wire n_404;
wire n_1177;
wire n_1025;
wire n_296;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_289;
wire n_716;
wire n_923;
wire n_642;
wire n_286;
wire n_933;
wire n_1037;
wire n_464;
wire n_838;
wire n_1021;
wire n_746;
wire n_1188;
wire n_261;
wire n_742;
wire n_1191;
wire n_221;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_490;
wire n_407;
wire n_595;
wire n_1001;
wire n_269;
wire n_570;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_246;
wire n_922;
wire n_851;
wire n_993;
wire n_253;
wire n_208;
wire n_300;
wire n_1135;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_1066;
wire n_1169;
wire n_245;
wire n_571;
wire n_229;
wire n_648;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_768;
wire n_839;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_976;
wire n_1063;
wire n_834;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_804;
wire n_484;
wire n_480;
wire n_354;
wire n_1057;
wire n_516;
wire n_329;
wire n_1149;
wire n_1176;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_248;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_218;
wire n_277;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_247;
wire n_237;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_782;
wire n_616;
wire n_833;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1221;
wire n_284;
wire n_1047;
wire n_792;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_302;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_298;
wire n_1256;
wire n_587;
wire n_764;
wire n_1206;
wire n_855;
wire n_812;
wire n_232;
wire n_1050;
wire n_599;
wire n_1060;
wire n_756;
wire n_1257;
wire n_274;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1097;
wire n_293;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_249;
wire n_478;
wire n_239;
wire n_336;
wire n_861;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_828;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1098;
wire n_584;
wire n_1187;
wire n_698;
wire n_1061;
wire n_682;
wire n_327;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_265;
wire n_1029;
wire n_470;
wire n_770;
wire n_210;
wire n_941;
wire n_1245;
wire n_243;
wire n_228;
wire n_632;
wire n_373;
wire n_854;
wire n_244;
wire n_343;
wire n_714;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_928;
wire n_898;
wire n_333;
wire n_967;
wire n_736;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_215;
wire n_987;
wire n_750;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1023;
wire n_568;
wire n_813;
wire n_1211;
wire n_1116;
wire n_791;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1074;
wire n_759;
wire n_953;
wire n_1180;
wire n_536;
wire n_1220;
wire n_467;
wire n_427;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_335;
wire n_263;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_735;
wire n_305;
wire n_566;
wire n_416;
wire n_581;
wire n_1089;
wire n_392;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_658;
wire n_1216;
wire n_1026;
wire n_283;
wire n_366;
wire n_1033;
wire n_627;
wire n_990;
wire n_322;
wire n_888;
wire n_582;
wire n_653;
wire n_1205;
wire n_238;
wire n_214;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_225;
wire n_511;
wire n_223;
wire n_381;
wire n_1002;
wire n_1111;
wire n_405;
wire n_612;
wire n_955;
wire n_440;
wire n_342;
wire n_233;
wire n_414;
wire n_378;
wire n_952;
wire n_264;
wire n_1145;
wire n_217;
wire n_537;
wire n_1113;
wire n_913;
wire n_509;
wire n_1164;
wire n_1016;
wire n_240;
wire n_680;
wire n_809;
wire n_856;
wire n_779;
wire n_294;
wire n_493;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_212;
wire n_860;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_297;
wire n_921;
wire n_489;
wire n_254;
wire n_908;
wire n_565;
wire n_1123;
wire n_271;
wire n_984;
wire n_394;
wire n_364;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

INVx2_ASAP7_75t_L g208 ( 
.A(n_17),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_205),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_127),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_38),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_162),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_192),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_16),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_3),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_90),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_145),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_174),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_170),
.Y(n_220)
);

CKINVDCx11_ASAP7_75t_R g221 ( 
.A(n_106),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_73),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_14),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_0),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_175),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_58),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_87),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_155),
.Y(n_228)
);

BUFx10_ASAP7_75t_L g229 ( 
.A(n_116),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_9),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_8),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_125),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_146),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_104),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_42),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_37),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_95),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_18),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_83),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_147),
.Y(n_240)
);

INVxp67_ASAP7_75t_SL g241 ( 
.A(n_100),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_139),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_158),
.Y(n_243)
);

BUFx2_ASAP7_75t_R g244 ( 
.A(n_194),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_188),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_132),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_20),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_69),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_160),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_75),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_199),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_105),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_76),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_82),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_131),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_37),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_206),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_167),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_161),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_159),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_60),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_14),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_183),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_156),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_151),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_52),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_13),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_111),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_17),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_5),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_71),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_178),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_86),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_102),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_48),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_94),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_198),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_57),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_204),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_68),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_177),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_144),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_7),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_30),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_154),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_186),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_45),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_66),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_72),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_112),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_129),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_130),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_120),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_150),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_138),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_108),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_53),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_107),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_84),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_62),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_143),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_20),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_119),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_190),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_97),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_118),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_176),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_9),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_2),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_34),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_23),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_99),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_171),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_91),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_148),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_121),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_54),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_179),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_25),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_197),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_109),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_61),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_74),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_80),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_113),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_202),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_59),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_L g328 ( 
.A(n_172),
.B(n_189),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_128),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_77),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_191),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_115),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_85),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_19),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_26),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_180),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_26),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_28),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_45),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_10),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_10),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_173),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_149),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_141),
.Y(n_344)
);

INVx2_ASAP7_75t_SL g345 ( 
.A(n_103),
.Y(n_345)
);

INVx2_ASAP7_75t_SL g346 ( 
.A(n_134),
.Y(n_346)
);

BUFx10_ASAP7_75t_L g347 ( 
.A(n_163),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_137),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_187),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_93),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_101),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_153),
.Y(n_352)
);

BUFx10_ASAP7_75t_L g353 ( 
.A(n_181),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_12),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_182),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_152),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_140),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_110),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_92),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_28),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_157),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_164),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_117),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_242),
.Y(n_364)
);

NAND2x1p5_ASAP7_75t_L g365 ( 
.A(n_223),
.B(n_1),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_263),
.B(n_1),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_208),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g368 ( 
.A(n_229),
.Y(n_368)
);

AND2x4_ASAP7_75t_L g369 ( 
.A(n_208),
.B(n_2),
.Y(n_369)
);

AND2x4_ASAP7_75t_L g370 ( 
.A(n_302),
.B(n_3),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_302),
.B(n_4),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_334),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_372)
);

BUFx12f_ASAP7_75t_L g373 ( 
.A(n_221),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_339),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_221),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_297),
.B(n_11),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_345),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_226),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_265),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_265),
.B(n_12),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_224),
.B(n_13),
.Y(n_381)
);

OAI22x1_ASAP7_75t_SL g382 ( 
.A1(n_360),
.A2(n_15),
.B1(n_16),
.B2(n_19),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_215),
.Y(n_383)
);

AOI22x1_ASAP7_75t_SL g384 ( 
.A1(n_360),
.A2(n_15),
.B1(n_21),
.B2(n_22),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_346),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_242),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g387 ( 
.A(n_271),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_210),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_245),
.Y(n_389)
);

INVx5_ASAP7_75t_L g390 ( 
.A(n_245),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_216),
.Y(n_391)
);

AND2x6_ASAP7_75t_L g392 ( 
.A(n_239),
.B(n_207),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_259),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_245),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_230),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_217),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_235),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_271),
.Y(n_398)
);

INVx5_ASAP7_75t_L g399 ( 
.A(n_245),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_220),
.Y(n_400)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_209),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_219),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_266),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_236),
.B(n_24),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_219),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_294),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_289),
.Y(n_407)
);

OA21x2_ASAP7_75t_L g408 ( 
.A1(n_212),
.A2(n_257),
.B(n_253),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_222),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_289),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_289),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_231),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_211),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_289),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_303),
.Y(n_415)
);

INVx6_ASAP7_75t_L g416 ( 
.A(n_277),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_303),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_211),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_303),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_294),
.A2(n_25),
.B1(n_27),
.B2(n_29),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_303),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_351),
.Y(n_422)
);

INVx5_ASAP7_75t_L g423 ( 
.A(n_351),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_211),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_351),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_347),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_238),
.B(n_29),
.Y(n_427)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_213),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_262),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_247),
.B(n_31),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_214),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_431)
);

AND2x6_ASAP7_75t_L g432 ( 
.A(n_239),
.B(n_55),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_347),
.B(n_32),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_353),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_233),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_262),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_267),
.B(n_287),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_256),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_330),
.A2(n_35),
.B1(n_36),
.B2(n_39),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_275),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_269),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_330),
.A2(n_35),
.B1(n_36),
.B2(n_39),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_351),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_275),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_237),
.B(n_40),
.Y(n_445)
);

CKINVDCx11_ASAP7_75t_R g446 ( 
.A(n_308),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_282),
.B(n_40),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_275),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_275),
.Y(n_449)
);

INVx6_ASAP7_75t_L g450 ( 
.A(n_282),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_243),
.Y(n_451)
);

NAND2xp33_ASAP7_75t_L g452 ( 
.A(n_363),
.B(n_56),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_304),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_270),
.Y(n_454)
);

INVx5_ASAP7_75t_L g455 ( 
.A(n_304),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_212),
.B(n_41),
.Y(n_456)
);

BUFx12f_ASAP7_75t_L g457 ( 
.A(n_284),
.Y(n_457)
);

BUFx8_ASAP7_75t_SL g458 ( 
.A(n_350),
.Y(n_458)
);

INVxp33_ASAP7_75t_L g459 ( 
.A(n_253),
.Y(n_459)
);

INVx6_ASAP7_75t_L g460 ( 
.A(n_314),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_257),
.B(n_41),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_279),
.Y(n_462)
);

OAI22x1_ASAP7_75t_SL g463 ( 
.A1(n_244),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_350),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_291),
.B(n_46),
.Y(n_465)
);

INVx5_ASAP7_75t_L g466 ( 
.A(n_291),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_246),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_326),
.Y(n_468)
);

BUFx8_ASAP7_75t_SL g469 ( 
.A(n_309),
.Y(n_469)
);

BUFx8_ASAP7_75t_SL g470 ( 
.A(n_310),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_369),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_458),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_369),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_373),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_375),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_456),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_378),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_370),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_393),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_403),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_469),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_395),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_470),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_371),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_456),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_405),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_406),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_388),
.B(n_326),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_408),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_408),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_462),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_446),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_462),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_374),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_462),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_381),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_457),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_412),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_383),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_468),
.Y(n_500)
);

BUFx10_ASAP7_75t_L g501 ( 
.A(n_416),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_438),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_381),
.Y(n_503)
);

INVx4_ASAP7_75t_L g504 ( 
.A(n_392),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_364),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_401),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_364),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_401),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_428),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_428),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_427),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_459),
.B(n_311),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_441),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_R g514 ( 
.A(n_434),
.B(n_218),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_454),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_427),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_397),
.B(n_319),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_380),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_433),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_434),
.B(n_249),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_379),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_398),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_377),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_426),
.Y(n_524)
);

AOI21x1_ASAP7_75t_L g525 ( 
.A1(n_461),
.A2(n_251),
.B(n_250),
.Y(n_525)
);

AND3x2_ASAP7_75t_L g526 ( 
.A(n_463),
.B(n_241),
.C(n_252),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_463),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_385),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_460),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_R g530 ( 
.A(n_368),
.B(n_225),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_447),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_387),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_460),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_R g534 ( 
.A(n_452),
.B(n_227),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_384),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_382),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_466),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_382),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_466),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_453),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_420),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_466),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_420),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_464),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_464),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_366),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_402),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_431),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_431),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_402),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_439),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_439),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_R g553 ( 
.A(n_392),
.B(n_228),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_442),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_376),
.Y(n_555)
);

BUFx6f_ASAP7_75t_SL g556 ( 
.A(n_388),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_372),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_391),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_372),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_391),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_396),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_450),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_R g563 ( 
.A(n_392),
.B(n_232),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_450),
.Y(n_564)
);

BUFx6f_ASAP7_75t_SL g565 ( 
.A(n_400),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_400),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_409),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_465),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_365),
.Y(n_569)
);

NOR2xp67_ASAP7_75t_L g570 ( 
.A(n_455),
.B(n_261),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_367),
.Y(n_571)
);

INVxp33_ASAP7_75t_SL g572 ( 
.A(n_437),
.Y(n_572)
);

BUFx10_ASAP7_75t_L g573 ( 
.A(n_432),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_435),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_435),
.Y(n_575)
);

INVxp33_ASAP7_75t_L g576 ( 
.A(n_404),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_430),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_451),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_467),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_467),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_445),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_367),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_453),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_455),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_455),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_390),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_432),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_390),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_399),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_399),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_423),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_423),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_423),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_413),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_418),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_444),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_424),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_429),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_436),
.Y(n_599)
);

NAND2xp33_ASAP7_75t_L g600 ( 
.A(n_386),
.B(n_234),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_440),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_444),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_448),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_R g604 ( 
.A(n_448),
.B(n_335),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_449),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_389),
.Y(n_606)
);

NOR3xp33_ASAP7_75t_L g607 ( 
.A(n_547),
.B(n_337),
.C(n_283),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_572),
.B(n_576),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_498),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_576),
.B(n_349),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_568),
.B(n_580),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_494),
.Y(n_612)
);

NOR3xp33_ASAP7_75t_L g613 ( 
.A(n_551),
.B(n_340),
.C(n_338),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_504),
.B(n_240),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_603),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_512),
.B(n_341),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_540),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_558),
.B(n_248),
.Y(n_618)
);

OAI221xp5_ASAP7_75t_L g619 ( 
.A1(n_546),
.A2(n_354),
.B1(n_362),
.B2(n_273),
.C(n_276),
.Y(n_619)
);

INVxp67_ASAP7_75t_L g620 ( 
.A(n_482),
.Y(n_620)
);

NOR3xp33_ASAP7_75t_SL g621 ( 
.A(n_535),
.B(n_527),
.C(n_536),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_506),
.B(n_254),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_508),
.B(n_509),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_540),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_510),
.B(n_255),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_523),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_560),
.B(n_258),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_R g628 ( 
.A(n_474),
.B(n_260),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_540),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_517),
.B(n_264),
.Y(n_630)
);

AND2x6_ASAP7_75t_L g631 ( 
.A(n_489),
.B(n_268),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_566),
.B(n_567),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_528),
.Y(n_633)
);

BUFx5_ASAP7_75t_L g634 ( 
.A(n_573),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_574),
.B(n_272),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_481),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_496),
.B(n_328),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_476),
.Y(n_638)
);

INVxp33_ASAP7_75t_L g639 ( 
.A(n_502),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_575),
.B(n_274),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_578),
.B(n_278),
.Y(n_641)
);

NOR3xp33_ASAP7_75t_L g642 ( 
.A(n_552),
.B(n_286),
.C(n_281),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_501),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_476),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_571),
.Y(n_645)
);

NAND2xp33_ASAP7_75t_L g646 ( 
.A(n_553),
.B(n_280),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_501),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_537),
.Y(n_648)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_518),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_503),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_519),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_581),
.B(n_285),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_503),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_579),
.B(n_288),
.Y(n_654)
);

BUFx10_ASAP7_75t_L g655 ( 
.A(n_556),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_511),
.B(n_292),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_582),
.B(n_293),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_516),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_516),
.Y(n_659)
);

INVxp67_ASAP7_75t_L g660 ( 
.A(n_556),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_531),
.B(n_520),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_485),
.B(n_471),
.Y(n_662)
);

BUFx8_ASAP7_75t_L g663 ( 
.A(n_565),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_555),
.B(n_298),
.Y(n_664)
);

NOR2xp67_ASAP7_75t_L g665 ( 
.A(n_584),
.B(n_539),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_542),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_563),
.B(n_299),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_573),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_532),
.B(n_300),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_565),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_569),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_529),
.B(n_305),
.Y(n_672)
);

AOI221xp5_ASAP7_75t_L g673 ( 
.A1(n_541),
.A2(n_290),
.B1(n_295),
.B2(n_296),
.C(n_301),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_493),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_473),
.B(n_307),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_478),
.B(n_313),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_484),
.B(n_315),
.Y(n_677)
);

NAND2xp33_ASAP7_75t_L g678 ( 
.A(n_587),
.B(n_316),
.Y(n_678)
);

BUFx5_ASAP7_75t_L g679 ( 
.A(n_573),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_533),
.B(n_317),
.Y(n_680)
);

NOR3xp33_ASAP7_75t_L g681 ( 
.A(n_554),
.B(n_545),
.C(n_543),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_534),
.B(n_318),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_514),
.B(n_320),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_488),
.B(n_322),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_490),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_525),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_570),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_594),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_530),
.B(n_324),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_521),
.B(n_331),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_522),
.B(n_333),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_564),
.Y(n_692)
);

NOR2x1p5_ASAP7_75t_L g693 ( 
.A(n_492),
.B(n_342),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_595),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_524),
.B(n_352),
.Y(n_695)
);

CKINVDCx16_ASAP7_75t_R g696 ( 
.A(n_499),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_577),
.B(n_355),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_585),
.B(n_357),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_583),
.B(n_359),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_544),
.A2(n_356),
.B1(n_312),
.B2(n_321),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_597),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_586),
.B(n_361),
.Y(n_702)
);

BUFx8_ASAP7_75t_L g703 ( 
.A(n_472),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_513),
.B(n_306),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_599),
.B(n_323),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_601),
.B(n_325),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_605),
.Y(n_707)
);

BUFx8_ASAP7_75t_L g708 ( 
.A(n_483),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_564),
.B(n_327),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_515),
.B(n_329),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_588),
.B(n_332),
.Y(n_711)
);

OR2x6_ASAP7_75t_L g712 ( 
.A(n_526),
.B(n_336),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_589),
.B(n_343),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_475),
.B(n_344),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_562),
.B(n_348),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_497),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_590),
.B(n_591),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_491),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_598),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_592),
.B(n_358),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_593),
.B(n_443),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_486),
.B(n_394),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_495),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_487),
.B(n_63),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_611),
.A2(n_544),
.B1(n_559),
.B2(n_557),
.Y(n_725)
);

NAND2xp33_ASAP7_75t_SL g726 ( 
.A(n_639),
.B(n_477),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_650),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_653),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_663),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_660),
.B(n_479),
.Y(n_730)
);

INVx5_ASAP7_75t_L g731 ( 
.A(n_655),
.Y(n_731)
);

BUFx2_ASAP7_75t_L g732 ( 
.A(n_609),
.Y(n_732)
);

INVx1_ASAP7_75t_SL g733 ( 
.A(n_615),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_658),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_608),
.B(n_480),
.Y(n_735)
);

OR2x6_ASAP7_75t_L g736 ( 
.A(n_692),
.B(n_550),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_659),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_638),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_632),
.B(n_606),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_644),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_685),
.Y(n_741)
);

NOR2xp67_ASAP7_75t_L g742 ( 
.A(n_686),
.B(n_64),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_663),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_620),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_610),
.B(n_500),
.Y(n_745)
);

BUFx2_ASAP7_75t_L g746 ( 
.A(n_696),
.Y(n_746)
);

BUFx2_ASAP7_75t_L g747 ( 
.A(n_671),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_661),
.B(n_500),
.Y(n_748)
);

NOR2x1p5_ASAP7_75t_L g749 ( 
.A(n_636),
.B(n_538),
.Y(n_749)
);

INVx1_ASAP7_75t_SL g750 ( 
.A(n_631),
.Y(n_750)
);

INVx1_ASAP7_75t_SL g751 ( 
.A(n_631),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_642),
.A2(n_548),
.B1(n_549),
.B2(n_600),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_645),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_648),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_613),
.A2(n_619),
.B1(n_673),
.B2(n_681),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_630),
.B(n_596),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_662),
.B(n_47),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_612),
.Y(n_758)
);

CKINVDCx11_ASAP7_75t_R g759 ( 
.A(n_716),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_666),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_700),
.B(n_48),
.Y(n_761)
);

INVx5_ASAP7_75t_L g762 ( 
.A(n_631),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_626),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_657),
.B(n_596),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_631),
.A2(n_604),
.B1(n_407),
.B2(n_410),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_633),
.Y(n_766)
);

BUFx2_ASAP7_75t_L g767 ( 
.A(n_649),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_719),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_651),
.B(n_49),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_618),
.B(n_602),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_670),
.B(n_616),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_664),
.B(n_50),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_703),
.Y(n_773)
);

HB1xp67_ASAP7_75t_L g774 ( 
.A(n_643),
.Y(n_774)
);

OR2x2_ASAP7_75t_SL g775 ( 
.A(n_703),
.B(n_50),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_708),
.Y(n_776)
);

HB1xp67_ASAP7_75t_L g777 ( 
.A(n_647),
.Y(n_777)
);

OR2x6_ASAP7_75t_L g778 ( 
.A(n_712),
.B(n_407),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_637),
.A2(n_410),
.B1(n_425),
.B2(n_411),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_668),
.Y(n_780)
);

BUFx10_ASAP7_75t_L g781 ( 
.A(n_693),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_708),
.Y(n_782)
);

INVx5_ASAP7_75t_L g783 ( 
.A(n_712),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_627),
.B(n_51),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_707),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_607),
.A2(n_414),
.B1(n_425),
.B2(n_415),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_715),
.Y(n_787)
);

INVx5_ASAP7_75t_L g788 ( 
.A(n_718),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_675),
.A2(n_414),
.B1(n_425),
.B2(n_415),
.Y(n_789)
);

INVx5_ASAP7_75t_L g790 ( 
.A(n_718),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_635),
.B(n_640),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_SL g792 ( 
.A1(n_704),
.A2(n_415),
.B1(n_417),
.B2(n_419),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_656),
.A2(n_417),
.B1(n_419),
.B2(n_421),
.Y(n_793)
);

NOR2x2_ASAP7_75t_L g794 ( 
.A(n_628),
.B(n_505),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_665),
.Y(n_795)
);

NOR2x2_ASAP7_75t_L g796 ( 
.A(n_621),
.B(n_507),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_665),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_721),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_668),
.Y(n_799)
);

NOR2x1p5_ASAP7_75t_L g800 ( 
.A(n_698),
.B(n_602),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_710),
.B(n_417),
.Y(n_801)
);

INVxp67_ASAP7_75t_SL g802 ( 
.A(n_709),
.Y(n_802)
);

BUFx12f_ASAP7_75t_L g803 ( 
.A(n_718),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_652),
.B(n_65),
.Y(n_804)
);

INVxp67_ASAP7_75t_L g805 ( 
.A(n_641),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_676),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_688),
.B(n_67),
.Y(n_807)
);

INVx5_ASAP7_75t_L g808 ( 
.A(n_668),
.Y(n_808)
);

INVx2_ASAP7_75t_SL g809 ( 
.A(n_722),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_669),
.B(n_422),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_677),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_623),
.B(n_70),
.Y(n_812)
);

BUFx4f_ASAP7_75t_L g813 ( 
.A(n_694),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_687),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_705),
.Y(n_815)
);

BUFx8_ASAP7_75t_L g816 ( 
.A(n_701),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_706),
.B(n_78),
.Y(n_817)
);

INVx3_ASAP7_75t_L g818 ( 
.A(n_617),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_711),
.Y(n_819)
);

NOR2x1p5_ASAP7_75t_L g820 ( 
.A(n_690),
.B(n_79),
.Y(n_820)
);

OAI21xp33_ASAP7_75t_L g821 ( 
.A1(n_684),
.A2(n_713),
.B(n_720),
.Y(n_821)
);

AND2x6_ASAP7_75t_SL g822 ( 
.A(n_724),
.B(n_81),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_717),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_699),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_654),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_714),
.B(n_88),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_731),
.B(n_702),
.Y(n_827)
);

INVxp67_ASAP7_75t_L g828 ( 
.A(n_767),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_744),
.B(n_691),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_802),
.A2(n_683),
.B1(n_689),
.B2(n_695),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_815),
.B(n_622),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_785),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_819),
.B(n_625),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_753),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_805),
.B(n_747),
.Y(n_835)
);

O2A1O1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_761),
.A2(n_667),
.B(n_646),
.C(n_682),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_803),
.Y(n_837)
);

OAI21xp33_ASAP7_75t_L g838 ( 
.A1(n_821),
.A2(n_680),
.B(n_672),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_791),
.A2(n_614),
.B(n_678),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_755),
.B(n_624),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_725),
.B(n_629),
.Y(n_841)
);

AND2x2_ASAP7_75t_SL g842 ( 
.A(n_807),
.B(n_634),
.Y(n_842)
);

BUFx2_ASAP7_75t_L g843 ( 
.A(n_732),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_806),
.B(n_723),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_R g845 ( 
.A(n_726),
.B(n_679),
.Y(n_845)
);

OR2x2_ASAP7_75t_L g846 ( 
.A(n_725),
.B(n_674),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_758),
.B(n_763),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_787),
.B(n_679),
.Y(n_848)
);

OAI21xp5_ASAP7_75t_L g849 ( 
.A1(n_742),
.A2(n_89),
.B(n_96),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_771),
.B(n_98),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_766),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_768),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_750),
.A2(n_114),
.B1(n_122),
.B2(n_123),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_761),
.B(n_124),
.Y(n_854)
);

AO21x1_ASAP7_75t_L g855 ( 
.A1(n_817),
.A2(n_126),
.B(n_133),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_751),
.A2(n_135),
.B1(n_136),
.B2(n_142),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_L g857 ( 
.A1(n_751),
.A2(n_165),
.B1(n_166),
.B2(n_168),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_R g858 ( 
.A(n_759),
.B(n_169),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_757),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_807),
.B(n_185),
.Y(n_860)
);

BUFx2_ASAP7_75t_L g861 ( 
.A(n_736),
.Y(n_861)
);

BUFx2_ASAP7_75t_L g862 ( 
.A(n_736),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_754),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_741),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_825),
.B(n_193),
.Y(n_865)
);

OAI321xp33_ASAP7_75t_L g866 ( 
.A1(n_786),
.A2(n_195),
.A3(n_196),
.B1(n_200),
.B2(n_201),
.C(n_203),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_760),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_748),
.Y(n_868)
);

O2A1O1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_772),
.A2(n_784),
.B(n_769),
.C(n_756),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_783),
.B(n_731),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_727),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_771),
.B(n_824),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_823),
.B(n_728),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_745),
.A2(n_770),
.B(n_764),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_734),
.B(n_737),
.Y(n_875)
);

BUFx2_ASAP7_75t_SL g876 ( 
.A(n_729),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_800),
.B(n_774),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_738),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_740),
.Y(n_879)
);

A2O1A1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_804),
.A2(n_826),
.B(n_795),
.C(n_797),
.Y(n_880)
);

OAI221xp5_ASAP7_75t_L g881 ( 
.A1(n_752),
.A2(n_736),
.B1(n_813),
.B2(n_733),
.C(n_746),
.Y(n_881)
);

AND2x4_ASAP7_75t_L g882 ( 
.A(n_777),
.B(n_808),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_780),
.Y(n_883)
);

BUFx8_ASAP7_75t_SL g884 ( 
.A(n_773),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_801),
.Y(n_885)
);

A2O1A1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_812),
.A2(n_820),
.B(n_810),
.C(n_814),
.Y(n_886)
);

BUFx2_ASAP7_75t_L g887 ( 
.A(n_743),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_SL g888 ( 
.A1(n_775),
.A2(n_776),
.B1(n_782),
.B2(n_730),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_813),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_809),
.B(n_739),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_765),
.A2(n_818),
.B(n_798),
.C(n_792),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_R g892 ( 
.A(n_781),
.B(n_816),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_816),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_799),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_730),
.B(n_781),
.Y(n_895)
);

O2A1O1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_778),
.A2(n_779),
.B(n_749),
.C(n_793),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_778),
.B(n_762),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_788),
.A2(n_790),
.B(n_789),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_822),
.Y(n_899)
);

A2O1A1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_822),
.A2(n_821),
.B(n_815),
.C(n_806),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_796),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_794),
.A2(n_504),
.B(n_791),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_803),
.Y(n_903)
);

INVx8_ASAP7_75t_L g904 ( 
.A(n_731),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_815),
.B(n_572),
.Y(n_905)
);

INVxp67_ASAP7_75t_L g906 ( 
.A(n_767),
.Y(n_906)
);

O2A1O1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_761),
.A2(n_619),
.B(n_815),
.C(n_632),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_767),
.A2(n_608),
.B1(n_544),
.B2(n_577),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_787),
.A2(n_544),
.B1(n_543),
.B2(n_541),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_744),
.B(n_608),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_744),
.B(n_639),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_785),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_815),
.B(n_572),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_815),
.B(n_572),
.Y(n_914)
);

O2A1O1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_761),
.A2(n_619),
.B(n_815),
.C(n_632),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_815),
.B(n_572),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_802),
.A2(n_815),
.B1(n_558),
.B2(n_561),
.Y(n_917)
);

OR2x2_ASAP7_75t_SL g918 ( 
.A(n_759),
.B(n_696),
.Y(n_918)
);

CKINVDCx20_ASAP7_75t_R g919 ( 
.A(n_759),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_803),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_815),
.B(n_572),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_802),
.A2(n_815),
.B1(n_558),
.B2(n_561),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_815),
.B(n_572),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_802),
.A2(n_815),
.B1(n_558),
.B2(n_561),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_741),
.Y(n_925)
);

CKINVDCx8_ASAP7_75t_R g926 ( 
.A(n_731),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_744),
.Y(n_927)
);

AOI21xp33_ASAP7_75t_L g928 ( 
.A1(n_735),
.A2(n_632),
.B(n_697),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_815),
.B(n_572),
.Y(n_929)
);

O2A1O1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_761),
.A2(n_619),
.B(n_815),
.C(n_632),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_729),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_731),
.B(n_783),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_R g933 ( 
.A(n_726),
.B(n_609),
.Y(n_933)
);

A2O1A1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_821),
.A2(n_815),
.B(n_806),
.C(n_811),
.Y(n_934)
);

INVx4_ASAP7_75t_L g935 ( 
.A(n_731),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_842),
.Y(n_936)
);

BUFx12f_ASAP7_75t_L g937 ( 
.A(n_918),
.Y(n_937)
);

NAND2x1p5_ASAP7_75t_L g938 ( 
.A(n_932),
.B(n_935),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_832),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_912),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_904),
.Y(n_941)
);

OAI21x1_ASAP7_75t_SL g942 ( 
.A1(n_849),
.A2(n_860),
.B(n_902),
.Y(n_942)
);

AO21x2_ASAP7_75t_L g943 ( 
.A1(n_891),
.A2(n_880),
.B(n_900),
.Y(n_943)
);

BUFx3_ASAP7_75t_L g944 ( 
.A(n_904),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_926),
.Y(n_945)
);

BUFx2_ASAP7_75t_SL g946 ( 
.A(n_893),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_934),
.B(n_868),
.Y(n_947)
);

INVx2_ASAP7_75t_SL g948 ( 
.A(n_932),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_851),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_882),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_892),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_882),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_852),
.B(n_847),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_837),
.Y(n_954)
);

INVx2_ASAP7_75t_SL g955 ( 
.A(n_837),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_878),
.Y(n_956)
);

OAI21xp5_ASAP7_75t_L g957 ( 
.A1(n_907),
.A2(n_930),
.B(n_915),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_905),
.B(n_913),
.Y(n_958)
);

NAND2x1p5_ASAP7_75t_L g959 ( 
.A(n_935),
.B(n_897),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_871),
.Y(n_960)
);

INVx1_ASAP7_75t_SL g961 ( 
.A(n_927),
.Y(n_961)
);

BUFx2_ASAP7_75t_R g962 ( 
.A(n_884),
.Y(n_962)
);

AO21x2_ASAP7_75t_L g963 ( 
.A1(n_855),
.A2(n_886),
.B(n_854),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_897),
.B(n_889),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_859),
.B(n_875),
.Y(n_965)
);

INVx5_ASAP7_75t_SL g966 ( 
.A(n_883),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_879),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_840),
.A2(n_839),
.B(n_885),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_914),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_869),
.A2(n_838),
.B(n_874),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_933),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_834),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_916),
.B(n_921),
.Y(n_973)
);

INVx1_ASAP7_75t_SL g974 ( 
.A(n_903),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_841),
.A2(n_901),
.B1(n_861),
.B2(n_862),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_830),
.A2(n_836),
.B(n_873),
.Y(n_976)
);

CKINVDCx11_ASAP7_75t_R g977 ( 
.A(n_919),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_863),
.B(n_867),
.Y(n_978)
);

AO21x1_ASAP7_75t_L g979 ( 
.A1(n_853),
.A2(n_857),
.B(n_856),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_844),
.A2(n_865),
.B(n_833),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_923),
.B(n_929),
.Y(n_981)
);

INVxp33_ASAP7_75t_L g982 ( 
.A(n_911),
.Y(n_982)
);

INVx6_ASAP7_75t_SL g983 ( 
.A(n_827),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_903),
.Y(n_984)
);

INVx1_ASAP7_75t_SL g985 ( 
.A(n_920),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_920),
.Y(n_986)
);

INVxp33_ASAP7_75t_L g987 ( 
.A(n_835),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_931),
.Y(n_988)
);

INVx2_ASAP7_75t_SL g989 ( 
.A(n_887),
.Y(n_989)
);

BUFx2_ASAP7_75t_SL g990 ( 
.A(n_870),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_876),
.Y(n_991)
);

INVx3_ASAP7_75t_SL g992 ( 
.A(n_877),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_908),
.B(n_909),
.Y(n_993)
);

BUFx12f_ASAP7_75t_L g994 ( 
.A(n_843),
.Y(n_994)
);

OAI21x1_ASAP7_75t_SL g995 ( 
.A1(n_896),
.A2(n_917),
.B(n_924),
.Y(n_995)
);

BUFx4_ASAP7_75t_SL g996 ( 
.A(n_846),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_894),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_827),
.B(n_877),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_831),
.B(n_922),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_864),
.Y(n_1000)
);

AOI22x1_ASAP7_75t_L g1001 ( 
.A1(n_925),
.A2(n_895),
.B1(n_866),
.B2(n_828),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_906),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_872),
.Y(n_1003)
);

OR2x6_ASAP7_75t_L g1004 ( 
.A(n_888),
.B(n_910),
.Y(n_1004)
);

CKINVDCx16_ASAP7_75t_R g1005 ( 
.A(n_858),
.Y(n_1005)
);

AO21x2_ASAP7_75t_L g1006 ( 
.A1(n_845),
.A2(n_928),
.B(n_850),
.Y(n_1006)
);

INVx4_ASAP7_75t_L g1007 ( 
.A(n_881),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_SL g1008 ( 
.A1(n_890),
.A2(n_848),
.B(n_829),
.Y(n_1008)
);

BUFx3_ASAP7_75t_L g1009 ( 
.A(n_904),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_934),
.B(n_868),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_832),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_934),
.A2(n_915),
.B(n_907),
.Y(n_1012)
);

INVx1_ASAP7_75t_SL g1013 ( 
.A(n_927),
.Y(n_1013)
);

AOI22x1_ASAP7_75t_L g1014 ( 
.A1(n_899),
.A2(n_820),
.B1(n_902),
.B2(n_898),
.Y(n_1014)
);

AOI22x1_ASAP7_75t_L g1015 ( 
.A1(n_899),
.A2(n_820),
.B1(n_902),
.B2(n_898),
.Y(n_1015)
);

NAND2x1p5_ASAP7_75t_L g1016 ( 
.A(n_842),
.B(n_932),
.Y(n_1016)
);

OR2x6_ASAP7_75t_L g1017 ( 
.A(n_904),
.B(n_876),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_927),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_832),
.Y(n_1019)
);

BUFx3_ASAP7_75t_L g1020 ( 
.A(n_904),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_926),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_904),
.Y(n_1022)
);

AND2x2_ASAP7_75t_SL g1023 ( 
.A(n_842),
.B(n_897),
.Y(n_1023)
);

OR2x2_ASAP7_75t_L g1024 ( 
.A(n_905),
.B(n_913),
.Y(n_1024)
);

INVx5_ASAP7_75t_L g1025 ( 
.A(n_904),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_904),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_926),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_904),
.Y(n_1028)
);

NAND2x1p5_ASAP7_75t_L g1029 ( 
.A(n_1023),
.B(n_1025),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_947),
.Y(n_1030)
);

INVx1_ASAP7_75t_SL g1031 ( 
.A(n_941),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_969),
.B(n_958),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_1018),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_966),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_961),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_947),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1010),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_981),
.B(n_973),
.Y(n_1038)
);

INVxp67_ASAP7_75t_L g1039 ( 
.A(n_1002),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_956),
.B(n_967),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_960),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_1023),
.A2(n_936),
.B1(n_999),
.B2(n_965),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_1025),
.Y(n_1043)
);

OAI22xp33_ASAP7_75t_L g1044 ( 
.A1(n_1005),
.A2(n_987),
.B1(n_999),
.B2(n_1004),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_978),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_995),
.A2(n_993),
.B1(n_1007),
.B2(n_937),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_978),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_L g1048 ( 
.A1(n_1007),
.A2(n_987),
.B1(n_975),
.B2(n_982),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_968),
.Y(n_1049)
);

CKINVDCx6p67_ASAP7_75t_R g1050 ( 
.A(n_1025),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_975),
.A2(n_982),
.B1(n_1004),
.B2(n_981),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_1025),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_1024),
.B(n_965),
.Y(n_1053)
);

OA21x2_ASAP7_75t_L g1054 ( 
.A1(n_970),
.A2(n_1012),
.B(n_957),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_957),
.B(n_936),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_968),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_1013),
.Y(n_1057)
);

CKINVDCx11_ASAP7_75t_R g1058 ( 
.A(n_977),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_949),
.B(n_953),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_939),
.Y(n_1060)
);

AOI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_1004),
.A2(n_1003),
.B1(n_953),
.B2(n_971),
.Y(n_1061)
);

HB1xp67_ASAP7_75t_L g1062 ( 
.A(n_1017),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_1008),
.A2(n_976),
.B1(n_994),
.B2(n_980),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_972),
.B(n_940),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1011),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1019),
.Y(n_1066)
);

INVx1_ASAP7_75t_SL g1067 ( 
.A(n_941),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1012),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_966),
.Y(n_1069)
);

AOI22xp33_ASAP7_75t_SL g1070 ( 
.A1(n_1001),
.A2(n_1016),
.B1(n_996),
.B2(n_990),
.Y(n_1070)
);

CKINVDCx6p67_ASAP7_75t_R g1071 ( 
.A(n_1017),
.Y(n_1071)
);

BUFx10_ASAP7_75t_L g1072 ( 
.A(n_1017),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_944),
.Y(n_1073)
);

INVx1_ASAP7_75t_SL g1074 ( 
.A(n_944),
.Y(n_1074)
);

CKINVDCx6p67_ASAP7_75t_R g1075 ( 
.A(n_1009),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_943),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_996),
.Y(n_1077)
);

AO21x2_ASAP7_75t_L g1078 ( 
.A1(n_942),
.A2(n_943),
.B(n_963),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_966),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_1055),
.B(n_1006),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1059),
.B(n_950),
.Y(n_1081)
);

BUFx2_ASAP7_75t_L g1082 ( 
.A(n_1029),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_1035),
.Y(n_1083)
);

NAND3xp33_ASAP7_75t_SL g1084 ( 
.A(n_1070),
.B(n_991),
.C(n_951),
.Y(n_1084)
);

NAND2xp33_ASAP7_75t_R g1085 ( 
.A(n_1071),
.B(n_1027),
.Y(n_1085)
);

OR2x6_ASAP7_75t_L g1086 ( 
.A(n_1029),
.B(n_938),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_1068),
.B(n_1006),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1054),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1030),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_1029),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1059),
.B(n_950),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1030),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_R g1093 ( 
.A(n_1050),
.B(n_977),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_SL g1094 ( 
.A1(n_1042),
.A2(n_1077),
.B1(n_1072),
.B2(n_1062),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1055),
.B(n_952),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1041),
.B(n_1040),
.Y(n_1096)
);

HB1xp67_ASAP7_75t_L g1097 ( 
.A(n_1057),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_1038),
.B(n_1032),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1041),
.B(n_997),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1036),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1040),
.B(n_1000),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_1075),
.Y(n_1102)
);

CKINVDCx16_ASAP7_75t_R g1103 ( 
.A(n_1073),
.Y(n_1103)
);

INVxp67_ASAP7_75t_L g1104 ( 
.A(n_1033),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_R g1105 ( 
.A(n_1050),
.B(n_1028),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1036),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1051),
.A2(n_998),
.B1(n_979),
.B2(n_989),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_1075),
.Y(n_1108)
);

NAND3xp33_ASAP7_75t_L g1109 ( 
.A(n_1063),
.B(n_1015),
.C(n_1014),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1037),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_1072),
.Y(n_1111)
);

BUFx3_ASAP7_75t_L g1112 ( 
.A(n_1073),
.Y(n_1112)
);

HB1xp67_ASAP7_75t_L g1113 ( 
.A(n_1064),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1037),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_R g1115 ( 
.A(n_1071),
.B(n_1028),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_R g1116 ( 
.A(n_1058),
.B(n_1026),
.Y(n_1116)
);

OR2x2_ASAP7_75t_L g1117 ( 
.A(n_1053),
.B(n_992),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_1072),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1087),
.B(n_1076),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1087),
.B(n_1096),
.Y(n_1120)
);

NOR2x1p5_ASAP7_75t_L g1121 ( 
.A(n_1090),
.B(n_1043),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1089),
.Y(n_1122)
);

INVx1_ASAP7_75t_SL g1123 ( 
.A(n_1112),
.Y(n_1123)
);

HB1xp67_ASAP7_75t_L g1124 ( 
.A(n_1113),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1089),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1096),
.B(n_1049),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1098),
.B(n_1060),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_1092),
.B(n_1049),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_1092),
.B(n_1056),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1100),
.B(n_1056),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1083),
.B(n_1060),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_1097),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_1112),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1104),
.B(n_1066),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1103),
.B(n_1066),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1106),
.B(n_1078),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_1082),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1101),
.B(n_1099),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1122),
.Y(n_1139)
);

HB1xp67_ASAP7_75t_L g1140 ( 
.A(n_1124),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1120),
.B(n_1080),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1120),
.B(n_1080),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1126),
.B(n_1110),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1126),
.B(n_1110),
.Y(n_1144)
);

INVx2_ASAP7_75t_SL g1145 ( 
.A(n_1133),
.Y(n_1145)
);

NAND2x1_ASAP7_75t_L g1146 ( 
.A(n_1137),
.B(n_1082),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1119),
.B(n_1080),
.Y(n_1147)
);

CKINVDCx20_ASAP7_75t_R g1148 ( 
.A(n_1135),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1132),
.B(n_1114),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1119),
.B(n_1088),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1136),
.B(n_1088),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_1123),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1122),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1125),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1139),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1141),
.B(n_1136),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1141),
.B(n_1138),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1142),
.B(n_1128),
.Y(n_1158)
);

NOR2x1_ASAP7_75t_L g1159 ( 
.A(n_1146),
.B(n_1121),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_1152),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1139),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1142),
.B(n_1128),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1148),
.B(n_1102),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1147),
.B(n_1129),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1153),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1147),
.B(n_1129),
.Y(n_1166)
);

OR2x2_ASAP7_75t_L g1167 ( 
.A(n_1140),
.B(n_1131),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1150),
.B(n_1130),
.Y(n_1168)
);

INVx1_ASAP7_75t_SL g1169 ( 
.A(n_1145),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1150),
.B(n_1130),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1153),
.Y(n_1171)
);

OR2x2_ASAP7_75t_L g1172 ( 
.A(n_1167),
.B(n_1149),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1155),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1164),
.B(n_1145),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_1159),
.B(n_1151),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1156),
.B(n_1158),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1164),
.B(n_1143),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1156),
.B(n_1151),
.Y(n_1178)
);

OAI322xp33_ASAP7_75t_L g1179 ( 
.A1(n_1167),
.A2(n_1127),
.A3(n_1144),
.B1(n_1134),
.B2(n_1044),
.C1(n_1039),
.C2(n_1154),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1155),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_1169),
.Y(n_1181)
);

INVxp67_ASAP7_75t_SL g1182 ( 
.A(n_1160),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1161),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1166),
.B(n_1154),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1161),
.Y(n_1185)
);

OAI31xp33_ASAP7_75t_L g1186 ( 
.A1(n_1160),
.A2(n_1121),
.A3(n_1123),
.B(n_1137),
.Y(n_1186)
);

OAI32xp33_ASAP7_75t_L g1187 ( 
.A1(n_1163),
.A2(n_1085),
.A3(n_1102),
.B1(n_1108),
.B2(n_1090),
.Y(n_1187)
);

INVx2_ASAP7_75t_SL g1188 ( 
.A(n_1181),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_SL g1189 ( 
.A1(n_1179),
.A2(n_1108),
.B(n_1084),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1182),
.A2(n_1187),
.B(n_1186),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1176),
.B(n_1166),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1173),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1176),
.B(n_1158),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1172),
.A2(n_1046),
.B1(n_1048),
.B2(n_1117),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1187),
.A2(n_1175),
.B(n_1094),
.Y(n_1195)
);

OAI21xp33_ASAP7_75t_L g1196 ( 
.A1(n_1175),
.A2(n_1162),
.B(n_1170),
.Y(n_1196)
);

OAI221xp5_ASAP7_75t_L g1197 ( 
.A1(n_1190),
.A2(n_1172),
.B1(n_1107),
.B2(n_1174),
.C(n_1184),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1188),
.Y(n_1198)
);

O2A1O1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1195),
.A2(n_985),
.B(n_974),
.C(n_1067),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_SL g1200 ( 
.A1(n_1194),
.A2(n_1031),
.B(n_1074),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1192),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1196),
.B(n_1175),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_SL g1203 ( 
.A1(n_1191),
.A2(n_1093),
.B1(n_1115),
.B2(n_1105),
.Y(n_1203)
);

OAI211xp5_ASAP7_75t_L g1204 ( 
.A1(n_1189),
.A2(n_1116),
.B(n_1061),
.C(n_1118),
.Y(n_1204)
);

OR2x2_ASAP7_75t_L g1205 ( 
.A(n_1193),
.B(n_1177),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_1194),
.B(n_1178),
.Y(n_1206)
);

AOI221xp5_ASAP7_75t_L g1207 ( 
.A1(n_1206),
.A2(n_1185),
.B1(n_1180),
.B2(n_1183),
.C(n_1171),
.Y(n_1207)
);

NOR2x1_ASAP7_75t_L g1208 ( 
.A(n_1204),
.B(n_1200),
.Y(n_1208)
);

OR2x2_ASAP7_75t_L g1209 ( 
.A(n_1205),
.B(n_1206),
.Y(n_1209)
);

AOI221xp5_ASAP7_75t_L g1210 ( 
.A1(n_1199),
.A2(n_1165),
.B1(n_1171),
.B2(n_1178),
.C(n_1162),
.Y(n_1210)
);

NOR3xp33_ASAP7_75t_L g1211 ( 
.A(n_1200),
.B(n_1203),
.C(n_1198),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1201),
.Y(n_1212)
);

NOR3xp33_ASAP7_75t_L g1213 ( 
.A(n_1197),
.B(n_1021),
.C(n_1027),
.Y(n_1213)
);

NOR3xp33_ASAP7_75t_SL g1214 ( 
.A(n_1208),
.B(n_962),
.C(n_1118),
.Y(n_1214)
);

NOR2x1_ASAP7_75t_L g1215 ( 
.A(n_1209),
.B(n_946),
.Y(n_1215)
);

OAI21xp33_ASAP7_75t_L g1216 ( 
.A1(n_1211),
.A2(n_1213),
.B(n_1207),
.Y(n_1216)
);

OAI21xp33_ASAP7_75t_L g1217 ( 
.A1(n_1212),
.A2(n_1202),
.B(n_1210),
.Y(n_1217)
);

OR3x1_ASAP7_75t_L g1218 ( 
.A(n_1208),
.B(n_962),
.C(n_1165),
.Y(n_1218)
);

AOI221xp5_ASAP7_75t_L g1219 ( 
.A1(n_1211),
.A2(n_1157),
.B1(n_1170),
.B2(n_1168),
.C(n_955),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1209),
.B(n_1157),
.Y(n_1220)
);

AOI211xp5_ASAP7_75t_L g1221 ( 
.A1(n_1216),
.A2(n_1217),
.B(n_1219),
.C(n_1214),
.Y(n_1221)
);

AOI211xp5_ASAP7_75t_L g1222 ( 
.A1(n_1218),
.A2(n_945),
.B(n_1026),
.C(n_1022),
.Y(n_1222)
);

AOI311xp33_ASAP7_75t_L g1223 ( 
.A1(n_1220),
.A2(n_1215),
.A3(n_1065),
.B(n_1045),
.C(n_1047),
.Y(n_1223)
);

AOI222xp33_ASAP7_75t_L g1224 ( 
.A1(n_1216),
.A2(n_945),
.B1(n_988),
.B2(n_1109),
.C1(n_1021),
.C2(n_984),
.Y(n_1224)
);

AOI211xp5_ASAP7_75t_L g1225 ( 
.A1(n_1216),
.A2(n_1009),
.B(n_1020),
.C(n_1022),
.Y(n_1225)
);

OAI32xp33_ASAP7_75t_L g1226 ( 
.A1(n_1216),
.A2(n_988),
.A3(n_1043),
.B1(n_1052),
.B2(n_1020),
.Y(n_1226)
);

OAI211xp5_ASAP7_75t_L g1227 ( 
.A1(n_1214),
.A2(n_1052),
.B(n_954),
.C(n_986),
.Y(n_1227)
);

AOI221x1_ASAP7_75t_SL g1228 ( 
.A1(n_1216),
.A2(n_998),
.B1(n_964),
.B2(n_1081),
.C(n_1091),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1221),
.B(n_1168),
.Y(n_1229)
);

AOI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1224),
.A2(n_1111),
.B1(n_992),
.B2(n_1086),
.Y(n_1230)
);

NOR2x1p5_ASAP7_75t_L g1231 ( 
.A(n_1226),
.B(n_954),
.Y(n_1231)
);

NOR2x1_ASAP7_75t_L g1232 ( 
.A(n_1227),
.B(n_986),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1225),
.Y(n_1233)
);

NOR2x1_ASAP7_75t_L g1234 ( 
.A(n_1223),
.B(n_1034),
.Y(n_1234)
);

AOI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1222),
.A2(n_1111),
.B1(n_1086),
.B2(n_1117),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1229),
.Y(n_1236)
);

NAND4xp25_ASAP7_75t_L g1237 ( 
.A(n_1233),
.B(n_1228),
.C(n_1234),
.D(n_1232),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1235),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1231),
.B(n_1095),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1238),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1239),
.Y(n_1241)
);

INVx1_ASAP7_75t_SL g1242 ( 
.A(n_1236),
.Y(n_1242)
);

CKINVDCx16_ASAP7_75t_R g1243 ( 
.A(n_1237),
.Y(n_1243)
);

XOR2xp5_ASAP7_75t_L g1244 ( 
.A(n_1243),
.B(n_1230),
.Y(n_1244)
);

XNOR2x2_ASAP7_75t_L g1245 ( 
.A(n_1242),
.B(n_983),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1240),
.B(n_1241),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1246),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1245),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1244),
.Y(n_1249)
);

INVxp67_ASAP7_75t_L g1250 ( 
.A(n_1246),
.Y(n_1250)
);

OAI22x1_ASAP7_75t_L g1251 ( 
.A1(n_1249),
.A2(n_948),
.B1(n_964),
.B2(n_959),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1247),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_1248),
.Y(n_1253)
);

OAI22x1_ASAP7_75t_L g1254 ( 
.A1(n_1250),
.A2(n_959),
.B1(n_1034),
.B2(n_1079),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_1253),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1252),
.Y(n_1256)
);

NAND3xp33_ASAP7_75t_L g1257 ( 
.A(n_1256),
.B(n_1250),
.C(n_1251),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1257),
.A2(n_1255),
.B1(n_1254),
.B2(n_1069),
.Y(n_1258)
);

OR2x6_ASAP7_75t_L g1259 ( 
.A(n_1258),
.B(n_1034),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1259),
.A2(n_983),
.B1(n_1079),
.B2(n_1069),
.Y(n_1260)
);


endmodule