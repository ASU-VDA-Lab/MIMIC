module fake_jpeg_31874_n_119 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_119);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_119;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx16f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx4f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_3),
.B(n_11),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_6),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_32),
.Y(n_44)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_0),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_5),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_11),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

CKINVDCx6p67_ASAP7_75t_R g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_21),
.B1(n_17),
.B2(n_13),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_36),
.B1(n_27),
.B2(n_21),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_10),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_26),
.B(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_30),
.B(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_44),
.B(n_20),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_53),
.B(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_60),
.Y(n_72)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_27),
.B1(n_41),
.B2(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_16),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_16),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_37),
.C(n_25),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_47),
.C(n_45),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_48),
.A2(n_14),
.B1(n_13),
.B2(n_36),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_29),
.B1(n_33),
.B2(n_31),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_40),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_67),
.Y(n_73)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_15),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_69),
.Y(n_78)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_75),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_67),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_58),
.A2(n_14),
.B1(n_47),
.B2(n_49),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_81),
.Y(n_83)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_85),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_53),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_78),
.B(n_61),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_87),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_73),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_64),
.C(n_59),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_89),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_61),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_90),
.A2(n_73),
.B(n_69),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_82),
.A2(n_77),
.B1(n_78),
.B2(n_70),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_91),
.A2(n_74),
.B1(n_55),
.B2(n_70),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_84),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_93),
.B(n_88),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_96),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_99),
.B(n_100),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_72),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_95),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_79),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_102),
.B(n_103),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_35),
.Y(n_110)
);

OAI321xp33_ASAP7_75t_L g108 ( 
.A1(n_101),
.A2(n_91),
.A3(n_97),
.B1(n_96),
.B2(n_8),
.C(n_10),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_108),
.A2(n_0),
.B(n_1),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_99),
.C(n_49),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_110),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_105),
.A2(n_106),
.B(n_8),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_111),
.A2(n_112),
.B(n_1),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_1),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_SL g116 ( 
.A1(n_115),
.A2(n_2),
.B(n_35),
.C(n_56),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_116),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_113),
.B1(n_56),
.B2(n_35),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_14),
.Y(n_119)
);


endmodule