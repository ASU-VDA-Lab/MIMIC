module real_jpeg_23783_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_173;
wire n_40;
wire n_105;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_258;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_0),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_0),
.B(n_34),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_0),
.B(n_46),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_0),
.B(n_48),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_0),
.B(n_53),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_0),
.B(n_63),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_0),
.B(n_28),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_0),
.B(n_17),
.Y(n_208)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_2),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_2),
.B(n_41),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_2),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_2),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_2),
.B(n_63),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_2),
.B(n_28),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_2),
.B(n_53),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_2),
.B(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_3),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_3),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_3),
.B(n_63),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_4),
.B(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_4),
.B(n_53),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_4),
.B(n_48),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_4),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_4),
.B(n_17),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_6),
.B(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_6),
.B(n_63),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_6),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_6),
.B(n_48),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_6),
.B(n_53),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_6),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_6),
.B(n_28),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_8),
.B(n_28),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_8),
.B(n_53),
.Y(n_93)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_10),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_13),
.B(n_53),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_13),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_13),
.B(n_41),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_13),
.B(n_28),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_13),
.B(n_182),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_14),
.B(n_48),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_14),
.B(n_41),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_14),
.B(n_63),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_14),
.B(n_28),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_14),
.B(n_46),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_16),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_16),
.B(n_63),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_16),
.B(n_48),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_16),
.B(n_53),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_16),
.B(n_28),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_16),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_16),
.B(n_41),
.Y(n_236)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_17),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_150),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_127),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_69),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_50),
.C(n_56),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_22),
.B(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.C(n_44),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_23),
.B(n_266),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_24),
.B(n_51),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_24),
.B(n_52),
.C(n_55),
.Y(n_115)
);

FAx1_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_30),
.CI(n_33),
.CON(n_24),
.SN(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_27),
.B(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_32),
.Y(n_218)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_35),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_36),
.A2(n_37),
.B(n_40),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_36),
.B(n_44),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_39),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_47),
.C(n_49),
.Y(n_44)
);

FAx1_ASAP7_75t_SL g131 ( 
.A(n_45),
.B(n_47),
.CI(n_49),
.CON(n_131),
.SN(n_131)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_50),
.B(n_56),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_53),
.Y(n_214)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_65),
.C(n_67),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_57),
.B(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_61),
.C(n_62),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_58),
.B(n_255),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_59),
.B(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_61),
.B(n_62),
.Y(n_255)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_65),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_94),
.B2(n_126),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_85),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_79),
.B1(n_83),
.B2(n_84),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_77),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_78),
.B(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_79),
.A2(n_83),
.B1(n_87),
.B2(n_114),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_87),
.C(n_88),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_87),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_89),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx24_ASAP7_75t_SL g273 ( 
.A(n_90),
.Y(n_273)
);

FAx1_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_92),
.CI(n_93),
.CON(n_90),
.SN(n_90)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

BUFx24_ASAP7_75t_SL g272 ( 
.A(n_94),
.Y(n_272)
);

FAx1_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_115),
.CI(n_116),
.CON(n_94),
.SN(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_105),
.C(n_111),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_96),
.B(n_147),
.Y(n_146)
);

BUFx24_ASAP7_75t_SL g277 ( 
.A(n_96),
.Y(n_277)
);

FAx1_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_100),
.CI(n_103),
.CON(n_96),
.SN(n_96)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_100),
.C(n_103),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_101),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_111),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.C(n_109),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_106),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_125),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_120),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_146),
.C(n_148),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_128),
.A2(n_129),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_142),
.C(n_144),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_130),
.B(n_262),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.C(n_138),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_131),
.B(n_248),
.Y(n_247)
);

BUFx24_ASAP7_75t_SL g274 ( 
.A(n_131),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_132),
.A2(n_133),
.B1(n_138),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_138),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.C(n_141),
.Y(n_138)
);

FAx1_ASAP7_75t_SL g229 ( 
.A(n_139),
.B(n_140),
.CI(n_141),
.CON(n_229),
.SN(n_229)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_142),
.B(n_144),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_146),
.B(n_148),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_268),
.C(n_269),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_258),
.C(n_259),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_241),
.C(n_242),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_223),
.C(n_224),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_185),
.C(n_197),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_169),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_164),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_157),
.B(n_164),
.C(n_169),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.C(n_162),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_158),
.A2(n_159),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_165),
.B(n_167),
.C(n_168),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_176),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_170),
.B(n_177),
.C(n_178),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_174),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_171),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_184),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_179),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_180),
.B(n_184),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.C(n_196),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_189),
.A2(n_190),
.B1(n_196),
.B2(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_201)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_196),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_219),
.C(n_220),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_206),
.C(n_211),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_204),
.C(n_205),
.Y(n_219)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.C(n_215),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_230),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_231),
.C(n_240),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_229),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_228),
.C(n_229),
.Y(n_245)
);

BUFx24_ASAP7_75t_SL g275 ( 
.A(n_229),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_240),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_238),
.B2(n_239),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_234),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_237),
.C(n_239),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_238),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_250),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_246),
.C(n_250),
.Y(n_258)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_254),
.C(n_256),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_256),
.B2(n_257),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_253),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_254),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_263),
.B2(n_267),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_264),
.C(n_265),
.Y(n_268)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_263),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_270),
.Y(n_271)
);


endmodule