module fake_netlist_1_7216_n_1044 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_1044);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1044;
wire n_663;
wire n_707;
wire n_791;
wire n_513;
wire n_361;
wire n_963;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_786;
wire n_724;
wire n_857;
wire n_345;
wire n_360;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_769;
wire n_927;
wire n_596;
wire n_286;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_572;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_975;
wire n_279;
wire n_303;
wire n_968;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_945;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_1011;
wire n_1025;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_624;
wire n_426;
wire n_725;
wire n_844;
wire n_818;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_634;
wire n_307;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_950;
wire n_460;
wire n_478;
wire n_415;
wire n_482;
wire n_703;
wire n_394;
wire n_813;
wire n_442;
wire n_331;
wire n_485;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_729;
wire n_519;
wire n_699;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_880;
wire n_799;
wire n_370;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_899;
wire n_260;
wire n_806;
wire n_881;
wire n_539;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_1029;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_721;
wire n_656;
wire n_438;
wire n_445;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_811;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_924;
wire n_912;
wire n_947;
wire n_1043;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1040;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_695;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_631;
wire n_453;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_992;
wire n_269;
INVx1_ASAP7_75t_L g257 ( .A(n_52), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_117), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_85), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_83), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_223), .Y(n_261) );
INVxp33_ASAP7_75t_L g262 ( .A(n_237), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g263 ( .A(n_241), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_42), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_244), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_218), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_20), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_159), .Y(n_268) );
CKINVDCx16_ASAP7_75t_R g269 ( .A(n_69), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_209), .Y(n_270) );
INVxp67_ASAP7_75t_SL g271 ( .A(n_33), .Y(n_271) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_230), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_28), .Y(n_273) );
CKINVDCx16_ASAP7_75t_R g274 ( .A(n_4), .Y(n_274) );
INVxp33_ASAP7_75t_SL g275 ( .A(n_71), .Y(n_275) );
NOR2xp67_ASAP7_75t_L g276 ( .A(n_169), .B(n_198), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_16), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_228), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_114), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_43), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_131), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_147), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_238), .Y(n_283) );
INVxp33_ASAP7_75t_SL g284 ( .A(n_15), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_252), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_157), .Y(n_286) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_13), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_108), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_135), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_216), .Y(n_290) );
INVxp33_ASAP7_75t_SL g291 ( .A(n_161), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_239), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_181), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_247), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_80), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_109), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_42), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_106), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_188), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_53), .Y(n_300) );
BUFx10_ASAP7_75t_L g301 ( .A(n_45), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_38), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_60), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_225), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_125), .Y(n_305) );
CKINVDCx14_ASAP7_75t_R g306 ( .A(n_178), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_229), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_170), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_212), .Y(n_309) );
INVx1_ASAP7_75t_SL g310 ( .A(n_141), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_165), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_59), .Y(n_312) );
CKINVDCx20_ASAP7_75t_R g313 ( .A(n_145), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_160), .Y(n_314) );
BUFx3_ASAP7_75t_L g315 ( .A(n_91), .Y(n_315) );
INVxp67_ASAP7_75t_SL g316 ( .A(n_72), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_179), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_32), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_27), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_103), .Y(n_320) );
INVxp67_ASAP7_75t_L g321 ( .A(n_62), .Y(n_321) );
INVxp33_ASAP7_75t_SL g322 ( .A(n_227), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_11), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_185), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_45), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_6), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_221), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_88), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_251), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_166), .Y(n_330) );
INVxp67_ASAP7_75t_L g331 ( .A(n_182), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_99), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_94), .Y(n_333) );
INVxp33_ASAP7_75t_SL g334 ( .A(n_87), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_47), .Y(n_335) );
INVxp33_ASAP7_75t_L g336 ( .A(n_245), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_201), .Y(n_337) );
INVxp33_ASAP7_75t_SL g338 ( .A(n_16), .Y(n_338) );
INVxp67_ASAP7_75t_L g339 ( .A(n_43), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_193), .Y(n_340) );
INVxp33_ASAP7_75t_SL g341 ( .A(n_118), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_78), .Y(n_342) );
BUFx3_ASAP7_75t_L g343 ( .A(n_205), .Y(n_343) );
BUFx2_ASAP7_75t_L g344 ( .A(n_208), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_206), .Y(n_345) );
INVxp67_ASAP7_75t_L g346 ( .A(n_248), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_191), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_171), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_250), .Y(n_349) );
INVx1_ASAP7_75t_SL g350 ( .A(n_111), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_90), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_168), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_137), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_58), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_220), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_105), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_33), .Y(n_357) );
CKINVDCx20_ASAP7_75t_R g358 ( .A(n_233), .Y(n_358) );
INVxp33_ASAP7_75t_SL g359 ( .A(n_96), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_207), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_77), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_55), .Y(n_362) );
INVxp67_ASAP7_75t_SL g363 ( .A(n_54), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_175), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_9), .Y(n_365) );
CKINVDCx20_ASAP7_75t_R g366 ( .A(n_124), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_8), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_144), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_232), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_5), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_98), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_107), .Y(n_372) );
INVx3_ASAP7_75t_L g373 ( .A(n_199), .Y(n_373) );
INVxp33_ASAP7_75t_SL g374 ( .A(n_155), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_64), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_311), .B(n_0), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_311), .B(n_0), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_344), .B(n_1), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_370), .B(n_1), .Y(n_379) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_324), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_373), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_258), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_258), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_344), .B(n_2), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_370), .B(n_2), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_265), .Y(n_386) );
BUFx2_ASAP7_75t_L g387 ( .A(n_315), .Y(n_387) );
AND2x4_ASAP7_75t_L g388 ( .A(n_373), .B(n_3), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_324), .Y(n_389) );
INVx4_ASAP7_75t_L g390 ( .A(n_373), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_265), .Y(n_391) );
AND2x4_ASAP7_75t_L g392 ( .A(n_264), .B(n_3), .Y(n_392) );
NAND2xp33_ASAP7_75t_L g393 ( .A(n_287), .B(n_100), .Y(n_393) );
AND2x4_ASAP7_75t_L g394 ( .A(n_264), .B(n_4), .Y(n_394) );
AND3x2_ASAP7_75t_L g395 ( .A(n_272), .B(n_5), .C(n_6), .Y(n_395) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_324), .Y(n_396) );
INVx6_ASAP7_75t_L g397 ( .A(n_343), .Y(n_397) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_324), .Y(n_398) );
AND2x4_ASAP7_75t_L g399 ( .A(n_300), .B(n_7), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_324), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_266), .Y(n_401) );
INVx4_ASAP7_75t_L g402 ( .A(n_287), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_289), .Y(n_403) );
INVx5_ASAP7_75t_L g404 ( .A(n_343), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_266), .Y(n_405) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_289), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_275), .A2(n_7), .B1(n_8), .B2(n_10), .Y(n_407) );
INVx2_ASAP7_75t_SL g408 ( .A(n_301), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_290), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_387), .B(n_301), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_408), .B(n_262), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_387), .B(n_301), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_408), .B(n_336), .Y(n_413) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_380), .Y(n_414) );
INVx4_ASAP7_75t_L g415 ( .A(n_388), .Y(n_415) );
BUFx2_ASAP7_75t_L g416 ( .A(n_379), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_390), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_390), .B(n_290), .Y(n_418) );
INVx2_ASAP7_75t_SL g419 ( .A(n_390), .Y(n_419) );
INVx4_ASAP7_75t_L g420 ( .A(n_388), .Y(n_420) );
AO22x2_ASAP7_75t_L g421 ( .A1(n_376), .A2(n_279), .B1(n_281), .B2(n_278), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_379), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_387), .B(n_315), .Y(n_423) );
INVx2_ASAP7_75t_SL g424 ( .A(n_390), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_390), .B(n_304), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_381), .Y(n_426) );
INVxp67_ASAP7_75t_L g427 ( .A(n_379), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_408), .B(n_331), .Y(n_428) );
INVx3_ASAP7_75t_L g429 ( .A(n_388), .Y(n_429) );
INVx1_ASAP7_75t_SL g430 ( .A(n_377), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_376), .A2(n_284), .B1(n_334), .B2(n_275), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_381), .Y(n_432) );
INVx4_ASAP7_75t_L g433 ( .A(n_388), .Y(n_433) );
AND2x4_ASAP7_75t_L g434 ( .A(n_376), .B(n_300), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_381), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_388), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g437 ( .A(n_376), .B(n_261), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_406), .Y(n_438) );
OAI22xp33_ASAP7_75t_L g439 ( .A1(n_407), .A2(n_269), .B1(n_274), .B2(n_303), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_376), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_406), .Y(n_441) );
CKINVDCx8_ASAP7_75t_R g442 ( .A(n_392), .Y(n_442) );
CKINVDCx8_ASAP7_75t_R g443 ( .A(n_392), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_406), .Y(n_444) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_380), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_406), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_382), .B(n_304), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_406), .Y(n_448) );
INVx2_ASAP7_75t_SL g449 ( .A(n_404), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_406), .Y(n_450) );
INVx1_ASAP7_75t_SL g451 ( .A(n_377), .Y(n_451) );
INVxp67_ASAP7_75t_SL g452 ( .A(n_385), .Y(n_452) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_380), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_382), .B(n_306), .Y(n_454) );
AND2x6_ASAP7_75t_L g455 ( .A(n_392), .B(n_278), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_406), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_452), .B(n_378), .Y(n_457) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_415), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_426), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_426), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_429), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_432), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_430), .B(n_392), .Y(n_463) );
BUFx2_ASAP7_75t_L g464 ( .A(n_421), .Y(n_464) );
OR2x6_ASAP7_75t_L g465 ( .A(n_421), .B(n_385), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_429), .Y(n_466) );
BUFx3_ASAP7_75t_L g467 ( .A(n_455), .Y(n_467) );
BUFx3_ASAP7_75t_L g468 ( .A(n_455), .Y(n_468) );
INVxp67_ASAP7_75t_L g469 ( .A(n_430), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_432), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_429), .Y(n_471) );
INVx3_ASAP7_75t_L g472 ( .A(n_415), .Y(n_472) );
INVx2_ASAP7_75t_SL g473 ( .A(n_415), .Y(n_473) );
NOR2xp67_ASAP7_75t_L g474 ( .A(n_431), .B(n_378), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_429), .Y(n_475) );
INVx5_ASAP7_75t_L g476 ( .A(n_455), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_435), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_415), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_435), .Y(n_479) );
INVx3_ASAP7_75t_L g480 ( .A(n_420), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_451), .B(n_392), .Y(n_481) );
INVx5_ASAP7_75t_L g482 ( .A(n_455), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_419), .A2(n_393), .B(n_386), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_436), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_436), .Y(n_485) );
AND2x4_ASAP7_75t_L g486 ( .A(n_451), .B(n_394), .Y(n_486) );
BUFx3_ASAP7_75t_L g487 ( .A(n_455), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_423), .Y(n_488) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_420), .Y(n_489) );
AND2x4_ASAP7_75t_L g490 ( .A(n_454), .B(n_394), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_427), .B(n_384), .Y(n_491) );
INVx2_ASAP7_75t_SL g492 ( .A(n_420), .Y(n_492) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_420), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_416), .B(n_394), .Y(n_494) );
INVx3_ASAP7_75t_L g495 ( .A(n_433), .Y(n_495) );
NOR2x1_ASAP7_75t_L g496 ( .A(n_410), .B(n_394), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_433), .B(n_394), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_427), .B(n_399), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_423), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_433), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_411), .B(n_383), .Y(n_501) );
AND3x1_ASAP7_75t_SL g502 ( .A(n_439), .B(n_260), .C(n_259), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_433), .Y(n_503) );
BUFx2_ASAP7_75t_L g504 ( .A(n_421), .Y(n_504) );
AND2x4_ASAP7_75t_L g505 ( .A(n_422), .B(n_399), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_410), .B(n_383), .Y(n_506) );
AND2x2_ASAP7_75t_SL g507 ( .A(n_434), .B(n_399), .Y(n_507) );
AND2x6_ASAP7_75t_L g508 ( .A(n_434), .B(n_399), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_434), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_442), .Y(n_510) );
AND2x6_ASAP7_75t_L g511 ( .A(n_442), .B(n_399), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_418), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_418), .Y(n_513) );
BUFx3_ASAP7_75t_L g514 ( .A(n_455), .Y(n_514) );
INVx3_ASAP7_75t_L g515 ( .A(n_443), .Y(n_515) );
AND2x4_ASAP7_75t_L g516 ( .A(n_412), .B(n_395), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_440), .B(n_386), .Y(n_517) );
INVx4_ASAP7_75t_L g518 ( .A(n_455), .Y(n_518) );
INVx2_ASAP7_75t_SL g519 ( .A(n_455), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_413), .B(n_391), .Y(n_520) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_443), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_428), .B(n_401), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_425), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_437), .B(n_401), .Y(n_524) );
OAI22xp33_ASAP7_75t_L g525 ( .A1(n_431), .A2(n_312), .B1(n_318), .B2(n_303), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_419), .B(n_405), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_419), .B(n_405), .Y(n_527) );
INVx4_ASAP7_75t_L g528 ( .A(n_421), .Y(n_528) );
INVx2_ASAP7_75t_SL g529 ( .A(n_421), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_424), .B(n_261), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_424), .B(n_285), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_438), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_417), .B(n_291), .Y(n_533) );
INVxp67_ASAP7_75t_L g534 ( .A(n_447), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_417), .B(n_291), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_425), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_438), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_447), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_469), .B(n_312), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_534), .B(n_395), .Y(n_540) );
AND2x4_ASAP7_75t_L g541 ( .A(n_488), .B(n_271), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_538), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_474), .A2(n_263), .B1(n_358), .B2(n_313), .Y(n_543) );
AND2x4_ASAP7_75t_L g544 ( .A(n_499), .B(n_316), .Y(n_544) );
INVx2_ASAP7_75t_SL g545 ( .A(n_457), .Y(n_545) );
AND2x4_ASAP7_75t_L g546 ( .A(n_516), .B(n_363), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_512), .B(n_375), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_512), .B(n_375), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_513), .B(n_322), .Y(n_549) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_467), .Y(n_550) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_467), .Y(n_551) );
INVx3_ASAP7_75t_L g552 ( .A(n_458), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_528), .A2(n_366), .B1(n_409), .B2(n_403), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_509), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_513), .B(n_322), .Y(n_555) );
INVx3_ASAP7_75t_L g556 ( .A(n_458), .Y(n_556) );
INVx6_ASAP7_75t_L g557 ( .A(n_458), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_477), .Y(n_558) );
OAI21x1_ASAP7_75t_SL g559 ( .A1(n_528), .A2(n_281), .B(n_279), .Y(n_559) );
INVx4_ASAP7_75t_L g560 ( .A(n_528), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_477), .Y(n_561) );
AND2x4_ASAP7_75t_L g562 ( .A(n_518), .B(n_267), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_498), .Y(n_563) );
INVx4_ASAP7_75t_L g564 ( .A(n_476), .Y(n_564) );
INVx3_ASAP7_75t_L g565 ( .A(n_458), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_498), .Y(n_566) );
INVx5_ASAP7_75t_L g567 ( .A(n_518), .Y(n_567) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_497), .A2(n_393), .B(n_449), .Y(n_568) );
AND2x4_ASAP7_75t_L g569 ( .A(n_518), .B(n_273), .Y(n_569) );
INVx2_ASAP7_75t_SL g570 ( .A(n_505), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_490), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_458), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_489), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_490), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_523), .B(n_341), .Y(n_575) );
CKINVDCx8_ASAP7_75t_R g576 ( .A(n_464), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_504), .A2(n_338), .B1(n_359), .B2(n_334), .Y(n_577) );
INVx3_ASAP7_75t_L g578 ( .A(n_489), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_507), .Y(n_579) );
INVx1_ASAP7_75t_SL g580 ( .A(n_504), .Y(n_580) );
CKINVDCx6p67_ASAP7_75t_R g581 ( .A(n_476), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_506), .Y(n_582) );
INVx1_ASAP7_75t_SL g583 ( .A(n_529), .Y(n_583) );
INVx4_ASAP7_75t_L g584 ( .A(n_476), .Y(n_584) );
AOI22xp33_ASAP7_75t_SL g585 ( .A1(n_529), .A2(n_359), .B1(n_338), .B2(n_341), .Y(n_585) );
BUFx3_ASAP7_75t_L g586 ( .A(n_508), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_536), .B(n_374), .Y(n_587) );
INVxp67_ASAP7_75t_L g588 ( .A(n_511), .Y(n_588) );
INVx4_ASAP7_75t_L g589 ( .A(n_476), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_463), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_489), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_489), .Y(n_592) );
BUFx3_ASAP7_75t_L g593 ( .A(n_508), .Y(n_593) );
NOR2xp67_ASAP7_75t_SL g594 ( .A(n_476), .B(n_286), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_491), .B(n_321), .Y(n_595) );
INVx3_ASAP7_75t_L g596 ( .A(n_489), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_463), .B(n_374), .Y(n_597) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_468), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g599 ( .A1(n_497), .A2(n_449), .B(n_456), .Y(n_599) );
A2O1A1Ixp33_ASAP7_75t_L g600 ( .A1(n_522), .A2(n_409), .B(n_403), .C(n_283), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_494), .Y(n_601) );
INVx5_ASAP7_75t_L g602 ( .A(n_465), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g603 ( .A1(n_505), .A2(n_325), .B1(n_326), .B2(n_323), .C(n_319), .Y(n_603) );
INVx4_ASAP7_75t_L g604 ( .A(n_482), .Y(n_604) );
AND2x4_ASAP7_75t_L g605 ( .A(n_505), .B(n_328), .Y(n_605) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_463), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_481), .Y(n_607) );
INVx3_ASAP7_75t_L g608 ( .A(n_493), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_481), .B(n_403), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_526), .A2(n_449), .B(n_456), .Y(n_610) );
INVx2_ASAP7_75t_SL g611 ( .A(n_496), .Y(n_611) );
AND2x4_ASAP7_75t_L g612 ( .A(n_482), .B(n_333), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_481), .Y(n_613) );
AOI33xp33_ASAP7_75t_L g614 ( .A1(n_525), .A2(n_354), .A3(n_342), .B1(n_335), .B2(n_295), .B3(n_297), .Y(n_614) );
INVxp67_ASAP7_75t_L g615 ( .A(n_511), .Y(n_615) );
NOR2x1_ASAP7_75t_R g616 ( .A(n_482), .B(n_286), .Y(n_616) );
AOI22xp33_ASAP7_75t_SL g617 ( .A1(n_465), .A2(n_277), .B1(n_280), .B2(n_257), .Y(n_617) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_468), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_484), .A2(n_409), .B1(n_277), .B2(n_280), .Y(n_619) );
BUFx6f_ASAP7_75t_L g620 ( .A(n_487), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_515), .B(n_339), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_486), .Y(n_622) );
OAI22xp5_ASAP7_75t_SL g623 ( .A1(n_502), .A2(n_314), .B1(n_317), .B2(n_309), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_511), .A2(n_397), .B1(n_295), .B2(n_297), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_515), .B(n_346), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_493), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_493), .Y(n_627) );
AND2x2_ASAP7_75t_SL g628 ( .A(n_521), .B(n_257), .Y(n_628) );
CKINVDCx8_ASAP7_75t_R g629 ( .A(n_511), .Y(n_629) );
AND2x6_ASAP7_75t_L g630 ( .A(n_514), .B(n_282), .Y(n_630) );
OR2x6_ASAP7_75t_L g631 ( .A(n_514), .B(n_302), .Y(n_631) );
CKINVDCx5p33_ASAP7_75t_R g632 ( .A(n_486), .Y(n_632) );
INVx3_ASAP7_75t_L g633 ( .A(n_493), .Y(n_633) );
A2O1A1Ixp33_ASAP7_75t_L g634 ( .A1(n_501), .A2(n_283), .B(n_288), .C(n_282), .Y(n_634) );
BUFx8_ASAP7_75t_SL g635 ( .A(n_521), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_493), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_527), .A2(n_444), .B(n_441), .Y(n_637) );
AND2x4_ASAP7_75t_L g638 ( .A(n_482), .B(n_302), .Y(n_638) );
BUFx6f_ASAP7_75t_L g639 ( .A(n_482), .Y(n_639) );
OAI221xp5_ASAP7_75t_L g640 ( .A1(n_520), .A2(n_361), .B1(n_365), .B2(n_362), .C(n_357), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_484), .B(n_357), .Y(n_641) );
INVx3_ASAP7_75t_L g642 ( .A(n_472), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_478), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_478), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_485), .B(n_361), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_461), .Y(n_646) );
O2A1O1Ixp33_ASAP7_75t_SL g647 ( .A1(n_485), .A2(n_517), .B(n_483), .C(n_524), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_508), .B(n_362), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_558), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_582), .A2(n_508), .B1(n_511), .B2(n_510), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_561), .Y(n_651) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_545), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_542), .Y(n_653) );
AO31x2_ASAP7_75t_L g654 ( .A1(n_600), .A2(n_400), .A3(n_389), .B(n_459), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_641), .Y(n_655) );
INVx1_ASAP7_75t_SL g656 ( .A(n_635), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_646), .Y(n_657) );
NAND2xp33_ASAP7_75t_L g658 ( .A(n_583), .B(n_521), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_643), .Y(n_659) );
BUFx3_ASAP7_75t_L g660 ( .A(n_639), .Y(n_660) );
BUFx3_ASAP7_75t_L g661 ( .A(n_639), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_617), .A2(n_462), .B1(n_470), .B2(n_460), .Y(n_662) );
BUFx6f_ASAP7_75t_L g663 ( .A(n_567), .Y(n_663) );
BUFx6f_ASAP7_75t_L g664 ( .A(n_567), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_617), .A2(n_479), .B1(n_519), .B2(n_533), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_547), .B(n_508), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_553), .A2(n_519), .B1(n_535), .B2(n_531), .Y(n_667) );
BUFx4_ASAP7_75t_SL g668 ( .A(n_631), .Y(n_668) );
BUFx3_ASAP7_75t_L g669 ( .A(n_639), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_644), .Y(n_670) );
CKINVDCx11_ASAP7_75t_R g671 ( .A(n_576), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_601), .A2(n_508), .B1(n_466), .B2(n_475), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_547), .B(n_530), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_579), .A2(n_466), .B1(n_475), .B2(n_471), .Y(n_674) );
OAI222xp33_ASAP7_75t_L g675 ( .A1(n_585), .A2(n_371), .B1(n_367), .B2(n_365), .C1(n_351), .C2(n_320), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_539), .B(n_500), .Y(n_676) );
AND2x4_ASAP7_75t_L g677 ( .A(n_560), .B(n_472), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_641), .Y(n_678) );
AOI22xp33_ASAP7_75t_SL g679 ( .A1(n_628), .A2(n_320), .B1(n_353), .B2(n_337), .Y(n_679) );
O2A1O1Ixp33_ASAP7_75t_SL g680 ( .A1(n_634), .A2(n_444), .B(n_446), .C(n_441), .Y(n_680) );
OAI21xp5_ASAP7_75t_L g681 ( .A1(n_568), .A2(n_503), .B(n_492), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_645), .Y(n_682) );
AND2x4_ASAP7_75t_L g683 ( .A(n_586), .B(n_472), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_647), .A2(n_473), .B(n_480), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_645), .Y(n_685) );
AND2x4_ASAP7_75t_L g686 ( .A(n_593), .B(n_480), .Y(n_686) );
AND2x4_ASAP7_75t_L g687 ( .A(n_567), .B(n_480), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_648), .Y(n_688) );
INVx3_ASAP7_75t_L g689 ( .A(n_629), .Y(n_689) );
AND2x4_ASAP7_75t_L g690 ( .A(n_588), .B(n_495), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_605), .A2(n_287), .B1(n_495), .B2(n_351), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_580), .A2(n_473), .B1(n_353), .B2(n_355), .Y(n_692) );
CKINVDCx5p33_ASAP7_75t_R g693 ( .A(n_623), .Y(n_693) );
OAI22xp33_ASAP7_75t_L g694 ( .A1(n_543), .A2(n_287), .B1(n_397), .B2(n_292), .Y(n_694) );
A2O1A1Ixp33_ASAP7_75t_L g695 ( .A1(n_614), .A2(n_288), .B(n_293), .C(n_292), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_548), .B(n_397), .Y(n_696) );
INVx3_ASAP7_75t_L g697 ( .A(n_564), .Y(n_697) );
AOI21xp33_ASAP7_75t_L g698 ( .A1(n_540), .A2(n_350), .B(n_310), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_605), .Y(n_699) );
INVx5_ASAP7_75t_L g700 ( .A(n_630), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_541), .Y(n_701) );
BUFx6f_ASAP7_75t_L g702 ( .A(n_550), .Y(n_702) );
INVx4_ASAP7_75t_L g703 ( .A(n_630), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_607), .A2(n_406), .B1(n_402), .B2(n_294), .Y(n_704) );
A2O1A1Ixp33_ASAP7_75t_L g705 ( .A1(n_613), .A2(n_293), .B(n_296), .C(n_294), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_549), .A2(n_298), .B1(n_299), .B2(n_296), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_549), .A2(n_369), .B1(n_372), .B2(n_364), .Y(n_707) );
NAND2x1p5_ASAP7_75t_L g708 ( .A(n_602), .B(n_364), .Y(n_708) );
OAI22xp33_ASAP7_75t_SL g709 ( .A1(n_632), .A2(n_372), .B1(n_369), .B2(n_270), .Y(n_709) );
AND2x4_ASAP7_75t_L g710 ( .A(n_588), .B(n_276), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_555), .B(n_402), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_555), .A2(n_307), .B1(n_308), .B2(n_268), .Y(n_712) );
BUFx3_ASAP7_75t_L g713 ( .A(n_557), .Y(n_713) );
CKINVDCx5p33_ASAP7_75t_R g714 ( .A(n_546), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_572), .Y(n_715) );
INVx2_ASAP7_75t_L g716 ( .A(n_573), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_637), .A2(n_537), .B(n_532), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_585), .B(n_402), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_591), .Y(n_719) );
CKINVDCx11_ASAP7_75t_R g720 ( .A(n_581), .Y(n_720) );
INVx4_ASAP7_75t_L g721 ( .A(n_630), .Y(n_721) );
BUFx2_ASAP7_75t_L g722 ( .A(n_630), .Y(n_722) );
CKINVDCx11_ASAP7_75t_R g723 ( .A(n_546), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_592), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_540), .B(n_327), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_626), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_622), .A2(n_402), .B1(n_329), .B2(n_332), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_595), .B(n_10), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g729 ( .A1(n_637), .A2(n_537), .B(n_532), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_541), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_571), .A2(n_345), .B1(n_347), .B2(n_340), .Y(n_731) );
A2O1A1Ixp33_ASAP7_75t_L g732 ( .A1(n_640), .A2(n_330), .B(n_356), .C(n_305), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_574), .A2(n_349), .B1(n_352), .B2(n_348), .Y(n_733) );
INVx3_ASAP7_75t_L g734 ( .A(n_564), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_627), .Y(n_735) );
BUFx3_ASAP7_75t_L g736 ( .A(n_557), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_577), .B(n_11), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_544), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_590), .A2(n_606), .B1(n_563), .B2(n_566), .Y(n_739) );
AND2x4_ASAP7_75t_L g740 ( .A(n_615), .B(n_305), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_636), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_552), .Y(n_742) );
INVx1_ASAP7_75t_SL g743 ( .A(n_638), .Y(n_743) );
NOR2xp33_ASAP7_75t_SL g744 ( .A(n_616), .B(n_404), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_575), .B(n_12), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_587), .B(n_12), .Y(n_746) );
OA21x2_ASAP7_75t_L g747 ( .A1(n_610), .A2(n_446), .B(n_438), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_554), .Y(n_748) );
INVx5_ASAP7_75t_L g749 ( .A(n_630), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_597), .B(n_570), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_603), .A2(n_368), .B1(n_360), .B2(n_389), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_603), .A2(n_389), .B1(n_400), .B2(n_404), .Y(n_752) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_597), .A2(n_404), .B1(n_450), .B2(n_448), .Y(n_753) );
AND2x2_ASAP7_75t_L g754 ( .A(n_562), .B(n_13), .Y(n_754) );
BUFx3_ASAP7_75t_L g755 ( .A(n_557), .Y(n_755) );
AO21x2_ASAP7_75t_L g756 ( .A1(n_684), .A2(n_559), .B(n_609), .Y(n_756) );
A2O1A1Ixp33_ASAP7_75t_L g757 ( .A1(n_655), .A2(n_625), .B(n_621), .C(n_624), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_737), .A2(n_619), .B1(n_611), .B2(n_569), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_678), .A2(n_619), .B1(n_569), .B2(n_562), .Y(n_759) );
AOI221xp5_ASAP7_75t_L g760 ( .A1(n_675), .A2(n_568), .B1(n_638), .B2(n_612), .C(n_642), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_662), .A2(n_612), .B1(n_551), .B2(n_598), .Y(n_761) );
INVx4_ASAP7_75t_L g762 ( .A(n_720), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_682), .A2(n_642), .B1(n_556), .B2(n_565), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_653), .Y(n_764) );
OAI221xp5_ASAP7_75t_L g765 ( .A1(n_725), .A2(n_610), .B1(n_599), .B2(n_633), .C(n_565), .Y(n_765) );
OAI22xp5_ASAP7_75t_L g766 ( .A1(n_685), .A2(n_551), .B1(n_598), .B2(n_550), .Y(n_766) );
BUFx6f_ASAP7_75t_SL g767 ( .A(n_668), .Y(n_767) );
INVx2_ASAP7_75t_L g768 ( .A(n_649), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_745), .A2(n_596), .B1(n_608), .B2(n_578), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_701), .Y(n_770) );
NAND3xp33_ASAP7_75t_L g771 ( .A(n_732), .B(n_400), .C(n_594), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_730), .Y(n_772) );
OAI221xp5_ASAP7_75t_L g773 ( .A1(n_695), .A2(n_604), .B1(n_589), .B2(n_584), .C(n_598), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_728), .A2(n_620), .B1(n_618), .B2(n_589), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_738), .Y(n_775) );
AND2x4_ASAP7_75t_L g776 ( .A(n_703), .B(n_14), .Y(n_776) );
BUFx2_ASAP7_75t_L g777 ( .A(n_652), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_665), .A2(n_404), .B1(n_450), .B2(n_448), .Y(n_778) );
OAI22xp5_ASAP7_75t_L g779 ( .A1(n_667), .A2(n_404), .B1(n_448), .B2(n_398), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_746), .A2(n_398), .B1(n_396), .B2(n_380), .Y(n_780) );
AND2x4_ASAP7_75t_L g781 ( .A(n_703), .B(n_14), .Y(n_781) );
INVx3_ASAP7_75t_L g782 ( .A(n_721), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_688), .A2(n_398), .B1(n_396), .B2(n_380), .Y(n_783) );
AOI221xp5_ASAP7_75t_L g784 ( .A1(n_712), .A2(n_398), .B1(n_396), .B2(n_380), .C(n_453), .Y(n_784) );
BUFx12f_ASAP7_75t_L g785 ( .A(n_671), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_671), .Y(n_786) );
AOI222xp33_ASAP7_75t_L g787 ( .A1(n_723), .A2(n_396), .B1(n_398), .B2(n_19), .C1(n_20), .C2(n_21), .Y(n_787) );
AOI22xp33_ASAP7_75t_SL g788 ( .A1(n_721), .A2(n_396), .B1(n_398), .B2(n_19), .Y(n_788) );
BUFx12f_ASAP7_75t_L g789 ( .A(n_714), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_748), .B(n_17), .Y(n_790) );
AOI21xp5_ASAP7_75t_L g791 ( .A1(n_717), .A2(n_729), .B(n_673), .Y(n_791) );
OAI22xp33_ASAP7_75t_L g792 ( .A1(n_700), .A2(n_17), .B1(n_18), .B2(n_22), .Y(n_792) );
AOI21xp33_ASAP7_75t_L g793 ( .A1(n_718), .A2(n_23), .B(n_24), .Y(n_793) );
O2A1O1Ixp33_ASAP7_75t_SL g794 ( .A1(n_732), .A2(n_122), .B(n_256), .C(n_255), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_676), .Y(n_795) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_691), .A2(n_25), .B1(n_26), .B2(n_27), .Y(n_796) );
CKINVDCx11_ASAP7_75t_R g797 ( .A(n_656), .Y(n_797) );
HB1xp67_ASAP7_75t_L g798 ( .A(n_754), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_666), .A2(n_453), .B1(n_445), .B2(n_414), .Y(n_799) );
AOI322xp5_ASAP7_75t_L g800 ( .A1(n_693), .A2(n_29), .A3(n_30), .B1(n_31), .B2(n_32), .C1(n_34), .C2(n_35), .Y(n_800) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_708), .A2(n_29), .B1(n_30), .B2(n_31), .Y(n_801) );
BUFx4f_ASAP7_75t_SL g802 ( .A(n_663), .Y(n_802) );
AOI222xp33_ASAP7_75t_L g803 ( .A1(n_699), .A2(n_34), .B1(n_35), .B2(n_36), .C1(n_37), .C2(n_38), .Y(n_803) );
OAI21xp5_ASAP7_75t_L g804 ( .A1(n_705), .A2(n_39), .B(n_40), .Y(n_804) );
AND2x4_ASAP7_75t_L g805 ( .A(n_749), .B(n_40), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_679), .B(n_41), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_695), .B(n_44), .Y(n_807) );
OAI22xp5_ASAP7_75t_L g808 ( .A1(n_749), .A2(n_46), .B1(n_47), .B2(n_48), .Y(n_808) );
AOI21xp5_ASAP7_75t_L g809 ( .A1(n_696), .A2(n_445), .B(n_414), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_651), .A2(n_453), .B1(n_445), .B2(n_414), .Y(n_810) );
AOI222xp33_ASAP7_75t_L g811 ( .A1(n_750), .A2(n_48), .B1(n_49), .B2(n_50), .C1(n_51), .C2(n_53), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_694), .A2(n_453), .B1(n_445), .B2(n_414), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_706), .A2(n_445), .B1(n_414), .B2(n_56), .Y(n_813) );
AOI222xp33_ASAP7_75t_L g814 ( .A1(n_751), .A2(n_54), .B1(n_55), .B2(n_56), .C1(n_57), .C2(n_58), .Y(n_814) );
OAI211xp5_ASAP7_75t_L g815 ( .A1(n_698), .A2(n_57), .B(n_59), .C(n_60), .Y(n_815) );
INVx2_ASAP7_75t_L g816 ( .A(n_657), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_657), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_707), .A2(n_61), .B1(n_62), .B2(n_63), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_710), .A2(n_65), .B1(n_66), .B2(n_67), .Y(n_819) );
OR2x6_ASAP7_75t_L g820 ( .A(n_722), .B(n_66), .Y(n_820) );
OAI21x1_ASAP7_75t_SL g821 ( .A1(n_650), .A2(n_67), .B(n_68), .Y(n_821) );
INVx2_ASAP7_75t_L g822 ( .A(n_659), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_710), .A2(n_69), .B1(n_70), .B2(n_71), .Y(n_823) );
OAI22xp33_ASAP7_75t_L g824 ( .A1(n_744), .A2(n_70), .B1(n_73), .B2(n_74), .Y(n_824) );
OAI211xp5_ASAP7_75t_L g825 ( .A1(n_731), .A2(n_73), .B(n_74), .C(n_75), .Y(n_825) );
OA21x2_ASAP7_75t_L g826 ( .A1(n_681), .A2(n_152), .B(n_253), .Y(n_826) );
OAI22xp5_ASAP7_75t_L g827 ( .A1(n_743), .A2(n_76), .B1(n_77), .B2(n_78), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_710), .A2(n_76), .B1(n_79), .B2(n_80), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_709), .A2(n_79), .B1(n_81), .B2(n_82), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_659), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_711), .Y(n_831) );
INVx4_ASAP7_75t_L g832 ( .A(n_663), .Y(n_832) );
O2A1O1Ixp33_ASAP7_75t_L g833 ( .A1(n_705), .A2(n_81), .B(n_83), .C(n_84), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_740), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_740), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_733), .A2(n_86), .B1(n_87), .B2(n_88), .Y(n_836) );
AOI221xp5_ASAP7_75t_L g837 ( .A1(n_733), .A2(n_89), .B1(n_90), .B2(n_91), .C(n_92), .Y(n_837) );
INVxp67_ASAP7_75t_L g838 ( .A(n_692), .Y(n_838) );
AOI21xp5_ASAP7_75t_L g839 ( .A1(n_680), .A2(n_164), .B(n_249), .Y(n_839) );
OR2x2_ASAP7_75t_L g840 ( .A(n_670), .B(n_89), .Y(n_840) );
OAI22xp5_ASAP7_75t_L g841 ( .A1(n_650), .A2(n_92), .B1(n_93), .B2(n_94), .Y(n_841) );
OAI22xp5_ASAP7_75t_L g842 ( .A1(n_672), .A2(n_93), .B1(n_95), .B2(n_96), .Y(n_842) );
AND2x2_ASAP7_75t_L g843 ( .A(n_739), .B(n_95), .Y(n_843) );
BUFx2_ASAP7_75t_L g844 ( .A(n_755), .Y(n_844) );
AOI222xp33_ASAP7_75t_L g845 ( .A1(n_752), .A2(n_97), .B1(n_98), .B2(n_101), .C1(n_102), .C2(n_104), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_740), .Y(n_846) );
BUFx3_ASAP7_75t_L g847 ( .A(n_663), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_764), .Y(n_848) );
INVx2_ASAP7_75t_L g849 ( .A(n_816), .Y(n_849) );
INVx2_ASAP7_75t_L g850 ( .A(n_817), .Y(n_850) );
OR2x6_ASAP7_75t_L g851 ( .A(n_820), .B(n_663), .Y(n_851) );
INVx2_ASAP7_75t_L g852 ( .A(n_768), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_795), .B(n_752), .Y(n_853) );
HB1xp67_ASAP7_75t_L g854 ( .A(n_777), .Y(n_854) );
AND2x2_ASAP7_75t_L g855 ( .A(n_822), .B(n_654), .Y(n_855) );
BUFx6f_ASAP7_75t_L g856 ( .A(n_847), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_770), .Y(n_857) );
OR2x2_ASAP7_75t_L g858 ( .A(n_798), .B(n_715), .Y(n_858) );
OAI22xp5_ASAP7_75t_L g859 ( .A1(n_759), .A2(n_672), .B1(n_674), .B2(n_727), .Y(n_859) );
INVx2_ASAP7_75t_L g860 ( .A(n_830), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_758), .A2(n_674), .B1(n_690), .B2(n_689), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_772), .Y(n_862) );
OAI211xp5_ASAP7_75t_L g863 ( .A1(n_811), .A2(n_704), .B(n_753), .C(n_680), .Y(n_863) );
AO221x2_ASAP7_75t_L g864 ( .A1(n_792), .A2(n_742), .B1(n_741), .B2(n_735), .C(n_726), .Y(n_864) );
AOI22xp5_ASAP7_75t_L g865 ( .A1(n_759), .A2(n_690), .B1(n_677), .B2(n_686), .Y(n_865) );
CKINVDCx20_ASAP7_75t_R g866 ( .A(n_786), .Y(n_866) );
NOR2xp33_ASAP7_75t_L g867 ( .A(n_838), .B(n_683), .Y(n_867) );
INVx3_ASAP7_75t_L g868 ( .A(n_802), .Y(n_868) );
AND2x4_ASAP7_75t_SL g869 ( .A(n_762), .B(n_664), .Y(n_869) );
AND2x4_ASAP7_75t_SL g870 ( .A(n_762), .B(n_664), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_775), .Y(n_871) );
AOI222xp33_ASAP7_75t_L g872 ( .A1(n_767), .A2(n_704), .B1(n_683), .B2(n_686), .C1(n_690), .C2(n_677), .Y(n_872) );
AOI211xp5_ASAP7_75t_L g873 ( .A1(n_824), .A2(n_683), .B(n_686), .C(n_677), .Y(n_873) );
NAND3xp33_ASAP7_75t_L g874 ( .A(n_787), .B(n_658), .C(n_742), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_843), .A2(n_747), .B1(n_697), .B2(n_734), .Y(n_875) );
INVx2_ASAP7_75t_L g876 ( .A(n_826), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_790), .Y(n_877) );
INVx2_ASAP7_75t_L g878 ( .A(n_826), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_804), .A2(n_747), .B1(n_734), .B2(n_713), .Y(n_879) );
OAI322xp33_ASAP7_75t_L g880 ( .A1(n_824), .A2(n_741), .A3(n_735), .B1(n_726), .B2(n_724), .C1(n_719), .C2(n_716), .Y(n_880) );
AOI221xp5_ASAP7_75t_L g881 ( .A1(n_833), .A2(n_687), .B1(n_715), .B2(n_716), .C(n_724), .Y(n_881) );
NAND3xp33_ASAP7_75t_L g882 ( .A(n_815), .B(n_755), .C(n_713), .Y(n_882) );
AND2x2_ASAP7_75t_L g883 ( .A(n_776), .B(n_654), .Y(n_883) );
INVx2_ASAP7_75t_L g884 ( .A(n_826), .Y(n_884) );
INVx2_ASAP7_75t_SL g885 ( .A(n_832), .Y(n_885) );
HB1xp67_ASAP7_75t_L g886 ( .A(n_781), .Y(n_886) );
AND2x2_ASAP7_75t_L g887 ( .A(n_806), .B(n_800), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_831), .B(n_736), .Y(n_888) );
AND2x2_ASAP7_75t_L g889 ( .A(n_840), .B(n_654), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_803), .B(n_687), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_805), .Y(n_891) );
AOI222xp33_ASAP7_75t_L g892 ( .A1(n_785), .A2(n_669), .B1(n_661), .B2(n_660), .C1(n_702), .C2(n_747), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_801), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_829), .A2(n_669), .B1(n_661), .B2(n_660), .Y(n_894) );
AOI21xp5_ASAP7_75t_L g895 ( .A1(n_791), .A2(n_702), .B(n_112), .Y(n_895) );
OR2x2_ASAP7_75t_L g896 ( .A(n_844), .B(n_702), .Y(n_896) );
OAI22xp5_ASAP7_75t_L g897 ( .A1(n_813), .A2(n_702), .B1(n_113), .B2(n_115), .Y(n_897) );
OAI22xp5_ASAP7_75t_L g898 ( .A1(n_813), .A2(n_110), .B1(n_116), .B2(n_119), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_814), .A2(n_120), .B1(n_121), .B2(n_123), .Y(n_899) );
OAI31xp33_ASAP7_75t_L g900 ( .A1(n_825), .A2(n_126), .A3(n_127), .B(n_128), .Y(n_900) );
OAI222xp33_ASAP7_75t_L g901 ( .A1(n_819), .A2(n_129), .B1(n_130), .B2(n_132), .C1(n_133), .C2(n_134), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_837), .A2(n_136), .B1(n_138), .B2(n_139), .Y(n_902) );
AOI22xp5_ASAP7_75t_L g903 ( .A1(n_841), .A2(n_140), .B1(n_142), .B2(n_143), .Y(n_903) );
AO21x2_ASAP7_75t_L g904 ( .A1(n_809), .A2(n_146), .B(n_148), .Y(n_904) );
AOI22xp5_ASAP7_75t_L g905 ( .A1(n_796), .A2(n_149), .B1(n_150), .B2(n_151), .Y(n_905) );
BUFx3_ASAP7_75t_L g906 ( .A(n_847), .Y(n_906) );
AO21x2_ASAP7_75t_L g907 ( .A1(n_839), .A2(n_153), .B(n_154), .Y(n_907) );
AND2x4_ASAP7_75t_SL g908 ( .A(n_782), .B(n_254), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_757), .B(n_156), .Y(n_909) );
INVx2_ASAP7_75t_SL g910 ( .A(n_782), .Y(n_910) );
INVx2_ASAP7_75t_L g911 ( .A(n_834), .Y(n_911) );
AOI22xp5_ASAP7_75t_L g912 ( .A1(n_842), .A2(n_158), .B1(n_162), .B2(n_163), .Y(n_912) );
AOI22xp33_ASAP7_75t_SL g913 ( .A1(n_821), .A2(n_167), .B1(n_172), .B2(n_173), .Y(n_913) );
INVx2_ASAP7_75t_L g914 ( .A(n_835), .Y(n_914) );
NAND3xp33_ASAP7_75t_SL g915 ( .A(n_823), .B(n_174), .C(n_176), .Y(n_915) );
INVx2_ASAP7_75t_L g916 ( .A(n_846), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_807), .Y(n_917) );
INVx2_ASAP7_75t_L g918 ( .A(n_756), .Y(n_918) );
OA21x2_ASAP7_75t_L g919 ( .A1(n_778), .A2(n_177), .B(n_180), .Y(n_919) );
OAI33xp33_ASAP7_75t_L g920 ( .A1(n_827), .A2(n_183), .A3(n_184), .B1(n_186), .B2(n_187), .B3(n_189), .Y(n_920) );
AOI221xp5_ASAP7_75t_L g921 ( .A1(n_793), .A2(n_190), .B1(n_192), .B2(n_194), .C(n_195), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_818), .B(n_196), .Y(n_922) );
AOI221xp5_ASAP7_75t_L g923 ( .A1(n_818), .A2(n_197), .B1(n_200), .B2(n_202), .C(n_203), .Y(n_923) );
INVx3_ASAP7_75t_L g924 ( .A(n_756), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_808), .Y(n_925) );
AOI33xp33_ASAP7_75t_L g926 ( .A1(n_836), .A2(n_246), .A3(n_210), .B1(n_211), .B2(n_213), .B3(n_214), .Y(n_926) );
INVx2_ASAP7_75t_L g927 ( .A(n_765), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_836), .A2(n_204), .B1(n_215), .B2(n_217), .Y(n_928) );
AOI21xp5_ASAP7_75t_L g929 ( .A1(n_880), .A2(n_761), .B(n_794), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_848), .Y(n_930) );
AND2x2_ASAP7_75t_L g931 ( .A(n_850), .B(n_823), .Y(n_931) );
NAND3xp33_ASAP7_75t_L g932 ( .A(n_892), .B(n_828), .C(n_845), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_887), .B(n_828), .Y(n_933) );
HB1xp67_ASAP7_75t_L g934 ( .A(n_854), .Y(n_934) );
NOR2xp33_ASAP7_75t_L g935 ( .A(n_890), .B(n_789), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_893), .A2(n_760), .B1(n_788), .B2(n_773), .Y(n_936) );
NOR2xp33_ASAP7_75t_SL g937 ( .A(n_866), .B(n_797), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_857), .B(n_862), .Y(n_938) );
OAI33xp33_ASAP7_75t_L g939 ( .A1(n_871), .A2(n_779), .A3(n_766), .B1(n_771), .B2(n_769), .B3(n_794), .Y(n_939) );
AND2x2_ASAP7_75t_L g940 ( .A(n_883), .B(n_763), .Y(n_940) );
AND2x2_ASAP7_75t_L g941 ( .A(n_855), .B(n_889), .Y(n_941) );
BUFx2_ASAP7_75t_L g942 ( .A(n_885), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_858), .Y(n_943) );
INVx4_ASAP7_75t_L g944 ( .A(n_851), .Y(n_944) );
BUFx2_ASAP7_75t_L g945 ( .A(n_885), .Y(n_945) );
NAND4xp25_ASAP7_75t_L g946 ( .A(n_867), .B(n_780), .C(n_774), .D(n_784), .Y(n_946) );
OR2x2_ASAP7_75t_L g947 ( .A(n_911), .B(n_799), .Y(n_947) );
INVx2_ASAP7_75t_L g948 ( .A(n_860), .Y(n_948) );
OR2x2_ASAP7_75t_L g949 ( .A(n_849), .B(n_783), .Y(n_949) );
AOI33xp33_ASAP7_75t_L g950 ( .A1(n_877), .A2(n_812), .A3(n_810), .B1(n_222), .B2(n_224), .B3(n_226), .Y(n_950) );
INVx1_ASAP7_75t_SL g951 ( .A(n_869), .Y(n_951) );
AND2x2_ASAP7_75t_L g952 ( .A(n_852), .B(n_219), .Y(n_952) );
INVx2_ASAP7_75t_L g953 ( .A(n_852), .Y(n_953) );
NOR2xp33_ASAP7_75t_L g954 ( .A(n_867), .B(n_231), .Y(n_954) );
AND2x4_ASAP7_75t_L g955 ( .A(n_851), .B(n_234), .Y(n_955) );
AND2x2_ASAP7_75t_L g956 ( .A(n_914), .B(n_235), .Y(n_956) );
INVx2_ASAP7_75t_L g957 ( .A(n_918), .Y(n_957) );
OAI33xp33_ASAP7_75t_L g958 ( .A1(n_925), .A2(n_236), .A3(n_240), .B1(n_242), .B2(n_243), .B3(n_917), .Y(n_958) );
OAI33xp33_ASAP7_75t_L g959 ( .A1(n_888), .A2(n_891), .A3(n_859), .B1(n_853), .B2(n_898), .B3(n_909), .Y(n_959) );
INVxp67_ASAP7_75t_L g960 ( .A(n_886), .Y(n_960) );
INVx4_ASAP7_75t_SL g961 ( .A(n_851), .Y(n_961) );
INVx2_ASAP7_75t_L g962 ( .A(n_918), .Y(n_962) );
OAI221xp5_ASAP7_75t_L g963 ( .A1(n_899), .A2(n_894), .B1(n_861), .B2(n_873), .C(n_872), .Y(n_963) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_916), .B(n_861), .Y(n_964) );
OAI33xp33_ASAP7_75t_L g965 ( .A1(n_927), .A2(n_922), .A3(n_897), .B1(n_874), .B2(n_916), .B3(n_896), .Y(n_965) );
OAI321xp33_ASAP7_75t_L g966 ( .A1(n_894), .A2(n_928), .A3(n_915), .B1(n_882), .B2(n_927), .C(n_879), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_910), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g968 ( .A(n_865), .B(n_870), .Y(n_968) );
AND2x2_ASAP7_75t_L g969 ( .A(n_875), .B(n_864), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_910), .Y(n_970) );
NOR3xp33_ASAP7_75t_SL g971 ( .A(n_901), .B(n_863), .C(n_920), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_875), .B(n_864), .Y(n_972) );
AND2x2_ASAP7_75t_L g973 ( .A(n_864), .B(n_924), .Y(n_973) );
INVx1_ASAP7_75t_L g974 ( .A(n_908), .Y(n_974) );
NOR2xp33_ASAP7_75t_L g975 ( .A(n_868), .B(n_870), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_906), .B(n_856), .Y(n_976) );
NOR2x1_ASAP7_75t_L g977 ( .A(n_942), .B(n_868), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_941), .B(n_878), .Y(n_978) );
BUFx3_ASAP7_75t_L g979 ( .A(n_945), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g980 ( .A(n_943), .B(n_868), .Y(n_980) );
AND2x2_ASAP7_75t_L g981 ( .A(n_940), .B(n_876), .Y(n_981) );
OR2x2_ASAP7_75t_L g982 ( .A(n_964), .B(n_884), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_948), .Y(n_983) );
INVx2_ASAP7_75t_L g984 ( .A(n_957), .Y(n_984) );
NOR2xp33_ASAP7_75t_L g985 ( .A(n_937), .B(n_866), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g986 ( .A(n_930), .B(n_881), .Y(n_986) );
AND2x2_ASAP7_75t_L g987 ( .A(n_940), .B(n_878), .Y(n_987) );
NAND2x1p5_ASAP7_75t_L g988 ( .A(n_955), .B(n_919), .Y(n_988) );
OAI21xp5_ASAP7_75t_L g989 ( .A1(n_932), .A2(n_902), .B(n_926), .Y(n_989) );
INVxp33_ASAP7_75t_L g990 ( .A(n_975), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_953), .Y(n_991) );
OAI31xp33_ASAP7_75t_SL g992 ( .A1(n_963), .A2(n_913), .A3(n_923), .B(n_921), .Y(n_992) );
OR2x2_ASAP7_75t_L g993 ( .A(n_934), .B(n_904), .Y(n_993) );
NOR2xp33_ASAP7_75t_L g994 ( .A(n_935), .B(n_905), .Y(n_994) );
BUFx2_ASAP7_75t_L g995 ( .A(n_976), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g996 ( .A(n_938), .B(n_900), .Y(n_996) );
OAI322xp33_ASAP7_75t_L g997 ( .A1(n_933), .A2(n_895), .A3(n_903), .B1(n_907), .B2(n_912), .C1(n_935), .C2(n_960), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_953), .Y(n_998) );
OR2x2_ASAP7_75t_L g999 ( .A(n_969), .B(n_972), .Y(n_999) );
INVx2_ASAP7_75t_L g1000 ( .A(n_957), .Y(n_1000) );
AOI322xp5_ASAP7_75t_L g1001 ( .A1(n_971), .A2(n_974), .A3(n_954), .B1(n_931), .B2(n_975), .C1(n_936), .C2(n_955), .Y(n_1001) );
INVx1_ASAP7_75t_SL g1002 ( .A(n_951), .Y(n_1002) );
NAND3xp33_ASAP7_75t_L g1003 ( .A(n_950), .B(n_970), .C(n_967), .Y(n_1003) );
AND2x4_ASAP7_75t_L g1004 ( .A(n_973), .B(n_961), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1005 ( .A(n_968), .B(n_954), .Y(n_1005) );
NAND4xp25_ASAP7_75t_L g1006 ( .A(n_946), .B(n_929), .C(n_950), .D(n_944), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_962), .B(n_947), .Y(n_1007) );
AOI221xp5_ASAP7_75t_L g1008 ( .A1(n_959), .A2(n_965), .B1(n_958), .B2(n_966), .C(n_939), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_980), .Y(n_1009) );
OR2x2_ASAP7_75t_L g1010 ( .A(n_995), .B(n_949), .Y(n_1010) );
INVx2_ASAP7_75t_L g1011 ( .A(n_984), .Y(n_1011) );
OR2x2_ASAP7_75t_L g1012 ( .A(n_999), .B(n_952), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_978), .B(n_956), .Y(n_1013) );
AND2x2_ASAP7_75t_L g1014 ( .A(n_978), .B(n_952), .Y(n_1014) );
INVx1_ASAP7_75t_L g1015 ( .A(n_979), .Y(n_1015) );
NAND2x1_ASAP7_75t_L g1016 ( .A(n_977), .B(n_1004), .Y(n_1016) );
NOR3xp33_ASAP7_75t_L g1017 ( .A(n_1006), .B(n_1008), .C(n_989), .Y(n_1017) );
NAND2xp5_ASAP7_75t_L g1018 ( .A(n_1007), .B(n_981), .Y(n_1018) );
OAI31xp33_ASAP7_75t_L g1019 ( .A1(n_994), .A2(n_988), .A3(n_985), .B(n_1003), .Y(n_1019) );
NOR3xp33_ASAP7_75t_L g1020 ( .A(n_997), .B(n_996), .C(n_1002), .Y(n_1020) );
NAND4xp25_ASAP7_75t_L g1021 ( .A(n_1001), .B(n_992), .C(n_1005), .D(n_986), .Y(n_1021) );
NAND4xp25_ASAP7_75t_L g1022 ( .A(n_1017), .B(n_1001), .C(n_992), .D(n_993), .Y(n_1022) );
NOR2xp33_ASAP7_75t_L g1023 ( .A(n_1021), .B(n_990), .Y(n_1023) );
INVx2_ASAP7_75t_L g1024 ( .A(n_1011), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_1009), .Y(n_1025) );
NAND2xp5_ASAP7_75t_SL g1026 ( .A(n_1019), .B(n_988), .Y(n_1026) );
NOR3xp33_ASAP7_75t_L g1027 ( .A(n_1020), .B(n_997), .C(n_993), .Y(n_1027) );
INVx2_ASAP7_75t_SL g1028 ( .A(n_1016), .Y(n_1028) );
OR2x2_ASAP7_75t_L g1029 ( .A(n_1018), .B(n_982), .Y(n_1029) );
OR2x2_ASAP7_75t_L g1030 ( .A(n_1010), .B(n_987), .Y(n_1030) );
INVx1_ASAP7_75t_SL g1031 ( .A(n_1014), .Y(n_1031) );
NOR5xp2_ASAP7_75t_L g1032 ( .A(n_1015), .B(n_983), .C(n_991), .D(n_998), .E(n_1000), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_1022), .A2(n_1023), .B1(n_1026), .B2(n_1027), .Y(n_1033) );
OR2x2_ASAP7_75t_L g1034 ( .A(n_1029), .B(n_1030), .Y(n_1034) );
INVx1_ASAP7_75t_L g1035 ( .A(n_1029), .Y(n_1035) );
OA22x2_ASAP7_75t_L g1036 ( .A1(n_1033), .A2(n_1028), .B1(n_1031), .B2(n_1025), .Y(n_1036) );
XOR2xp5_ASAP7_75t_L g1037 ( .A(n_1035), .B(n_1012), .Y(n_1037) );
NAND3xp33_ASAP7_75t_SL g1038 ( .A(n_1036), .B(n_1032), .C(n_1034), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_1038), .Y(n_1039) );
NAND2xp5_ASAP7_75t_L g1040 ( .A(n_1039), .B(n_1037), .Y(n_1040) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1040), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1041), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_1042), .Y(n_1043) );
AO21x2_ASAP7_75t_L g1044 ( .A1(n_1043), .A2(n_1024), .B(n_1013), .Y(n_1044) );
endmodule