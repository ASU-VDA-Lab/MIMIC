module fake_jpeg_20080_n_175 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_175);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_127;
wire n_76;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_61;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_22),
.B(n_5),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_24),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_48),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_23),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_18),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_44),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_5),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_28),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_9),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_12),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_15),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_42),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_1),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_9),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_81),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_19),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_68),
.Y(n_97)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

INVx4_ASAP7_75t_SL g88 ( 
.A(n_79),
.Y(n_88)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_85),
.Y(n_105)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_99),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_100),
.A2(n_81),
.B1(n_73),
.B2(n_74),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_83),
.Y(n_101)
);

FAx1_ASAP7_75t_SL g121 ( 
.A(n_101),
.B(n_77),
.CI(n_75),
.CON(n_121),
.SN(n_121)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_109),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_105),
.B(n_110),
.Y(n_130)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_90),
.A2(n_88),
.B(n_79),
.Y(n_107)
);

AOI32xp33_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_112),
.A3(n_93),
.B1(n_104),
.B2(n_108),
.Y(n_120)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_80),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

INVx3_ASAP7_75t_SL g117 ( 
.A(n_111),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_79),
.B(n_68),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_112),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_113),
.B(n_118),
.Y(n_145)
);

MAJx2_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_77),
.C(n_66),
.Y(n_114)
);

MAJx2_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_77),
.C(n_75),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_54),
.C(n_59),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_128),
.C(n_65),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_107),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_120),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_122),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_67),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_55),
.B1(n_82),
.B2(n_69),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_123),
.A2(n_125),
.B1(n_127),
.B2(n_66),
.Y(n_139)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_57),
.B1(n_53),
.B2(n_76),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_126),
.A2(n_72),
.B1(n_78),
.B2(n_71),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_62),
.B1(n_58),
.B2(n_60),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_105),
.B(n_51),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_103),
.Y(n_129)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_133),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_52),
.Y(n_152)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_139),
.A2(n_140),
.B1(n_144),
.B2(n_70),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_113),
.A2(n_61),
.B1(n_56),
.B2(n_70),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_115),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_141),
.Y(n_154)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_142),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_125),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_143),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_136),
.A2(n_122),
.B1(n_130),
.B2(n_114),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_146),
.A2(n_148),
.B1(n_141),
.B2(n_1),
.Y(n_159)
);

AOI322xp5_ASAP7_75t_L g149 ( 
.A1(n_136),
.A2(n_121),
.A3(n_21),
.B1(n_26),
.B2(n_32),
.C1(n_49),
.C2(n_47),
.Y(n_149)
);

OAI32xp33_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_152),
.A3(n_134),
.B1(n_137),
.B2(n_20),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_14),
.C(n_41),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_153),
.A2(n_38),
.B(n_16),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_157),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_147),
.A2(n_135),
.B(n_131),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_159),
.C(n_160),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_150),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_152),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_162),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_151),
.B(n_155),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_29),
.C(n_45),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_166),
.A2(n_17),
.B(n_13),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_133),
.B(n_31),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_40),
.C(n_39),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_33),
.B(n_2),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_0),
.B(n_3),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_153),
.B(n_154),
.Y(n_172)
);

AO21x1_ASAP7_75t_SL g173 ( 
.A1(n_172),
.A2(n_154),
.B(n_3),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_146),
.B1(n_4),
.B2(n_6),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_0),
.B(n_4),
.Y(n_175)
);


endmodule