module real_aes_598_n_382 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_382);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_382;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_577;
wire n_1004;
wire n_469;
wire n_987;
wire n_979;
wire n_759;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_666;
wire n_551;
wire n_884;
wire n_537;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_948;
wire n_399;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_816;
wire n_539;
wire n_400;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_994;
wire n_384;
wire n_744;
wire n_938;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_981;
wire n_791;
wire n_559;
wire n_466;
wire n_1049;
wire n_872;
wire n_636;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_1025;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_725;
wire n_455;
wire n_504;
wire n_960;
wire n_671;
wire n_973;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_722;
wire n_867;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_449;
wire n_417;
wire n_754;
wire n_607;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_947;
wire n_561;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1031;
wire n_1037;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_488;
wire n_501;
wire n_1041;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_954;
wire n_702;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_756;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_1028;
wire n_727;
wire n_1014;
wire n_397;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_845;
wire n_850;
wire n_1043;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_698;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_603;
wire n_854;
wire n_403;
wire n_1039;
wire n_424;
wire n_802;
wire n_868;
wire n_877;
wire n_574;
wire n_1024;
wire n_842;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_0), .A2(n_333), .B1(n_588), .B2(n_589), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_1), .A2(n_219), .B1(n_594), .B2(n_626), .Y(n_625) );
AOI22xp33_ASAP7_75t_SL g685 ( .A1(n_2), .A2(n_283), .B1(n_610), .B2(n_686), .Y(n_685) );
AOI22xp33_ASAP7_75t_SL g911 ( .A1(n_3), .A2(n_170), .B1(n_430), .B2(n_912), .Y(n_911) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_4), .A2(n_117), .B1(n_487), .B2(n_683), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_5), .A2(n_125), .B1(n_651), .B2(n_678), .Y(n_677) );
CKINVDCx20_ASAP7_75t_R g696 ( .A(n_6), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_7), .A2(n_79), .B1(n_503), .B2(n_642), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g889 ( .A1(n_8), .A2(n_198), .B1(n_499), .B2(n_890), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_9), .B(n_576), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_10), .A2(n_345), .B1(n_646), .B2(n_666), .Y(n_1060) );
AOI22xp33_ASAP7_75t_SL g800 ( .A1(n_11), .A2(n_254), .B1(n_588), .B2(n_589), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g1036 ( .A1(n_12), .A2(n_92), .B1(n_535), .B2(n_580), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_13), .A2(n_190), .B1(n_895), .B2(n_896), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_14), .A2(n_289), .B1(n_666), .B2(n_754), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_15), .A2(n_205), .B1(n_596), .B2(n_597), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_16), .A2(n_239), .B1(n_1042), .B2(n_1044), .Y(n_1041) );
AOI22xp33_ASAP7_75t_SL g729 ( .A1(n_17), .A2(n_78), .B1(n_583), .B2(n_584), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_18), .A2(n_142), .B1(n_426), .B2(n_611), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_19), .A2(n_195), .B1(n_526), .B2(n_683), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_20), .A2(n_244), .B1(n_483), .B2(n_486), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_21), .A2(n_220), .B1(n_581), .B2(n_705), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_22), .A2(n_185), .B1(n_559), .B2(n_674), .Y(n_864) );
AOI22xp33_ASAP7_75t_SL g803 ( .A1(n_23), .A2(n_183), .B1(n_594), .B2(n_712), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_24), .A2(n_153), .B1(n_614), .B2(n_839), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_25), .A2(n_285), .B1(n_563), .B2(n_671), .Y(n_1057) );
XOR2x2_ASAP7_75t_L g807 ( .A(n_26), .B(n_808), .Y(n_807) );
AO222x2_ASAP7_75t_L g699 ( .A1(n_27), .A2(n_148), .B1(n_240), .B2(n_397), .C1(n_417), .C2(n_700), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_28), .A2(n_340), .B1(n_705), .B2(n_706), .Y(n_704) );
INVx1_ASAP7_75t_SL g402 ( .A(n_29), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g1021 ( .A(n_29), .B(n_40), .Y(n_1021) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_30), .Y(n_725) );
OA22x2_ASAP7_75t_L g978 ( .A1(n_31), .A2(n_979), .B1(n_980), .B2(n_981), .Y(n_978) );
CKINVDCx20_ASAP7_75t_R g979 ( .A(n_31), .Y(n_979) );
AOI22xp5_ASAP7_75t_L g844 ( .A1(n_32), .A2(n_179), .B1(n_667), .B2(n_753), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_33), .A2(n_378), .B1(n_678), .B2(n_818), .Y(n_972) );
AOI22xp33_ASAP7_75t_SL g425 ( .A1(n_34), .A2(n_137), .B1(n_426), .B2(n_430), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_35), .A2(n_85), .B1(n_487), .B2(n_1007), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_36), .A2(n_298), .B1(n_596), .B2(n_597), .Y(n_595) );
AOI22x1_ASAP7_75t_L g736 ( .A1(n_37), .A2(n_200), .B1(n_454), .B2(n_596), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_38), .A2(n_116), .B1(n_705), .B2(n_706), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_39), .A2(n_368), .B1(n_839), .B2(n_990), .Y(n_989) );
AO22x2_ASAP7_75t_L g404 ( .A1(n_40), .A2(n_359), .B1(n_401), .B2(n_405), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_41), .A2(n_178), .B1(n_466), .B2(n_469), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_42), .A2(n_214), .B1(n_754), .B2(n_816), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_43), .A2(n_54), .B1(n_610), .B2(n_686), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g986 ( .A1(n_44), .A2(n_113), .B1(n_678), .B2(n_758), .Y(n_986) );
AOI22xp5_ASAP7_75t_L g924 ( .A1(n_45), .A2(n_332), .B1(n_754), .B2(n_816), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_46), .A2(n_367), .B1(n_751), .B2(n_818), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_47), .A2(n_154), .B1(n_494), .B2(n_496), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_48), .A2(n_234), .B1(n_610), .B2(n_686), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_49), .A2(n_290), .B1(n_462), .B2(n_751), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_50), .A2(n_344), .B1(n_446), .B2(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g403 ( .A(n_51), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_52), .A2(n_245), .B1(n_667), .B2(n_751), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g804 ( .A1(n_53), .A2(n_314), .B1(n_593), .B2(n_597), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_55), .A2(n_236), .B1(n_498), .B2(n_500), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_56), .A2(n_310), .B1(n_596), .B2(n_711), .Y(n_801) );
AOI22xp33_ASAP7_75t_SL g920 ( .A1(n_57), .A2(n_318), .B1(n_751), .B2(n_921), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_58), .A2(n_132), .B1(n_823), .B2(n_824), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_59), .A2(n_356), .B1(n_459), .B2(n_619), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g932 ( .A1(n_60), .A2(n_249), .B1(n_683), .B2(n_933), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_61), .A2(n_355), .B1(n_758), .B2(n_926), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_62), .A2(n_216), .B1(n_896), .B2(n_926), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_63), .A2(n_348), .B1(n_446), .B2(n_449), .Y(n_970) );
AO22x2_ASAP7_75t_L g411 ( .A1(n_64), .A2(n_196), .B1(n_401), .B2(n_412), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_65), .A2(n_315), .B1(n_674), .B2(n_754), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_66), .A2(n_202), .B1(n_551), .B2(n_674), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g1048 ( .A1(n_67), .A2(n_82), .B1(n_551), .B2(n_1049), .Y(n_1048) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_68), .A2(n_238), .B1(n_446), .B2(n_500), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_69), .A2(n_107), .B1(n_415), .B2(n_421), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_70), .A2(n_165), .B1(n_583), .B2(n_584), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_71), .A2(n_297), .B1(n_452), .B2(n_651), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_72), .A2(n_328), .B1(n_452), .B2(n_454), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_73), .A2(n_171), .B1(n_597), .B2(n_711), .Y(n_737) );
AOI22xp5_ASAP7_75t_L g942 ( .A1(n_74), .A2(n_204), .B1(n_496), .B2(n_751), .Y(n_942) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_75), .A2(n_159), .B1(n_454), .B2(n_466), .Y(n_590) );
AOI22xp33_ASAP7_75t_SL g709 ( .A1(n_76), .A2(n_114), .B1(n_588), .B2(n_589), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_77), .A2(n_294), .B1(n_711), .B2(n_712), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_80), .A2(n_255), .B1(n_538), .B2(n_540), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_81), .A2(n_253), .B1(n_417), .B2(n_421), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_83), .A2(n_100), .B1(n_459), .B2(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_84), .B(n_607), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_86), .A2(n_370), .B1(n_487), .B2(n_683), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_87), .A2(n_227), .B1(n_449), .B2(n_648), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g1005 ( .A1(n_88), .A2(n_308), .B1(n_540), .B2(n_990), .Y(n_1005) );
AOI22xp5_ASAP7_75t_L g842 ( .A1(n_89), .A2(n_286), .B1(n_756), .B2(n_843), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_90), .A2(n_139), .B1(n_556), .B2(n_946), .Y(n_945) );
AO222x2_ASAP7_75t_L g794 ( .A1(n_91), .A2(n_213), .B1(n_362), .B2(n_397), .C1(n_581), .C2(n_584), .Y(n_794) );
AOI22xp33_ASAP7_75t_SL g668 ( .A1(n_93), .A2(n_127), .B1(n_669), .B2(n_671), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_94), .A2(n_231), .B1(n_580), .B2(n_581), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g875 ( .A1(n_95), .A2(n_235), .B1(n_604), .B2(n_747), .Y(n_875) );
AOI22xp33_ASAP7_75t_SL g797 ( .A1(n_96), .A2(n_258), .B1(n_417), .B2(n_421), .Y(n_797) );
CKINVDCx20_ASAP7_75t_R g560 ( .A(n_97), .Y(n_560) );
AOI222xp33_ASAP7_75t_L g1006 ( .A1(n_98), .A2(n_180), .B1(n_347), .B2(n_487), .C1(n_745), .C2(n_1007), .Y(n_1006) );
OA22x2_ASAP7_75t_L g514 ( .A1(n_99), .A2(n_515), .B1(n_516), .B2(n_517), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_99), .Y(n_515) );
AOI222xp33_ASAP7_75t_L g744 ( .A1(n_101), .A2(n_145), .B1(n_282), .B2(n_614), .C1(n_689), .C2(n_745), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_102), .A2(n_160), .B1(n_584), .B2(n_703), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g1037 ( .A1(n_103), .A2(n_277), .B1(n_1038), .B2(n_1039), .Y(n_1037) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_104), .A2(n_237), .B1(n_823), .B2(n_824), .Y(n_1045) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_105), .A2(n_197), .B1(n_644), .B2(n_646), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_106), .A2(n_126), .B1(n_506), .B2(n_821), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_108), .A2(n_339), .B1(n_459), .B2(n_462), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_109), .B(n_476), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_110), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_111), .A2(n_241), .B1(n_446), .B2(n_449), .Y(n_985) );
AO22x2_ASAP7_75t_L g408 ( .A1(n_112), .A2(n_293), .B1(n_401), .B2(n_409), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_115), .A2(n_306), .B1(n_688), .B2(n_839), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_118), .A2(n_157), .B1(n_688), .B2(n_689), .Y(n_687) );
AO21x2_ASAP7_75t_L g636 ( .A1(n_119), .A2(n_637), .B(n_657), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_119), .B(n_639), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_120), .A2(n_122), .B1(n_525), .B2(n_528), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_121), .A2(n_272), .B1(n_651), .B2(n_678), .Y(n_863) );
AOI22xp5_ASAP7_75t_L g973 ( .A1(n_123), .A2(n_147), .B1(n_666), .B2(n_667), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_124), .A2(n_270), .B1(n_490), .B2(n_491), .Y(n_489) );
INVx1_ASAP7_75t_L g1008 ( .A(n_128), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_129), .A2(n_354), .B1(n_589), .B2(n_771), .Y(n_770) );
OA22x2_ASAP7_75t_L g869 ( .A1(n_130), .A2(n_870), .B1(n_871), .B2(n_872), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_130), .Y(n_870) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_131), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_133), .A2(n_207), .B1(n_594), .B2(n_626), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_134), .A2(n_337), .B1(n_525), .B2(n_528), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_135), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_136), .B(n_477), .Y(n_958) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_138), .A2(n_230), .B1(n_426), .B2(n_686), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_140), .A2(n_177), .B1(n_495), .B2(n_893), .Y(n_892) );
CKINVDCx20_ASAP7_75t_R g598 ( .A(n_141), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_143), .A2(n_276), .B1(n_487), .B2(n_683), .Y(n_917) );
OA22x2_ASAP7_75t_L g471 ( .A1(n_144), .A2(n_472), .B1(n_473), .B2(n_508), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_144), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g815 ( .A1(n_146), .A2(n_330), .B1(n_667), .B2(n_816), .Y(n_815) );
AOI22xp5_ASAP7_75t_L g938 ( .A1(n_149), .A2(n_175), .B1(n_614), .B2(n_689), .Y(n_938) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_150), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_151), .A2(n_158), .B1(n_711), .B2(n_712), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g934 ( .A1(n_152), .A2(n_336), .B1(n_430), .B2(n_912), .Y(n_934) );
CKINVDCx20_ASAP7_75t_R g878 ( .A(n_155), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_156), .A2(n_181), .B1(n_538), .B2(n_540), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g888 ( .A1(n_161), .A2(n_377), .B1(n_496), .B2(n_645), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_162), .B(n_607), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g983 ( .A1(n_163), .A2(n_242), .B1(n_666), .B2(n_921), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_164), .A2(n_295), .B1(n_449), .B2(n_499), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_166), .A2(n_265), .B1(n_551), .B2(n_1049), .Y(n_1058) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_167), .B(n_521), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_168), .A2(n_189), .B1(n_452), .B2(n_506), .Y(n_505) );
AOI22xp33_ASAP7_75t_SL g445 ( .A1(n_169), .A2(n_327), .B1(n_446), .B2(n_448), .Y(n_445) );
AOI22xp33_ASAP7_75t_SL g922 ( .A1(n_172), .A2(n_307), .B1(n_446), .B2(n_500), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_173), .A2(n_349), .B1(n_481), .B2(n_614), .Y(n_811) );
OA22x2_ASAP7_75t_L g739 ( .A1(n_174), .A2(n_740), .B1(n_741), .B2(n_742), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_174), .Y(n_740) );
INVx1_ASAP7_75t_L g905 ( .A(n_176), .Y(n_905) );
CKINVDCx20_ASAP7_75t_R g883 ( .A(n_182), .Y(n_883) );
AOI22xp33_ASAP7_75t_SL g991 ( .A1(n_184), .A2(n_229), .B1(n_426), .B2(n_686), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_186), .A2(n_211), .B1(n_430), .B2(n_610), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_187), .A2(n_303), .B1(n_532), .B2(n_535), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_188), .A2(n_259), .B1(n_610), .B2(n_686), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_191), .A2(n_366), .B1(n_487), .B2(n_683), .Y(n_812) );
CKINVDCx20_ASAP7_75t_R g880 ( .A(n_192), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_193), .A2(n_381), .B1(n_559), .B2(n_753), .Y(n_1047) );
AOI22xp33_ASAP7_75t_SL g673 ( .A1(n_194), .A2(n_316), .B1(n_674), .B2(n_675), .Y(n_673) );
INVx1_ASAP7_75t_L g1020 ( .A(n_196), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_199), .A2(n_228), .B1(n_596), .B2(n_597), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_201), .A2(n_260), .B1(n_588), .B2(n_589), .Y(n_733) );
XNOR2xp5_ASAP7_75t_L g720 ( .A(n_203), .B(n_721), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_206), .A2(n_360), .B1(n_610), .B2(n_611), .Y(n_609) );
INVx1_ASAP7_75t_L g681 ( .A(n_208), .Y(n_681) );
AOI22xp33_ASAP7_75t_SL g796 ( .A1(n_209), .A2(n_326), .B1(n_703), .B2(n_705), .Y(n_796) );
AO21x1_ASAP7_75t_L g1022 ( .A1(n_210), .A2(n_1023), .B(n_1030), .Y(n_1022) );
CKINVDCx20_ASAP7_75t_R g567 ( .A(n_212), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_215), .A2(n_273), .B1(n_683), .B2(n_747), .Y(n_988) );
XNOR2x1_ASAP7_75t_L g953 ( .A(n_217), .B(n_954), .Y(n_953) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_218), .A2(n_373), .B1(n_683), .B2(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g1029 ( .A(n_221), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_222), .A2(n_369), .B1(n_593), .B2(n_594), .Y(n_714) );
OA22x2_ASAP7_75t_L g928 ( .A1(n_223), .A2(n_929), .B1(n_947), .B2(n_948), .Y(n_928) );
CKINVDCx20_ASAP7_75t_R g947 ( .A(n_223), .Y(n_947) );
AOI22xp33_ASAP7_75t_SL g846 ( .A1(n_224), .A2(n_278), .B1(n_551), .B2(n_678), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g1059 ( .A1(n_225), .A2(n_311), .B1(n_674), .B2(n_1044), .Y(n_1059) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_226), .A2(n_246), .B1(n_469), .B2(n_926), .Y(n_1002) );
XOR2xp5_ASAP7_75t_L g1031 ( .A(n_232), .B(n_1032), .Y(n_1031) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_233), .A2(n_323), .B1(n_753), .B2(n_754), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_243), .A2(n_288), .B1(n_499), .B2(n_756), .Y(n_941) );
CKINVDCx16_ASAP7_75t_R g776 ( .A(n_247), .Y(n_776) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_248), .A2(n_661), .B1(n_662), .B2(n_690), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_248), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g790 ( .A1(n_250), .A2(n_791), .B1(n_792), .B2(n_805), .Y(n_790) );
INVx1_ASAP7_75t_L g805 ( .A(n_250), .Y(n_805) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_251), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_252), .A2(n_346), .B1(n_435), .B2(n_439), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_256), .A2(n_341), .B1(n_417), .B2(n_700), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_257), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g916 ( .A(n_261), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_262), .B(n_521), .Y(n_1065) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_263), .A2(n_274), .B1(n_487), .B2(n_683), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_264), .A2(n_324), .B1(n_435), .B2(n_481), .Y(n_480) );
AOI22xp33_ASAP7_75t_SL g702 ( .A1(n_266), .A2(n_291), .B1(n_584), .B2(n_703), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_267), .A2(n_380), .B1(n_594), .B2(n_626), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_268), .A2(n_353), .B1(n_624), .B2(n_751), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_269), .B(n_607), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_271), .A2(n_305), .B1(n_487), .B2(n_604), .Y(n_603) );
XNOR2x1_ASAP7_75t_L g829 ( .A(n_275), .B(n_830), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g960 ( .A(n_279), .Y(n_960) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_280), .A2(n_358), .B1(n_623), .B2(n_624), .Y(n_622) );
XNOR2x1_ASAP7_75t_L g1054 ( .A(n_281), .B(n_1055), .Y(n_1054) );
INVxp67_ASAP7_75t_L g1068 ( .A(n_281), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_284), .B(n_477), .Y(n_810) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_287), .Y(n_549) );
AOI22xp33_ASAP7_75t_SL g665 ( .A1(n_292), .A2(n_335), .B1(n_666), .B2(n_667), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g1018 ( .A(n_293), .B(n_1019), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_296), .A2(n_375), .B1(n_615), .B2(n_688), .Y(n_1063) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_299), .B(n_477), .Y(n_936) );
CKINVDCx20_ASAP7_75t_R g966 ( .A(n_300), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_301), .A2(n_379), .B1(n_446), .B2(n_448), .Y(n_862) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_302), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_304), .A2(n_338), .B1(n_532), .B2(n_535), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_309), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_312), .A2(n_334), .B1(n_678), .B2(n_758), .Y(n_757) );
INVx3_ASAP7_75t_L g401 ( .A(n_313), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_317), .A2(n_329), .B1(n_593), .B2(n_594), .Y(n_592) );
AOI222xp33_ASAP7_75t_L g1050 ( .A1(n_319), .A2(n_357), .B1(n_364), .B2(n_477), .C1(n_525), .C2(n_528), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_320), .A2(n_365), .B1(n_481), .B2(n_539), .Y(n_913) );
OAI22x1_ASAP7_75t_L g853 ( .A1(n_321), .A2(n_854), .B1(n_865), .B2(n_866), .Y(n_853) );
INVx1_ASAP7_75t_L g866 ( .A(n_321), .Y(n_866) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_322), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g965 ( .A(n_325), .Y(n_965) );
CKINVDCx20_ASAP7_75t_R g627 ( .A(n_331), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_342), .B(n_745), .Y(n_992) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_343), .Y(n_413) );
CKINVDCx20_ASAP7_75t_R g885 ( .A(n_350), .Y(n_885) );
INVx1_ASAP7_75t_L g392 ( .A(n_351), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_352), .A2(n_376), .B1(n_614), .B2(n_615), .Y(n_613) );
INVx1_ASAP7_75t_L g1015 ( .A(n_361), .Y(n_1015) );
NAND2xp5_ASAP7_75t_SL g1028 ( .A(n_361), .B(n_1029), .Y(n_1028) );
INVx1_ASAP7_75t_L g1016 ( .A(n_363), .Y(n_1016) );
AND2x2_ASAP7_75t_R g1052 ( .A(n_363), .B(n_1015), .Y(n_1052) );
INVxp67_ASAP7_75t_L g1027 ( .A(n_371), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_372), .B(n_397), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g962 ( .A(n_374), .Y(n_962) );
AOI21xp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_1011), .B(n_1022), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_781), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AOI21xp33_ASAP7_75t_L g1011 ( .A1(n_385), .A2(n_782), .B(n_1012), .Y(n_1011) );
AOI22xp33_ASAP7_75t_SL g385 ( .A1(n_386), .A2(n_632), .B1(n_633), .B2(n_780), .Y(n_385) );
INVx1_ASAP7_75t_SL g780 ( .A(n_386), .Y(n_780) );
OAI21x1_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_510), .B(n_631), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_387), .B(n_512), .Y(n_631) );
AO22x1_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_389), .B1(n_471), .B2(n_509), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
XNOR2x1_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
NAND2x1_ASAP7_75t_L g393 ( .A(n_394), .B(n_443), .Y(n_393) );
NOR2xp67_ASAP7_75t_L g394 ( .A(n_395), .B(n_424), .Y(n_394) );
OAI21xp5_ASAP7_75t_SL g395 ( .A1(n_396), .A2(n_413), .B(n_414), .Y(n_395) );
OAI222xp33_ASAP7_75t_L g723 ( .A1(n_396), .A2(n_416), .B1(n_724), .B2(n_725), .C1(n_726), .C2(n_727), .Y(n_723) );
INVx2_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
AND2x4_ASAP7_75t_L g397 ( .A(n_398), .B(n_406), .Y(n_397) );
AND2x4_ASAP7_75t_L g431 ( .A(n_398), .B(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_L g441 ( .A(n_398), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g479 ( .A(n_398), .B(n_406), .Y(n_479) );
AND2x2_ASAP7_75t_L g581 ( .A(n_398), .B(n_432), .Y(n_581) );
AND2x2_ASAP7_75t_L g584 ( .A(n_398), .B(n_442), .Y(n_584) );
AND2x2_ASAP7_75t_L g706 ( .A(n_398), .B(n_432), .Y(n_706) );
AND2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_404), .Y(n_398) );
AND2x2_ASAP7_75t_L g419 ( .A(n_399), .B(n_420), .Y(n_419) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_399), .Y(n_422) );
INVx2_ASAP7_75t_L g438 ( .A(n_399), .Y(n_438) );
OAI22x1_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B1(n_402), .B2(n_403), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g405 ( .A(n_401), .Y(n_405) );
INVx2_ASAP7_75t_L g409 ( .A(n_401), .Y(n_409) );
INVx1_ASAP7_75t_L g412 ( .A(n_401), .Y(n_412) );
INVx2_ASAP7_75t_L g420 ( .A(n_404), .Y(n_420) );
AND2x2_ASAP7_75t_L g437 ( .A(n_404), .B(n_438), .Y(n_437) );
BUFx2_ASAP7_75t_L g450 ( .A(n_404), .Y(n_450) );
AND2x4_ASAP7_75t_L g453 ( .A(n_406), .B(n_419), .Y(n_453) );
AND2x2_ASAP7_75t_L g461 ( .A(n_406), .B(n_437), .Y(n_461) );
AND2x4_ASAP7_75t_L g468 ( .A(n_406), .B(n_456), .Y(n_468) );
AND2x2_ASAP7_75t_L g593 ( .A(n_406), .B(n_419), .Y(n_593) );
AND2x6_ASAP7_75t_L g596 ( .A(n_406), .B(n_437), .Y(n_596) );
AND2x2_ASAP7_75t_L g626 ( .A(n_406), .B(n_419), .Y(n_626) );
AND2x2_ASAP7_75t_L g711 ( .A(n_406), .B(n_456), .Y(n_711) );
AND2x4_ASAP7_75t_L g406 ( .A(n_407), .B(n_410), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AND2x4_ASAP7_75t_L g418 ( .A(n_408), .B(n_410), .Y(n_418) );
AND2x2_ASAP7_75t_L g423 ( .A(n_408), .B(n_411), .Y(n_423) );
INVx1_ASAP7_75t_L g429 ( .A(n_408), .Y(n_429) );
INVxp67_ASAP7_75t_L g442 ( .A(n_410), .Y(n_442) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g428 ( .A(n_411), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
AND2x4_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
AND2x4_ASAP7_75t_L g436 ( .A(n_418), .B(n_437), .Y(n_436) );
AND2x4_ASAP7_75t_L g455 ( .A(n_418), .B(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g485 ( .A(n_418), .B(n_419), .Y(n_485) );
AND2x2_ASAP7_75t_L g583 ( .A(n_418), .B(n_437), .Y(n_583) );
AND2x2_ASAP7_75t_L g703 ( .A(n_418), .B(n_437), .Y(n_703) );
AND2x2_ASAP7_75t_L g712 ( .A(n_418), .B(n_456), .Y(n_712) );
AND2x2_ASAP7_75t_L g427 ( .A(n_419), .B(n_428), .Y(n_427) );
AND2x4_ASAP7_75t_L g705 ( .A(n_419), .B(n_428), .Y(n_705) );
AND2x4_ASAP7_75t_L g456 ( .A(n_420), .B(n_438), .Y(n_456) );
INVxp67_ASAP7_75t_L g727 ( .A(n_421), .Y(n_727) );
AND2x2_ASAP7_75t_SL g421 ( .A(n_422), .B(n_423), .Y(n_421) );
AND2x2_ASAP7_75t_L g488 ( .A(n_422), .B(n_423), .Y(n_488) );
AND2x2_ASAP7_75t_SL g700 ( .A(n_422), .B(n_423), .Y(n_700) );
AND2x4_ASAP7_75t_L g449 ( .A(n_423), .B(n_450), .Y(n_449) );
AND2x4_ASAP7_75t_L g470 ( .A(n_423), .B(n_456), .Y(n_470) );
AND2x4_ASAP7_75t_L g589 ( .A(n_423), .B(n_450), .Y(n_589) );
AND2x4_ASAP7_75t_L g594 ( .A(n_423), .B(n_456), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_425), .B(n_434), .Y(n_424) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_426), .Y(n_490) );
INVx1_ASAP7_75t_L g879 ( .A(n_426), .Y(n_879) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx3_ASAP7_75t_L g534 ( .A(n_427), .Y(n_534) );
BUFx6f_ASAP7_75t_L g610 ( .A(n_427), .Y(n_610) );
AND2x2_ASAP7_75t_L g447 ( .A(n_428), .B(n_437), .Y(n_447) );
AND2x4_ASAP7_75t_L g464 ( .A(n_428), .B(n_456), .Y(n_464) );
AND2x2_ASAP7_75t_SL g588 ( .A(n_428), .B(n_437), .Y(n_588) );
AND2x6_ASAP7_75t_L g597 ( .A(n_428), .B(n_456), .Y(n_597) );
AND2x2_ASAP7_75t_L g771 ( .A(n_428), .B(n_437), .Y(n_771) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_429), .Y(n_433) );
BUFx2_ASAP7_75t_SL g491 ( .A(n_430), .Y(n_491) );
INVxp67_ASAP7_75t_L g881 ( .A(n_430), .Y(n_881) );
BUFx6f_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
BUFx3_ASAP7_75t_L g536 ( .A(n_431), .Y(n_536) );
INVx2_ASAP7_75t_L g612 ( .A(n_431), .Y(n_612) );
BUFx4f_ASAP7_75t_L g686 ( .A(n_431), .Y(n_686) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_436), .Y(n_539) );
BUFx3_ASAP7_75t_L g614 ( .A(n_436), .Y(n_614) );
BUFx2_ASAP7_75t_L g990 ( .A(n_436), .Y(n_990) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g481 ( .A(n_440), .Y(n_481) );
INVx2_ASAP7_75t_L g540 ( .A(n_440), .Y(n_540) );
INVx2_ASAP7_75t_L g615 ( .A(n_440), .Y(n_615) );
INVx2_ASAP7_75t_SL g689 ( .A(n_440), .Y(n_689) );
INVx2_ASAP7_75t_SL g839 ( .A(n_440), .Y(n_839) );
OAI22xp5_ASAP7_75t_L g882 ( .A1(n_440), .A2(n_883), .B1(n_884), .B2(n_885), .Y(n_882) );
OAI22xp5_ASAP7_75t_L g964 ( .A1(n_440), .A2(n_884), .B1(n_965), .B2(n_966), .Y(n_964) );
INVx2_ASAP7_75t_L g1039 ( .A(n_440), .Y(n_1039) );
INVx6_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_457), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_451), .Y(n_444) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx3_ASAP7_75t_L g499 ( .A(n_447), .Y(n_499) );
INVx2_ASAP7_75t_L g566 ( .A(n_447), .Y(n_566) );
BUFx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx5_ASAP7_75t_SL g501 ( .A(n_449), .Y(n_501) );
BUFx2_ASAP7_75t_L g824 ( .A(n_449), .Y(n_824) );
BUFx3_ASAP7_75t_L g890 ( .A(n_449), .Y(n_890) );
BUFx3_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx6_ASAP7_75t_L g544 ( .A(n_453), .Y(n_544) );
BUFx3_ASAP7_75t_L g895 ( .A(n_453), .Y(n_895) );
INVx2_ASAP7_75t_L g504 ( .A(n_454), .Y(n_504) );
BUFx6f_ASAP7_75t_L g1044 ( .A(n_454), .Y(n_1044) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_455), .Y(n_624) );
INVx2_ASAP7_75t_L g676 ( .A(n_455), .Y(n_676) );
BUFx3_ASAP7_75t_L g754 ( .A(n_455), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_465), .Y(n_457) );
INVx3_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g556 ( .A(n_460), .Y(n_556) );
INVx2_ASAP7_75t_SL g666 ( .A(n_460), .Y(n_666) );
INVx2_ASAP7_75t_SL g753 ( .A(n_460), .Y(n_753) );
INVx2_ASAP7_75t_L g816 ( .A(n_460), .Y(n_816) );
INVx3_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx2_ASAP7_75t_L g645 ( .A(n_461), .Y(n_645) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g496 ( .A(n_463), .Y(n_496) );
INVx2_ASAP7_75t_L g559 ( .A(n_463), .Y(n_559) );
INVx2_ASAP7_75t_SL g619 ( .A(n_463), .Y(n_619) );
INVx2_ASAP7_75t_L g646 ( .A(n_463), .Y(n_646) );
INVx2_ASAP7_75t_SL g667 ( .A(n_463), .Y(n_667) );
INVx1_ASAP7_75t_SL g921 ( .A(n_463), .Y(n_921) );
INVx8_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx3_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_SL g495 ( .A(n_467), .Y(n_495) );
INVx2_ASAP7_75t_L g623 ( .A(n_467), .Y(n_623) );
INVx4_ASAP7_75t_L g642 ( .A(n_467), .Y(n_642) );
INVx2_ASAP7_75t_SL g751 ( .A(n_467), .Y(n_751) );
INVx8_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g507 ( .A(n_470), .Y(n_507) );
BUFx2_ASAP7_75t_SL g551 ( .A(n_470), .Y(n_551) );
BUFx2_ASAP7_75t_SL g651 ( .A(n_470), .Y(n_651) );
BUFx3_ASAP7_75t_L g896 ( .A(n_470), .Y(n_896) );
INVx1_ASAP7_75t_L g509 ( .A(n_471), .Y(n_509) );
INVx1_ASAP7_75t_L g508 ( .A(n_473), .Y(n_508) );
OR2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_492), .Y(n_473) );
NAND4xp25_ASAP7_75t_SL g474 ( .A(n_475), .B(n_480), .C(n_482), .D(n_489), .Y(n_474) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx3_ASAP7_75t_SL g522 ( .A(n_478), .Y(n_522) );
INVx4_ASAP7_75t_SL g576 ( .A(n_478), .Y(n_576) );
INVx3_ASAP7_75t_L g607 ( .A(n_478), .Y(n_607) );
INVx4_ASAP7_75t_SL g745 ( .A(n_478), .Y(n_745) );
INVx6_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx3_ASAP7_75t_L g529 ( .A(n_485), .Y(n_529) );
INVx2_ASAP7_75t_L g605 ( .A(n_485), .Y(n_605) );
BUFx5_ASAP7_75t_L g683 ( .A(n_485), .Y(n_683) );
BUFx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx12f_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx3_ASAP7_75t_L g527 ( .A(n_488), .Y(n_527) );
NAND4xp25_ASAP7_75t_L g492 ( .A(n_493), .B(n_497), .C(n_502), .D(n_505), .Y(n_492) );
INVx1_ASAP7_75t_L g548 ( .A(n_494), .Y(n_548) );
BUFx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
OAI22xp33_ASAP7_75t_SL g561 ( .A1(n_501), .A2(n_562), .B1(n_567), .B2(n_568), .Y(n_561) );
INVx2_ASAP7_75t_L g671 ( .A(n_501), .Y(n_671) );
INVx3_ASAP7_75t_L g756 ( .A(n_501), .Y(n_756) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
OAI22xp33_ASAP7_75t_L g542 ( .A1(n_504), .A2(n_543), .B1(n_544), .B2(n_545), .Y(n_542) );
INVx2_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_SL g758 ( .A(n_507), .Y(n_758) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
OAI22x1_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_569), .B1(n_570), .B2(n_630), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g630 ( .A(n_514), .Y(n_630) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND3x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_541), .C(n_552), .Y(n_517) );
NOR2xp67_ASAP7_75t_SL g518 ( .A(n_519), .B(n_530), .Y(n_518) );
OAI21xp5_ASAP7_75t_SL g519 ( .A1(n_520), .A2(n_523), .B(n_524), .Y(n_519) );
OAI21xp33_ASAP7_75t_L g680 ( .A1(n_520), .A2(n_681), .B(n_682), .Y(n_680) );
INVx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
BUFx6f_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g747 ( .A(n_527), .Y(n_747) );
INVx2_ASAP7_75t_L g933 ( .A(n_527), .Y(n_933) );
BUFx6f_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_531), .B(n_537), .Y(n_530) );
BUFx3_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx4_ASAP7_75t_L g580 ( .A(n_534), .Y(n_580) );
INVx2_ASAP7_75t_L g912 ( .A(n_534), .Y(n_912) );
BUFx6f_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
BUFx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx4f_ASAP7_75t_SL g688 ( .A(n_539), .Y(n_688) );
INVx1_ASAP7_75t_L g884 ( .A(n_539), .Y(n_884) );
BUFx2_ASAP7_75t_L g1038 ( .A(n_539), .Y(n_1038) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_546), .Y(n_541) );
INVx2_ASAP7_75t_L g678 ( .A(n_544), .Y(n_678) );
INVx3_ASAP7_75t_L g821 ( .A(n_544), .Y(n_821) );
INVx2_ASAP7_75t_L g926 ( .A(n_544), .Y(n_926) );
INVx2_ASAP7_75t_L g1049 ( .A(n_544), .Y(n_1049) );
OAI22xp33_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B1(n_549), .B2(n_550), .Y(n_546) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_553), .B(n_561), .Y(n_552) );
OAI22xp33_ASAP7_75t_SL g553 ( .A1(n_554), .A2(n_557), .B1(n_558), .B2(n_560), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
BUFx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g843 ( .A(n_564), .Y(n_843) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g670 ( .A(n_565), .Y(n_670) );
BUFx6f_ASAP7_75t_L g823 ( .A(n_565), .Y(n_823) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g649 ( .A(n_566), .Y(n_649) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AO22x2_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_599), .B1(n_628), .B2(n_629), .Y(n_570) );
INVx1_ASAP7_75t_SL g629 ( .A(n_571), .Y(n_629) );
XOR2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_598), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_573), .B(n_585), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_578), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
INVx1_ASAP7_75t_SL g915 ( .A(n_576), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_582), .Y(n_578) );
INVx2_ASAP7_75t_SL g961 ( .A(n_580), .Y(n_961) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_586), .B(n_591), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_590), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_595), .Y(n_591) );
INVx2_ASAP7_75t_L g628 ( .A(n_599), .Y(n_628) );
XOR2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_627), .Y(n_599) );
NAND2x1p5_ASAP7_75t_L g600 ( .A(n_601), .B(n_616), .Y(n_600) );
NOR2x1_ASAP7_75t_L g601 ( .A(n_602), .B(n_608), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_606), .Y(n_602) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g1007 ( .A(n_605), .Y(n_1007) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_613), .Y(n_608) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NOR2x1_ASAP7_75t_L g616 ( .A(n_617), .B(n_621), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_625), .Y(n_621) );
INVx1_ASAP7_75t_L g819 ( .A(n_624), .Y(n_819) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
XNOR2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_692), .Y(n_633) );
AO22x1_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_636), .B1(n_658), .B2(n_691), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_640), .B(n_652), .Y(n_639) );
NAND4xp25_ASAP7_75t_SL g640 ( .A(n_641), .B(n_643), .C(n_647), .D(n_650), .Y(n_640) );
BUFx6f_ASAP7_75t_L g674 ( .A(n_642), .Y(n_674) );
INVx2_ASAP7_75t_L g1043 ( .A(n_642), .Y(n_1043) );
BUFx3_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND4xp25_ASAP7_75t_SL g652 ( .A(n_653), .B(n_654), .C(n_655), .D(n_656), .Y(n_652) );
INVx2_ASAP7_75t_L g691 ( .A(n_658), .Y(n_691) );
BUFx3_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVxp33_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g690 ( .A(n_662), .Y(n_690) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_679), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_672), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_668), .Y(n_664) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_677), .Y(n_672) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g893 ( .A(n_676), .Y(n_893) );
INVx2_ASAP7_75t_L g946 ( .A(n_676), .Y(n_946) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_680), .B(n_684), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_687), .Y(n_684) );
INVxp67_ASAP7_75t_L g963 ( .A(n_686), .Y(n_963) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_716), .B1(n_778), .B2(n_779), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
HB1xp67_ASAP7_75t_L g778 ( .A(n_694), .Y(n_778) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
XNOR2x1_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
AND2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_707), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_699), .B(n_701), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_704), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_713), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
INVx1_ASAP7_75t_L g779 ( .A(n_716), .Y(n_779) );
OAI22x1_ASAP7_75t_SL g716 ( .A1(n_717), .A2(n_718), .B1(n_738), .B2(n_777), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NAND2x1p5_ASAP7_75t_L g721 ( .A(n_722), .B(n_731), .Y(n_721) );
NOR2x1_ASAP7_75t_L g722 ( .A(n_723), .B(n_728), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
NOR2x1_ASAP7_75t_L g731 ( .A(n_732), .B(n_735), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
INVx2_ASAP7_75t_L g777 ( .A(n_738), .Y(n_777) );
XNOR2x1_ASAP7_75t_L g738 ( .A(n_739), .B(n_759), .Y(n_738) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
NOR2x1_ASAP7_75t_L g742 ( .A(n_743), .B(n_749), .Y(n_742) );
NAND3xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_746), .C(n_748), .Y(n_743) );
INVx1_ASAP7_75t_L g833 ( .A(n_745), .Y(n_833) );
NAND4xp25_ASAP7_75t_L g749 ( .A(n_750), .B(n_752), .C(n_755), .D(n_757), .Y(n_749) );
AO22x2_ASAP7_75t_L g868 ( .A1(n_759), .A2(n_869), .B1(n_897), .B2(n_898), .Y(n_868) );
INVx1_ASAP7_75t_L g898 ( .A(n_759), .Y(n_898) );
XOR2x2_ASAP7_75t_L g759 ( .A(n_760), .B(n_776), .Y(n_759) );
NAND2x1p5_ASAP7_75t_L g760 ( .A(n_761), .B(n_768), .Y(n_760) );
NOR2x1_ASAP7_75t_L g761 ( .A(n_762), .B(n_765), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
NOR2x1_ASAP7_75t_L g768 ( .A(n_769), .B(n_773), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_772), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_774), .B(n_775), .Y(n_773) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
XOR2xp5_ASAP7_75t_L g782 ( .A(n_783), .B(n_901), .Y(n_782) );
AOI22xp5_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_785), .B1(n_849), .B2(n_900), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
OAI22xp5_ASAP7_75t_SL g786 ( .A1(n_787), .A2(n_788), .B1(n_826), .B2(n_848), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
AO22x2_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_806), .B1(n_807), .B2(n_825), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
BUFx2_ASAP7_75t_L g825 ( .A(n_790), .Y(n_825) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
NAND2xp5_ASAP7_75t_SL g792 ( .A(n_793), .B(n_798), .Y(n_792) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .Y(n_795) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_799), .B(n_802), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_800), .B(n_801), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_803), .B(n_804), .Y(n_802) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
NOR2xp67_ASAP7_75t_L g808 ( .A(n_809), .B(n_814), .Y(n_808) );
NAND4xp25_ASAP7_75t_SL g809 ( .A(n_810), .B(n_811), .C(n_812), .D(n_813), .Y(n_809) );
NAND4xp25_ASAP7_75t_L g814 ( .A(n_815), .B(n_817), .C(n_820), .D(n_822), .Y(n_814) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g848 ( .A(n_828), .Y(n_848) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
AND2x4_ASAP7_75t_L g830 ( .A(n_831), .B(n_840), .Y(n_830) );
NOR2xp67_ASAP7_75t_L g831 ( .A(n_832), .B(n_836), .Y(n_831) );
OAI21xp5_ASAP7_75t_SL g832 ( .A1(n_833), .A2(n_834), .B(n_835), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_837), .B(n_838), .Y(n_836) );
NOR2x1_ASAP7_75t_L g840 ( .A(n_841), .B(n_845), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_842), .B(n_844), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_846), .B(n_847), .Y(n_845) );
INVx1_ASAP7_75t_L g900 ( .A(n_849), .Y(n_900) );
AOI22xp5_ASAP7_75t_L g849 ( .A1(n_850), .A2(n_851), .B1(n_867), .B2(n_899), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
HB1xp67_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g865 ( .A(n_854), .Y(n_865) );
OR2x2_ASAP7_75t_L g854 ( .A(n_855), .B(n_860), .Y(n_854) );
NAND4xp25_ASAP7_75t_L g855 ( .A(n_856), .B(n_857), .C(n_858), .D(n_859), .Y(n_855) );
NAND4xp25_ASAP7_75t_L g860 ( .A(n_861), .B(n_862), .C(n_863), .D(n_864), .Y(n_860) );
INVx1_ASAP7_75t_L g899 ( .A(n_867), .Y(n_899) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx1_ASAP7_75t_L g897 ( .A(n_869), .Y(n_897) );
INVx2_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
AND2x2_ASAP7_75t_L g872 ( .A(n_873), .B(n_886), .Y(n_872) );
NOR3xp33_ASAP7_75t_L g873 ( .A(n_874), .B(n_877), .C(n_882), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_875), .B(n_876), .Y(n_874) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_878), .A2(n_879), .B1(n_880), .B2(n_881), .Y(n_877) );
NOR2xp33_ASAP7_75t_L g886 ( .A(n_887), .B(n_891), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_888), .B(n_889), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_892), .B(n_894), .Y(n_891) );
OAI22xp5_ASAP7_75t_L g901 ( .A1(n_902), .A2(n_975), .B1(n_1009), .B2(n_1010), .Y(n_901) );
INVx1_ASAP7_75t_L g1009 ( .A(n_902), .Y(n_1009) );
OAI22xp5_ASAP7_75t_SL g902 ( .A1(n_903), .A2(n_952), .B1(n_953), .B2(n_974), .Y(n_902) );
INVx1_ASAP7_75t_L g974 ( .A(n_903), .Y(n_974) );
AO22x2_ASAP7_75t_SL g903 ( .A1(n_904), .A2(n_928), .B1(n_950), .B2(n_951), .Y(n_903) );
INVx2_ASAP7_75t_L g950 ( .A(n_904), .Y(n_950) );
OAI21x1_ASAP7_75t_L g904 ( .A1(n_905), .A2(n_906), .B(n_927), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_905), .B(n_908), .Y(n_927) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_909), .B(n_918), .Y(n_908) );
NOR2xp33_ASAP7_75t_L g909 ( .A(n_910), .B(n_914), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_911), .B(n_913), .Y(n_910) );
OAI21xp33_ASAP7_75t_L g914 ( .A1(n_915), .A2(n_916), .B(n_917), .Y(n_914) );
NOR2xp33_ASAP7_75t_L g918 ( .A(n_919), .B(n_923), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_920), .B(n_922), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_924), .B(n_925), .Y(n_923) );
INVx2_ASAP7_75t_L g951 ( .A(n_928), .Y(n_951) );
AOI22xp5_ASAP7_75t_L g977 ( .A1(n_928), .A2(n_951), .B1(n_978), .B2(n_993), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_930), .B(n_939), .Y(n_929) );
NOR3xp33_ASAP7_75t_L g930 ( .A(n_931), .B(n_935), .C(n_937), .Y(n_930) );
NOR4xp25_ASAP7_75t_L g948 ( .A(n_931), .B(n_940), .C(n_943), .D(n_949), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_932), .B(n_934), .Y(n_931) );
INVxp67_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_936), .B(n_938), .Y(n_949) );
INVxp67_ASAP7_75t_SL g937 ( .A(n_938), .Y(n_937) );
NOR2xp33_ASAP7_75t_L g939 ( .A(n_940), .B(n_943), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_941), .B(n_942), .Y(n_940) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_944), .B(n_945), .Y(n_943) );
INVx1_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_955), .B(n_967), .Y(n_954) );
NOR3xp33_ASAP7_75t_L g955 ( .A(n_956), .B(n_959), .C(n_964), .Y(n_955) );
NAND2xp5_ASAP7_75t_SL g956 ( .A(n_957), .B(n_958), .Y(n_956) );
OAI22xp5_ASAP7_75t_L g959 ( .A1(n_960), .A2(n_961), .B1(n_962), .B2(n_963), .Y(n_959) );
NOR2xp33_ASAP7_75t_L g967 ( .A(n_968), .B(n_971), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g968 ( .A(n_969), .B(n_970), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_972), .B(n_973), .Y(n_971) );
INVx2_ASAP7_75t_SL g1010 ( .A(n_975), .Y(n_1010) );
OA22x2_ASAP7_75t_L g975 ( .A1(n_976), .A2(n_977), .B1(n_994), .B2(n_995), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
INVx1_ASAP7_75t_L g993 ( .A(n_978), .Y(n_993) );
INVx1_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
NOR2x1_ASAP7_75t_L g981 ( .A(n_982), .B(n_987), .Y(n_981) );
NAND4xp25_ASAP7_75t_L g982 ( .A(n_983), .B(n_984), .C(n_985), .D(n_986), .Y(n_982) );
NAND4xp25_ASAP7_75t_L g987 ( .A(n_988), .B(n_989), .C(n_991), .D(n_992), .Y(n_987) );
INVx3_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
XOR2x2_ASAP7_75t_L g995 ( .A(n_996), .B(n_1008), .Y(n_995) );
NAND4xp75_ASAP7_75t_L g996 ( .A(n_997), .B(n_1000), .C(n_1003), .D(n_1006), .Y(n_996) );
AND2x2_ASAP7_75t_L g997 ( .A(n_998), .B(n_999), .Y(n_997) );
AND2x2_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1002), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1005), .Y(n_1003) );
INVx1_ASAP7_75t_SL g1012 ( .A(n_1013), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1017), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1066 ( .A(n_1014), .B(n_1018), .Y(n_1066) );
NOR2xp33_ASAP7_75t_L g1014 ( .A(n_1015), .B(n_1016), .Y(n_1014) );
INVx1_ASAP7_75t_L g1025 ( .A(n_1016), .Y(n_1025) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
NAND2xp5_ASAP7_75t_L g1019 ( .A(n_1020), .B(n_1021), .Y(n_1019) );
AND2x4_ASAP7_75t_SL g1023 ( .A(n_1024), .B(n_1026), .Y(n_1023) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
OR2x2_ASAP7_75t_L g1067 ( .A(n_1025), .B(n_1026), .Y(n_1067) );
NOR2xp33_ASAP7_75t_L g1026 ( .A(n_1027), .B(n_1028), .Y(n_1026) );
OAI222xp33_ASAP7_75t_R g1030 ( .A1(n_1031), .A2(n_1051), .B1(n_1053), .B2(n_1066), .C1(n_1067), .C2(n_1068), .Y(n_1030) );
CKINVDCx14_ASAP7_75t_R g1032 ( .A(n_1033), .Y(n_1032) );
HB1xp67_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
NAND4xp75_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1040), .C(n_1046), .D(n_1050), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_1036), .B(n_1037), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1045), .Y(n_1040) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_1047), .B(n_1048), .Y(n_1046) );
INVx1_ASAP7_75t_SL g1051 ( .A(n_1052), .Y(n_1051) );
HB1xp67_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
OR2x2_ASAP7_75t_L g1055 ( .A(n_1056), .B(n_1061), .Y(n_1055) );
NAND4xp25_ASAP7_75t_L g1056 ( .A(n_1057), .B(n_1058), .C(n_1059), .D(n_1060), .Y(n_1056) );
NAND4xp25_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1063), .C(n_1064), .D(n_1065), .Y(n_1061) );
endmodule