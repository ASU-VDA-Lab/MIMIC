module fake_jpeg_13500_n_661 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_661);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_661;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_525;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_332;
wire n_92;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_442;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_7),
.B(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_11),
.B(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_14),
.B(n_10),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_11),
.Y(n_59)
);

INVx11_ASAP7_75t_SL g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_64),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_67),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_68),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_69),
.B(n_73),
.Y(n_138)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_70),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_71),
.Y(n_148)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_72),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_18),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_74),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_75),
.B(n_79),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_76),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_77),
.Y(n_182)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_78),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_21),
.B(n_17),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_80),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_21),
.B(n_17),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_81),
.B(n_83),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_85),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_86),
.Y(n_189)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_87),
.Y(n_216)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_88),
.Y(n_194)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_89),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_60),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_90),
.B(n_91),
.Y(n_177)
);

BUFx12f_ASAP7_75t_SL g91 ( 
.A(n_60),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_92),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_93),
.Y(n_176)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_29),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_96),
.B(n_107),
.Y(n_181)
);

INVx3_ASAP7_75t_SL g97 ( 
.A(n_27),
.Y(n_97)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_97),
.Y(n_195)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_98),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_99),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_100),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_101),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_20),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_20),
.Y(n_103)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_103),
.Y(n_170)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_34),
.Y(n_104)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_104),
.Y(n_153)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_105),
.Y(n_172)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_22),
.Y(n_106)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_106),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_29),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_24),
.B(n_29),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_108),
.B(n_111),
.Y(n_217)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_109),
.Y(n_200)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_110),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_24),
.B(n_16),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_20),
.Y(n_112)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_112),
.Y(n_168)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_19),
.Y(n_113)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_30),
.Y(n_114)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_36),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_115),
.B(n_128),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_34),
.Y(n_116)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_116),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_27),
.Y(n_117)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_117),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_23),
.B(n_16),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_123),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_27),
.Y(n_119)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_119),
.Y(n_192)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_28),
.Y(n_120)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_120),
.Y(n_205)
);

INVx2_ASAP7_75t_R g121 ( 
.A(n_36),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_41),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_28),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_23),
.B(n_0),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_20),
.Y(n_124)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_37),
.Y(n_125)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_125),
.Y(n_204)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_30),
.Y(n_126)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_127),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_35),
.B(n_0),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_28),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_55),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_130),
.B(n_37),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_139),
.B(n_214),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_80),
.A2(n_53),
.B1(n_56),
.B2(n_37),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_142),
.A2(n_86),
.B1(n_85),
.B2(n_77),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_121),
.B(n_59),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_149),
.B(n_166),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g157 ( 
.A(n_68),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_157),
.Y(n_274)
);

BUFx12_ASAP7_75t_L g159 ( 
.A(n_94),
.Y(n_159)
);

BUFx8_ASAP7_75t_L g225 ( 
.A(n_159),
.Y(n_225)
);

INVx11_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g252 ( 
.A(n_160),
.Y(n_252)
);

OAI21xp33_ASAP7_75t_L g161 ( 
.A1(n_91),
.A2(n_59),
.B(n_54),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_161),
.B(n_35),
.Y(n_235)
);

NAND2x1_ASAP7_75t_SL g294 ( 
.A(n_163),
.B(n_1),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_102),
.Y(n_166)
);

BUFx2_ASAP7_75t_SL g173 ( 
.A(n_125),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_173),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_66),
.B(n_54),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_175),
.B(n_186),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_97),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_180),
.B(n_188),
.Y(n_255)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_103),
.Y(n_184)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_184),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_89),
.B(n_46),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_109),
.Y(n_187)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_95),
.B(n_46),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_105),
.B(n_39),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_196),
.B(n_198),
.Y(n_268)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_110),
.Y(n_197)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_197),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_95),
.B(n_39),
.Y(n_198)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_117),
.Y(n_207)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_120),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_208),
.B(n_211),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_104),
.B(n_44),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_209),
.B(n_48),
.Y(n_283)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_119),
.Y(n_210)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_210),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_82),
.B(n_44),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_122),
.Y(n_212)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_212),
.Y(n_253)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_72),
.Y(n_213)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_213),
.Y(n_276)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_87),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g215 ( 
.A(n_93),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_215),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_135),
.A2(n_129),
.B1(n_116),
.B2(n_101),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_218),
.A2(n_279),
.B1(n_142),
.B2(n_183),
.Y(n_310)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_176),
.Y(n_220)
);

INVx6_ASAP7_75t_L g296 ( 
.A(n_220),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_174),
.A2(n_99),
.B1(n_100),
.B2(n_63),
.Y(n_222)
);

OAI21xp33_ASAP7_75t_SL g309 ( 
.A1(n_222),
.A2(n_240),
.B(n_294),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_181),
.B(n_43),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_223),
.B(n_238),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_136),
.B(n_43),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_224),
.B(n_260),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_177),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_226),
.B(n_231),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_141),
.A2(n_112),
.B1(n_56),
.B2(n_53),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_228),
.A2(n_134),
.B(n_154),
.Y(n_314)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_172),
.Y(n_229)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_229),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_177),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_230),
.B(n_258),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_133),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_234),
.A2(n_280),
.B1(n_286),
.B2(n_250),
.Y(n_340)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_235),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_131),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_237),
.Y(n_322)
);

AOI21xp33_ASAP7_75t_L g238 ( 
.A1(n_138),
.A2(n_41),
.B(n_57),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_194),
.A2(n_76),
.B1(n_65),
.B2(n_42),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_133),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_241),
.B(n_261),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_181),
.B(n_137),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_244),
.B(n_262),
.Y(n_301)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_145),
.Y(n_245)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_245),
.Y(n_295)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_156),
.Y(n_246)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_246),
.Y(n_337)
);

CKINVDCx12_ASAP7_75t_R g247 ( 
.A(n_132),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_247),
.Y(n_319)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_147),
.Y(n_248)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_248),
.Y(n_306)
);

OR2x4_ASAP7_75t_L g249 ( 
.A(n_161),
.B(n_37),
.Y(n_249)
);

NAND2xp33_ASAP7_75t_SL g326 ( 
.A(n_249),
.B(n_282),
.Y(n_326)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_176),
.Y(n_251)
);

INVx5_ASAP7_75t_L g316 ( 
.A(n_251),
.Y(n_316)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_206),
.Y(n_254)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_254),
.Y(n_339)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_195),
.Y(n_256)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_256),
.Y(n_347)
);

BUFx4f_ASAP7_75t_L g257 ( 
.A(n_190),
.Y(n_257)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_257),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_163),
.B(n_38),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_131),
.Y(n_259)
);

INVx5_ASAP7_75t_L g341 ( 
.A(n_259),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_138),
.B(n_38),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_187),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_158),
.B(n_57),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_158),
.B(n_51),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_263),
.B(n_275),
.Y(n_321)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_203),
.Y(n_264)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_264),
.Y(n_333)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_205),
.Y(n_265)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_265),
.Y(n_352)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_144),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_266),
.Y(n_304)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_169),
.Y(n_267)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_267),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_171),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_269),
.B(n_271),
.Y(n_330)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_183),
.Y(n_270)
);

INVx8_ASAP7_75t_L g312 ( 
.A(n_270),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_159),
.Y(n_271)
);

CKINVDCx12_ASAP7_75t_R g272 ( 
.A(n_173),
.Y(n_272)
);

BUFx8_ASAP7_75t_L g354 ( 
.A(n_272),
.Y(n_354)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_147),
.Y(n_273)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_273),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_165),
.B(n_51),
.Y(n_275)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_155),
.Y(n_277)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_277),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_199),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_278),
.B(n_284),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_162),
.A2(n_56),
.B1(n_53),
.B2(n_32),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_171),
.A2(n_50),
.B1(n_48),
.B2(n_45),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_162),
.Y(n_281)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_281),
.Y(n_355)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_217),
.B(n_50),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_283),
.B(n_290),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_165),
.B(n_45),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_217),
.B(n_42),
.Y(n_285)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_285),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_179),
.A2(n_32),
.B1(n_37),
.B2(n_6),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_202),
.B(n_150),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_287),
.B(n_200),
.Y(n_317)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_140),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_289),
.Y(n_298)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_155),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_170),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_291),
.Y(n_307)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_157),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_292),
.Y(n_353)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_168),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_293),
.B(n_148),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_287),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_302),
.B(n_305),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_224),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g363 ( 
.A1(n_310),
.A2(n_335),
.B1(n_185),
.B2(n_146),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_235),
.A2(n_190),
.B1(n_201),
.B2(n_191),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_311),
.A2(n_323),
.B1(n_329),
.B2(n_346),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_314),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_317),
.B(n_324),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_236),
.B(n_167),
.C(n_151),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_318),
.B(n_343),
.C(n_351),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_235),
.A2(n_201),
.B1(n_191),
.B2(n_143),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_219),
.B(n_204),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_218),
.A2(n_153),
.B1(n_193),
.B2(n_216),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_245),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_332),
.B(n_345),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_228),
.A2(n_249),
.B1(n_279),
.B2(n_282),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_260),
.B(n_152),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_336),
.B(n_267),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_340),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_342),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_246),
.B(n_200),
.C(n_216),
.Y(n_343)
);

OAI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_258),
.A2(n_265),
.B1(n_288),
.B2(n_294),
.Y(n_344)
);

OA22x2_ASAP7_75t_L g389 ( 
.A1(n_344),
.A2(n_348),
.B1(n_293),
.B2(n_264),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_227),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_268),
.A2(n_193),
.B1(n_164),
.B2(n_192),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_281),
.A2(n_164),
.B1(n_185),
.B2(n_182),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_232),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_349),
.B(n_295),
.Y(n_368)
);

FAx1_ASAP7_75t_SL g350 ( 
.A(n_255),
.B(n_1),
.CI(n_4),
.CON(n_350),
.SN(n_350)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_350),
.B(n_1),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_266),
.B(n_1),
.Y(n_351)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_350),
.B(n_221),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_357),
.B(n_364),
.Y(n_424)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_352),
.Y(n_359)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_359),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_326),
.A2(n_233),
.B(n_276),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_362),
.A2(n_380),
.B(n_327),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_363),
.A2(n_400),
.B1(n_297),
.B2(n_319),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_330),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_295),
.Y(n_365)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_365),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_366),
.B(n_367),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_300),
.B(n_243),
.Y(n_367)
);

CKINVDCx14_ASAP7_75t_R g410 ( 
.A(n_368),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_300),
.B(n_239),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_369),
.B(n_375),
.Y(n_422)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_352),
.Y(n_370)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_370),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_371),
.B(n_378),
.Y(n_441)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_337),
.Y(n_372)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_372),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_314),
.A2(n_250),
.B(n_269),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_373),
.A2(n_379),
.B(n_362),
.Y(n_425)
);

INVx8_ASAP7_75t_L g374 ( 
.A(n_322),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_374),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_317),
.B(n_253),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g377 ( 
.A1(n_310),
.A2(n_254),
.B1(n_229),
.B2(n_189),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g419 ( 
.A(n_377),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_301),
.B(n_233),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_326),
.A2(n_320),
.B(n_303),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_331),
.B(n_256),
.Y(n_381)
);

CKINVDCx14_ASAP7_75t_R g433 ( 
.A(n_381),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_329),
.A2(n_178),
.B1(n_189),
.B2(n_182),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_383),
.A2(n_398),
.B1(n_341),
.B2(n_237),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_336),
.B(n_318),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_384),
.B(n_396),
.Y(n_437)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_337),
.Y(n_385)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_385),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_321),
.B(n_291),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_386),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_324),
.B(n_289),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_387),
.Y(n_428)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_347),
.Y(n_388)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_388),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_389),
.B(n_394),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_335),
.B(n_313),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_390),
.B(n_342),
.C(n_351),
.Y(n_429)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_308),
.Y(n_391)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_391),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_353),
.Y(n_392)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_392),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_341),
.Y(n_393)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_393),
.Y(n_436)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_347),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_355),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_395),
.B(n_397),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_351),
.B(n_220),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_315),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_346),
.A2(n_178),
.B1(n_146),
.B2(n_251),
.Y(n_398)
);

BUFx5_ASAP7_75t_L g399 ( 
.A(n_334),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_399),
.Y(n_412)
);

AO21x2_ASAP7_75t_SL g400 ( 
.A1(n_309),
.A2(n_343),
.B(n_350),
.Y(n_400)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_316),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_SL g439 ( 
.A1(n_402),
.A2(n_403),
.B1(n_242),
.B2(n_353),
.Y(n_439)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_316),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_384),
.B(n_313),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_404),
.B(n_429),
.C(n_432),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_405),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_358),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_406),
.B(n_407),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_356),
.Y(n_407)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_416),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_379),
.A2(n_313),
.B(n_342),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_417),
.A2(n_425),
.B(n_440),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_426),
.A2(n_438),
.B1(n_376),
.B2(n_360),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_375),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_427),
.B(n_367),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_390),
.B(n_328),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_380),
.B(n_304),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_435),
.B(n_442),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_400),
.A2(n_270),
.B1(n_296),
.B2(n_312),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_439),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_401),
.A2(n_333),
.B1(n_308),
.B2(n_338),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_382),
.B(n_369),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_382),
.B(n_299),
.C(n_339),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_443),
.B(n_376),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_437),
.A2(n_400),
.B1(n_401),
.B2(n_361),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_445),
.B(n_454),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_441),
.B(n_424),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_446),
.B(n_451),
.Y(n_502)
);

CKINVDCx14_ASAP7_75t_R g493 ( 
.A(n_447),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_448),
.A2(n_450),
.B1(n_467),
.B2(n_458),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_410),
.B(n_397),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_422),
.B(n_361),
.Y(n_452)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_452),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_422),
.B(n_366),
.Y(n_453)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_453),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_420),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_413),
.B(n_385),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_455),
.B(n_458),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_420),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_408),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_459),
.Y(n_499)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_408),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_460),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_437),
.A2(n_400),
.B1(n_373),
.B2(n_357),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_461),
.B(n_463),
.Y(n_506)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_430),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_462),
.Y(n_489)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_411),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_416),
.A2(n_396),
.B1(n_389),
.B2(n_365),
.Y(n_464)
);

A2O1A1Ixp33_ASAP7_75t_SL g508 ( 
.A1(n_464),
.A2(n_409),
.B(n_389),
.C(n_419),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_433),
.B(n_392),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_465),
.B(n_467),
.Y(n_500)
);

CKINVDCx10_ASAP7_75t_R g466 ( 
.A(n_412),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_466),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_420),
.Y(n_467)
);

INVx13_ASAP7_75t_L g469 ( 
.A(n_434),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_469),
.B(n_473),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_470),
.B(n_471),
.C(n_476),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_442),
.B(n_372),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_425),
.B(n_389),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_472),
.B(n_479),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_413),
.B(n_394),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_404),
.B(n_399),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_474),
.B(n_475),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_418),
.B(n_388),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_443),
.B(n_395),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_418),
.B(n_333),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_477),
.B(n_307),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_417),
.B(n_371),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_478),
.A2(n_428),
.B(n_409),
.Y(n_490)
);

INVx1_ASAP7_75t_SL g479 ( 
.A(n_435),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_468),
.B(n_432),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_482),
.B(n_484),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_468),
.B(n_429),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_457),
.B(n_405),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_485),
.B(n_486),
.C(n_487),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_457),
.B(n_426),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_471),
.B(n_476),
.Y(n_487)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_488),
.Y(n_526)
);

AOI21xp33_ASAP7_75t_L g524 ( 
.A1(n_490),
.A2(n_456),
.B(n_475),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_446),
.B(n_428),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_491),
.B(n_498),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_492),
.A2(n_509),
.B1(n_445),
.B2(n_460),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_444),
.B(n_434),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_470),
.B(n_438),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_504),
.B(n_515),
.C(n_494),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_452),
.B(n_359),
.Y(n_507)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_507),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_508),
.A2(n_450),
.B1(n_464),
.B2(n_456),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_448),
.A2(n_440),
.B1(n_409),
.B2(n_411),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_454),
.B(n_307),
.Y(n_510)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_510),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_472),
.B(n_449),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_512),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_449),
.A2(n_415),
.B(n_421),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_513),
.A2(n_514),
.B(n_414),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_472),
.A2(n_415),
.B(n_421),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_479),
.B(n_423),
.C(n_436),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_483),
.Y(n_516)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_516),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_499),
.B(n_455),
.Y(n_517)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_517),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_499),
.B(n_503),
.Y(n_518)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_518),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_SL g566 ( 
.A1(n_519),
.A2(n_508),
.B1(n_398),
.B2(n_383),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_503),
.B(n_473),
.Y(n_521)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_521),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_524),
.B(n_525),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_SL g525 ( 
.A(n_512),
.B(n_478),
.C(n_461),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_528),
.A2(n_531),
.B1(n_391),
.B2(n_469),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_485),
.B(n_453),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_529),
.B(n_539),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_495),
.A2(n_478),
.B1(n_480),
.B2(n_459),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_530),
.A2(n_490),
.B1(n_506),
.B2(n_495),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_509),
.A2(n_492),
.B1(n_512),
.B2(n_511),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_532),
.B(n_523),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_501),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_533),
.B(n_543),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_494),
.B(n_463),
.C(n_423),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_534),
.B(n_536),
.C(n_538),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_502),
.B(n_466),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g573 ( 
.A(n_535),
.B(n_306),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_484),
.B(n_436),
.C(n_403),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_486),
.B(n_402),
.C(n_370),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_487),
.B(n_430),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_482),
.B(n_431),
.C(n_414),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_540),
.B(n_547),
.C(n_513),
.Y(n_558)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_501),
.Y(n_541)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_541),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_L g564 ( 
.A1(n_542),
.A2(n_546),
.B(n_508),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_489),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_500),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_544),
.B(n_505),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_514),
.A2(n_462),
.B(n_431),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_515),
.B(n_338),
.C(n_339),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_529),
.B(n_493),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_SL g594 ( 
.A(n_549),
.B(n_552),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_516),
.B(n_481),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_517),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_553),
.B(n_559),
.Y(n_574)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_554),
.Y(n_581)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_556),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_558),
.B(n_566),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_534),
.B(n_504),
.C(n_511),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_530),
.A2(n_506),
.B1(n_497),
.B2(n_496),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_561),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_536),
.B(n_511),
.C(n_496),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_562),
.B(n_540),
.C(n_547),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_545),
.B(n_393),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_563),
.B(n_567),
.Y(n_595)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_564),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_532),
.B(n_508),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_569),
.B(n_523),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_570),
.A2(n_527),
.B1(n_537),
.B2(n_521),
.Y(n_577)
);

CKINVDCx16_ASAP7_75t_R g572 ( 
.A(n_518),
.Y(n_572)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_572),
.Y(n_586)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_573),
.Y(n_590)
);

AOI21xp33_ASAP7_75t_SL g575 ( 
.A1(n_560),
.A2(n_525),
.B(n_522),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_SL g602 ( 
.A1(n_575),
.A2(n_589),
.B(n_561),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_577),
.A2(n_587),
.B1(n_591),
.B2(n_564),
.Y(n_597)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_579),
.B(n_565),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_580),
.B(n_306),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g584 ( 
.A(n_571),
.B(n_526),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_584),
.A2(n_568),
.B(n_557),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_555),
.B(n_538),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_585),
.B(n_588),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_550),
.A2(n_528),
.B1(n_531),
.B2(n_546),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_555),
.B(n_520),
.C(n_539),
.Y(n_588)
);

NOR2xp67_ASAP7_75t_SL g589 ( 
.A(n_569),
.B(n_520),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_571),
.A2(n_542),
.B1(n_374),
.B2(n_312),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_551),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_592),
.B(n_593),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_558),
.B(n_325),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_SL g596 ( 
.A1(n_583),
.A2(n_570),
.B1(n_560),
.B2(n_548),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_596),
.B(n_598),
.Y(n_621)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_597),
.Y(n_620)
);

OAI21xp5_ASAP7_75t_L g598 ( 
.A1(n_582),
.A2(n_548),
.B(n_557),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_599),
.B(n_601),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_583),
.A2(n_562),
.B1(n_559),
.B2(n_556),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_600),
.A2(n_576),
.B1(n_578),
.B2(n_590),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_594),
.B(n_565),
.Y(n_601)
);

XOR2xp5_ASAP7_75t_L g629 ( 
.A(n_602),
.B(n_605),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_SL g603 ( 
.A(n_574),
.B(n_567),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_SL g624 ( 
.A(n_603),
.B(n_606),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_585),
.B(n_566),
.C(n_325),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_607),
.B(n_608),
.C(n_610),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_588),
.B(n_322),
.C(n_259),
.Y(n_608)
);

OAI21xp5_ASAP7_75t_SL g609 ( 
.A1(n_580),
.A2(n_354),
.B(n_225),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_609),
.B(n_613),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_593),
.B(n_242),
.C(n_296),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_595),
.B(n_298),
.C(n_257),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_611),
.B(n_614),
.C(n_225),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_581),
.B(n_354),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_579),
.B(n_298),
.C(n_257),
.Y(n_614)
);

OAI21xp5_ASAP7_75t_SL g615 ( 
.A1(n_596),
.A2(n_584),
.B(n_586),
.Y(n_615)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_615),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_617),
.B(n_618),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_SL g618 ( 
.A1(n_604),
.A2(n_578),
.B(n_576),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_612),
.B(n_252),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_619),
.B(n_623),
.Y(n_636)
);

NOR2xp67_ASAP7_75t_L g622 ( 
.A(n_600),
.B(n_354),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_622),
.B(n_611),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_608),
.B(n_252),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_627),
.B(n_628),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_605),
.B(n_277),
.C(n_290),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_620),
.B(n_625),
.C(n_629),
.Y(n_631)
);

XNOR2xp5_ASAP7_75t_L g641 ( 
.A(n_631),
.B(n_634),
.Y(n_641)
);

OA22x2_ASAP7_75t_L g632 ( 
.A1(n_621),
.A2(n_598),
.B1(n_599),
.B2(n_607),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_632),
.B(n_629),
.Y(n_644)
);

OAI21x1_ASAP7_75t_SL g643 ( 
.A1(n_633),
.A2(n_635),
.B(n_616),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_626),
.A2(n_614),
.B1(n_610),
.B2(n_292),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_624),
.A2(n_273),
.B1(n_248),
.B2(n_274),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g639 ( 
.A(n_625),
.B(n_225),
.C(n_274),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_639),
.B(n_628),
.C(n_627),
.Y(n_642)
);

OAI21xp5_ASAP7_75t_SL g640 ( 
.A1(n_615),
.A2(n_4),
.B(n_6),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_L g645 ( 
.A1(n_640),
.A2(n_4),
.B(n_6),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_642),
.B(n_647),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_SL g652 ( 
.A1(n_643),
.A2(n_644),
.B(n_646),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_645),
.B(n_648),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_L g646 ( 
.A1(n_637),
.A2(n_13),
.B(n_9),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_631),
.B(n_6),
.C(n_9),
.Y(n_647)
);

XOR2xp5_ASAP7_75t_L g648 ( 
.A(n_638),
.B(n_9),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g650 ( 
.A(n_641),
.B(n_630),
.C(n_632),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_650),
.B(n_653),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_L g653 ( 
.A1(n_642),
.A2(n_636),
.B(n_632),
.Y(n_653)
);

MAJx2_ASAP7_75t_L g654 ( 
.A(n_651),
.B(n_647),
.C(n_639),
.Y(n_654)
);

OAI21x1_ASAP7_75t_SL g657 ( 
.A1(n_654),
.A2(n_655),
.B(n_652),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_649),
.B(n_648),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_657),
.A2(n_656),
.B(n_640),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_658),
.B(n_635),
.C(n_12),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g660 ( 
.A(n_659),
.B(n_11),
.C(n_12),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_660),
.A2(n_13),
.B(n_358),
.Y(n_661)
);


endmodule