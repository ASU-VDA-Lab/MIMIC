module fake_jpeg_26366_n_414 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_414);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_414;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_9),
.B(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_44),
.B(n_60),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_25),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_46),
.B(n_47),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_31),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_25),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_50),
.B(n_53),
.Y(n_124)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_35),
.B(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_59),
.B(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_62),
.Y(n_123)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_15),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_33),
.B(n_14),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_74),
.B(n_77),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_33),
.B(n_13),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_21),
.B(n_11),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_37),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_23),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_79),
.B(n_82),
.Y(n_105)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_36),
.Y(n_92)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_26),
.B(n_11),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_92),
.B(n_97),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_43),
.B(n_23),
.C(n_16),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_44),
.B(n_36),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_99),
.B(n_114),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_27),
.B1(n_32),
.B2(n_37),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_100),
.A2(n_30),
.B1(n_18),
.B2(n_24),
.Y(n_130)
);

NAND2x1_ASAP7_75t_L g110 ( 
.A(n_55),
.B(n_37),
.Y(n_110)
);

OR2x2_ASAP7_75t_SL g133 ( 
.A(n_110),
.B(n_41),
.Y(n_133)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_62),
.A2(n_32),
.B1(n_27),
.B2(n_41),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_112),
.A2(n_76),
.B1(n_41),
.B2(n_24),
.Y(n_142)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_119),
.Y(n_128)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_127),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_78),
.B(n_18),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_125),
.B(n_96),
.Y(n_135)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_60),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_135),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_130),
.A2(n_142),
.B1(n_147),
.B2(n_150),
.Y(n_199)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_131),
.Y(n_184)
);

CKINVDCx12_ASAP7_75t_R g132 ( 
.A(n_110),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_132),
.Y(n_202)
);

OA21x2_ASAP7_75t_L g207 ( 
.A1(n_133),
.A2(n_166),
.B(n_113),
.Y(n_207)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_136),
.Y(n_175)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_137),
.B(n_158),
.Y(n_188)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_139),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_80),
.Y(n_140)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_140),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_90),
.B(n_91),
.Y(n_141)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_143),
.Y(n_182)
);

CKINVDCx12_ASAP7_75t_R g146 ( 
.A(n_94),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_98),
.A2(n_73),
.B1(n_48),
.B2(n_63),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_91),
.B(n_58),
.Y(n_148)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_101),
.Y(n_149)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_100),
.A2(n_68),
.B1(n_51),
.B2(n_56),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_23),
.Y(n_151)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_106),
.Y(n_153)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_153),
.Y(n_197)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_89),
.Y(n_154)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_154),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_20),
.B1(n_24),
.B2(n_17),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_155),
.A2(n_161),
.B1(n_115),
.B2(n_84),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_87),
.Y(n_156)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_156),
.Y(n_203)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_114),
.A2(n_30),
.B(n_20),
.C(n_17),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_116),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_104),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_163),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_112),
.A2(n_17),
.B1(n_20),
.B2(n_22),
.Y(n_161)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_93),
.Y(n_162)
);

INVx4_ASAP7_75t_SL g170 ( 
.A(n_162),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_10),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_86),
.B(n_10),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_165),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_100),
.B(n_16),
.Y(n_165)
);

O2A1O1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_85),
.A2(n_108),
.B(n_107),
.C(n_122),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_103),
.B(n_16),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_103),
.Y(n_186)
);

INVx11_ASAP7_75t_L g169 ( 
.A(n_93),
.Y(n_169)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_153),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_186),
.Y(n_208)
);

AOI32xp33_ASAP7_75t_L g174 ( 
.A1(n_132),
.A2(n_55),
.A3(n_57),
.B1(n_52),
.B2(n_45),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_SL g241 ( 
.A(n_174),
.B(n_113),
.C(n_57),
.Y(n_241)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_185),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_146),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_194),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_190),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_134),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_128),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_196),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_144),
.B(n_123),
.Y(n_196)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_169),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_205),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_147),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_206),
.A2(n_166),
.B1(n_159),
.B2(n_83),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_207),
.A2(n_28),
.B(n_155),
.Y(n_239)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_170),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_209),
.A2(n_221),
.B1(n_181),
.B2(n_104),
.Y(n_268)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_173),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_210),
.B(n_212),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_175),
.Y(n_211)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_211),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_201),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_179),
.B(n_165),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_28),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_199),
.A2(n_145),
.B1(n_157),
.B2(n_139),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_215),
.A2(n_232),
.B1(n_238),
.B2(n_197),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_144),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_216),
.B(n_217),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_207),
.Y(n_217)
);

NOR2x1_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_130),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_218),
.B(n_229),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_192),
.A2(n_168),
.B1(n_161),
.B2(n_129),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_220),
.A2(n_225),
.B1(n_230),
.B2(n_156),
.Y(n_262)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_167),
.C(n_137),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_228),
.C(n_172),
.Y(n_249)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_223),
.B(n_231),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_178),
.A2(n_145),
.B1(n_115),
.B2(n_136),
.Y(n_225)
);

INVx13_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_226),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_177),
.B(n_167),
.C(n_131),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_176),
.B(n_133),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_203),
.A2(n_138),
.B1(n_84),
.B2(n_83),
.Y(n_230)
);

NAND3xp33_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_135),
.C(n_158),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_170),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

CKINVDCx11_ASAP7_75t_R g235 ( 
.A(n_180),
.Y(n_235)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_191),
.Y(n_236)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_236),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_187),
.B(n_160),
.Y(n_237)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_185),
.A2(n_152),
.B1(n_143),
.B2(n_123),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_171),
.B1(n_197),
.B2(n_200),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_162),
.Y(n_240)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_240),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_241),
.A2(n_242),
.B(n_113),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_172),
.B(n_49),
.Y(n_242)
);

AOI32xp33_ASAP7_75t_L g243 ( 
.A1(n_229),
.A2(n_191),
.A3(n_204),
.B1(n_180),
.B2(n_61),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_243),
.B(n_273),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_228),
.B(n_184),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_244),
.B(n_253),
.Y(n_281)
);

MAJx2_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_61),
.C(n_28),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_245),
.B(n_246),
.Y(n_279)
);

NOR2xp67_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_22),
.Y(n_248)
);

NOR2xp67_ASAP7_75t_L g295 ( 
.A(n_248),
.B(n_225),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_249),
.B(n_261),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_250),
.A2(n_252),
.B1(n_262),
.B2(n_270),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_217),
.A2(n_182),
.B1(n_183),
.B2(n_200),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_183),
.Y(n_254)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_254),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_214),
.B(n_182),
.C(n_193),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_255),
.B(n_259),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_258),
.A2(n_239),
.B1(n_211),
.B2(n_208),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_210),
.B(n_224),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_218),
.A2(n_156),
.B1(n_181),
.B2(n_175),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_263),
.A2(n_269),
.B1(n_232),
.B2(n_211),
.Y(n_284)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_240),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_272),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_268),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_218),
.A2(n_22),
.B1(n_72),
.B2(n_71),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_209),
.A2(n_93),
.B1(n_1),
.B2(n_2),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_227),
.A2(n_22),
.B(n_1),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_237),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_251),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_276),
.B(n_281),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_277),
.A2(n_271),
.B1(n_267),
.B2(n_255),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_224),
.Y(n_282)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_282),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_260),
.B(n_259),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_283),
.B(n_219),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_284),
.A2(n_257),
.B1(n_230),
.B2(n_213),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_220),
.Y(n_285)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_285),
.Y(n_310)
);

OA22x2_ASAP7_75t_L g287 ( 
.A1(n_269),
.A2(n_235),
.B1(n_221),
.B2(n_241),
.Y(n_287)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_287),
.Y(n_318)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_265),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_288),
.B(n_296),
.Y(n_323)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_251),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_289),
.B(n_297),
.Y(n_320)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_252),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_292),
.Y(n_304)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_254),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_254),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_294),
.Y(n_307)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_262),
.Y(n_294)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_295),
.Y(n_317)
);

AND2x6_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_242),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_274),
.Y(n_297)
);

AND2x6_ASAP7_75t_L g298 ( 
.A(n_264),
.B(n_242),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_256),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_256),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_303),
.A2(n_306),
.B1(n_324),
.B2(n_285),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_301),
.B(n_246),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_305),
.B(n_315),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_294),
.A2(n_266),
.B1(n_208),
.B2(n_249),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_279),
.B(n_245),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_309),
.B(n_314),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_311),
.B(n_234),
.Y(n_342)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_312),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_279),
.B(n_261),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_272),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_316),
.A2(n_291),
.B1(n_293),
.B2(n_287),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_282),
.B(n_257),
.Y(n_319)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_319),
.Y(n_340)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_275),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_325),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_275),
.Y(n_322)
);

INVxp33_ASAP7_75t_L g329 ( 
.A(n_322),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_286),
.A2(n_219),
.B1(n_247),
.B2(n_265),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_278),
.B(n_234),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_323),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_327),
.B(n_0),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_280),
.C(n_290),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_328),
.B(n_330),
.C(n_341),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_290),
.C(n_292),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_331),
.A2(n_332),
.B1(n_334),
.B2(n_304),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_308),
.A2(n_299),
.B1(n_284),
.B2(n_285),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_333),
.A2(n_310),
.B1(n_302),
.B2(n_316),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_308),
.A2(n_321),
.B1(n_318),
.B2(n_317),
.Y(n_334)
);

OA21x2_ASAP7_75t_L g336 ( 
.A1(n_318),
.A2(n_296),
.B(n_298),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_336),
.A2(n_213),
.B(n_11),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_314),
.B(n_300),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_337),
.B(n_338),
.Y(n_348)
);

XNOR2x1_ASAP7_75t_L g338 ( 
.A(n_309),
.B(n_287),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_312),
.B(n_223),
.C(n_287),
.Y(n_341)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_342),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_313),
.B(n_320),
.Y(n_343)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_343),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_319),
.B(n_288),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_345),
.B(n_226),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_327),
.B(n_302),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g366 ( 
.A(n_346),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_347),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_338),
.A2(n_310),
.B1(n_307),
.B2(n_304),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_349),
.A2(n_357),
.B1(n_360),
.B2(n_335),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_326),
.B(n_307),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_350),
.B(n_359),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_353),
.B(n_362),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_354),
.A2(n_361),
.B(n_340),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_345),
.B(n_226),
.C(n_10),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_355),
.B(n_330),
.C(n_328),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_356),
.B(n_339),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_341),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_357)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_336),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_336),
.A2(n_2),
.B(n_4),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_337),
.B(n_4),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_355),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_363),
.B(n_365),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_367),
.B(n_369),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_368),
.B(n_348),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_351),
.B(n_344),
.C(n_339),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_371),
.B(n_372),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_351),
.B(n_344),
.C(n_329),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_352),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_374),
.B(n_375),
.Y(n_380)
);

NOR3xp33_ASAP7_75t_SL g375 ( 
.A(n_361),
.B(n_329),
.C(n_6),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_372),
.A2(n_354),
.B(n_358),
.Y(n_377)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_377),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_366),
.A2(n_349),
.B(n_356),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_379),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_367),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_381),
.B(n_387),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_382),
.B(n_384),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_365),
.B(n_348),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_383),
.B(n_386),
.Y(n_391)
);

INVxp33_ASAP7_75t_SL g384 ( 
.A(n_375),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_370),
.B(n_362),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_370),
.B(n_347),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_385),
.B(n_371),
.C(n_374),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_388),
.B(n_395),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_382),
.B(n_368),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_393),
.B(n_396),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_376),
.B(n_364),
.C(n_373),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_381),
.B(n_5),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_391),
.B(n_378),
.C(n_380),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_398),
.B(n_400),
.C(n_402),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_396),
.B(n_384),
.Y(n_399)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_399),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_389),
.A2(n_392),
.B(n_394),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_390),
.B(n_5),
.Y(n_402)
);

NOR3xp33_ASAP7_75t_SL g403 ( 
.A(n_401),
.B(n_390),
.C(n_393),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_403),
.B(n_405),
.Y(n_407)
);

AOI32xp33_ASAP7_75t_L g405 ( 
.A1(n_397),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_399),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_406),
.B(n_7),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_408),
.B(n_7),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_409),
.B(n_407),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_410),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_411),
.B(n_404),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_412),
.B(n_8),
.Y(n_413)
);

BUFx24_ASAP7_75t_SL g414 ( 
.A(n_413),
.Y(n_414)
);


endmodule