module fake_jpeg_8636_n_207 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_207);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_207;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_38),
.Y(n_49)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_0),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_L g64 ( 
.A1(n_36),
.A2(n_37),
.B(n_41),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_16),
.B(n_2),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_39),
.Y(n_65)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_43),
.Y(n_52)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_37),
.B(n_20),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_45),
.B(n_58),
.Y(n_72)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_24),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_51),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_24),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_21),
.B(n_27),
.C(n_16),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_21),
.B(n_32),
.C(n_27),
.Y(n_68)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_61),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_32),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_24),
.B1(n_18),
.B2(n_28),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_25),
.B1(n_28),
.B2(n_19),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_31),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_62),
.Y(n_71)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_67),
.A2(n_30),
.B1(n_31),
.B2(n_22),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_83),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_65),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_73),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_17),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_76),
.Y(n_102)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_28),
.B1(n_25),
.B2(n_17),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_74),
.A2(n_30),
.B1(n_63),
.B2(n_47),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_31),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_56),
.A2(n_50),
.B1(n_60),
.B2(n_62),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_60),
.B1(n_47),
.B2(n_57),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_54),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_82),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_44),
.C(n_38),
.Y(n_83)
);

NAND2xp33_ASAP7_75t_SL g85 ( 
.A(n_65),
.B(n_26),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_85),
.A2(n_26),
.B(n_54),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_89),
.B(n_105),
.Y(n_109)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_92),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_96),
.Y(n_110)
);

OAI22x1_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_65),
.B1(n_31),
.B2(n_29),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_95),
.A2(n_106),
.B(n_85),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_100),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_73),
.A2(n_44),
.B1(n_58),
.B2(n_26),
.Y(n_98)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_68),
.A2(n_26),
.B1(n_29),
.B2(n_38),
.Y(n_99)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_26),
.B1(n_22),
.B2(n_29),
.Y(n_101)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_53),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_104),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g104 ( 
.A(n_80),
.B(n_54),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_71),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_103),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_118),
.C(n_120),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_104),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_114),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_81),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_77),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_81),
.Y(n_120)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_76),
.Y(n_121)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

NOR2xp67_ASAP7_75t_R g132 ( 
.A(n_122),
.B(n_95),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_87),
.B(n_72),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_66),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_70),
.Y(n_126)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_66),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_127),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_123),
.A2(n_96),
.B1(n_101),
.B2(n_106),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_129),
.A2(n_131),
.B1(n_134),
.B2(n_124),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_116),
.A2(n_99),
.B1(n_89),
.B2(n_98),
.Y(n_131)
);

AOI321xp33_ASAP7_75t_L g151 ( 
.A1(n_132),
.A2(n_122),
.A3(n_121),
.B1(n_115),
.B2(n_26),
.C(n_23),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_123),
.A2(n_116),
.B1(n_124),
.B2(n_109),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_141),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_86),
.Y(n_136)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_144),
.C(n_82),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_110),
.Y(n_141)
);

A2O1A1O1Ixp25_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_102),
.B(n_70),
.C(n_97),
.D(n_69),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_126),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_78),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_143),
.B(n_119),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_102),
.C(n_71),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_128),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_147),
.Y(n_166)
);

AOI221xp5_ASAP7_75t_L g161 ( 
.A1(n_148),
.A2(n_160),
.B1(n_139),
.B2(n_142),
.C(n_141),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_149),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_112),
.Y(n_150)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_158),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_115),
.B1(n_91),
.B2(n_107),
.Y(n_152)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_156),
.C(n_159),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_144),
.C(n_140),
.Y(n_156)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_157),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_23),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_38),
.Y(n_159)
);

OAI321xp33_ASAP7_75t_L g160 ( 
.A1(n_133),
.A2(n_23),
.A3(n_15),
.B1(n_13),
.B2(n_12),
.C(n_11),
.Y(n_160)
);

AOI321xp33_ASAP7_75t_L g176 ( 
.A1(n_161),
.A2(n_157),
.A3(n_23),
.B1(n_53),
.B2(n_6),
.C(n_7),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_140),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_173),
.C(n_159),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_130),
.B(n_138),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_171),
.B1(n_149),
.B2(n_158),
.Y(n_174)
);

AOI321xp33_ASAP7_75t_L g170 ( 
.A1(n_151),
.A2(n_145),
.A3(n_138),
.B1(n_131),
.B2(n_23),
.C(n_12),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_53),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_154),
.A2(n_145),
.B(n_155),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_53),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_176),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_178),
.C(n_180),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_3),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_177),
.A2(n_4),
.B(n_5),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_173),
.C(n_165),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_183),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_3),
.Y(n_180)
);

INVxp33_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_169),
.Y(n_184)
);

MAJx2_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_170),
.C(n_167),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_182),
.A2(n_168),
.B1(n_162),
.B2(n_172),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_10),
.C(n_5),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_188),
.Y(n_193)
);

FAx1_ASAP7_75t_SL g196 ( 
.A(n_186),
.B(n_10),
.CI(n_8),
.CON(n_196),
.SN(n_196)
);

INVx11_ASAP7_75t_L g188 ( 
.A(n_181),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_189),
.A2(n_4),
.B(n_6),
.Y(n_192)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_190),
.A2(n_182),
.B1(n_6),
.B2(n_7),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_192),
.A2(n_197),
.B(n_189),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_185),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_4),
.C(n_7),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_191),
.C(n_186),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_196),
.A2(n_187),
.B(n_9),
.Y(n_200)
);

OAI21x1_ASAP7_75t_L g197 ( 
.A1(n_190),
.A2(n_185),
.B(n_184),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_199),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_200),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_201),
.B(n_193),
.C(n_196),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_204),
.B(n_202),
.C(n_8),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_203),
.A2(n_193),
.B(n_188),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_205),
.B(n_206),
.Y(n_207)
);


endmodule