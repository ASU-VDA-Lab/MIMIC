module real_jpeg_18876_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_0),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_0),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_0),
.A2(n_101),
.B1(n_267),
.B2(n_269),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_0),
.A2(n_101),
.B1(n_327),
.B2(n_329),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_1),
.A2(n_66),
.B1(n_70),
.B2(n_71),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_1),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_1),
.A2(n_31),
.B1(n_70),
.B2(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_1),
.A2(n_70),
.B1(n_341),
.B2(n_344),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_1),
.A2(n_70),
.B1(n_352),
.B2(n_354),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_2),
.A2(n_217),
.B1(n_220),
.B2(n_221),
.Y(n_216)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_2),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_3),
.Y(n_88)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_4),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_4),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_4),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_4),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_5),
.A2(n_171),
.B1(n_175),
.B2(n_177),
.Y(n_170)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_5),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_6),
.A2(n_110),
.B1(n_111),
.B2(n_114),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_6),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_6),
.A2(n_110),
.B1(n_248),
.B2(n_250),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_6),
.A2(n_110),
.B1(n_285),
.B2(n_290),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_7),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_7),
.Y(n_146)
);

OAI22x1_ASAP7_75t_SL g200 ( 
.A1(n_7),
.A2(n_146),
.B1(n_201),
.B2(n_203),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_8),
.A2(n_26),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_8),
.A2(n_58),
.B1(n_193),
.B2(n_197),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_8),
.A2(n_58),
.B1(n_317),
.B2(n_322),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_8),
.A2(n_58),
.B1(n_176),
.B2(n_374),
.Y(n_373)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_9),
.Y(n_157)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_9),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g379 ( 
.A(n_9),
.Y(n_379)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_10),
.B(n_62),
.Y(n_210)
);

OAI32xp33_ASAP7_75t_L g276 ( 
.A1(n_10),
.A2(n_75),
.A3(n_111),
.B1(n_277),
.B2(n_280),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_10),
.B(n_107),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_10),
.A2(n_154),
.B1(n_225),
.B2(n_373),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_10),
.A2(n_28),
.B1(n_393),
.B2(n_395),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_11),
.Y(n_93)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_11),
.Y(n_98)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_11),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_11),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_11),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_11),
.Y(n_235)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_11),
.Y(n_321)
);

OAI22xp33_ASAP7_75t_L g160 ( 
.A1(n_12),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_12),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_12),
.A2(n_162),
.B1(n_230),
.B2(n_232),
.Y(n_229)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_14),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_15),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_15),
.Y(n_128)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_15),
.Y(n_167)
);

BUFx4f_ASAP7_75t_L g174 ( 
.A(n_15),
.Y(n_174)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_255),
.B1(n_256),
.B2(n_411),
.Y(n_18)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_19),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_254),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_211),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_22),
.B(n_211),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_152),
.C(n_189),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_23),
.B(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_63),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_24),
.B(n_64),
.C(n_108),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_34),
.B1(n_57),
.B2(n_62),
.Y(n_24)
);

OAI21xp33_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_28),
.B(n_29),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_28),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_28),
.B(n_302),
.Y(n_301)
);

OAI21xp33_ASAP7_75t_SL g312 ( 
.A1(n_28),
.A2(n_301),
.B(n_313),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_28),
.B(n_207),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_28),
.B(n_151),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_29),
.A2(n_179),
.B1(n_186),
.B2(n_188),
.Y(n_178)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_34),
.A2(n_57),
.B1(n_62),
.B2(n_241),
.Y(n_240)
);

OA21x2_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_42),
.B(n_45),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_39),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_42),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_43),
.Y(n_180)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

AOI22x1_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_49),
.B1(n_52),
.B2(n_55),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_51),
.Y(n_196)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_61),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_108),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_73),
.B1(n_99),
.B2(n_107),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_65),
.A2(n_73),
.B1(n_107),
.B2(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_69),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_74),
.A2(n_246),
.B1(n_247),
.B2(n_252),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_74),
.A2(n_192),
.B1(n_252),
.B2(n_392),
.Y(n_391)
);

AO21x2_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_84),
.B(n_92),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_83),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_89),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g231 ( 
.A(n_93),
.Y(n_231)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_93),
.Y(n_268)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx6_ASAP7_75t_L g298 ( 
.A(n_97),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVxp67_ASAP7_75t_SL g113 ( 
.A(n_98),
.Y(n_113)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_99),
.Y(n_246)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_105),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_106),
.Y(n_185)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_107),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_119),
.B1(n_142),
.B2(n_150),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_109),
.Y(n_273)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_116),
.Y(n_281)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_119),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_119),
.A2(n_150),
.B1(n_312),
.B2(n_316),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_119),
.A2(n_150),
.B1(n_316),
.B2(n_340),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_119),
.A2(n_150),
.B1(n_266),
.B2(n_340),
.Y(n_401)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_131),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_124),
.B1(n_126),
.B2(n_129),
.Y(n_120)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_125),
.Y(n_202)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_125),
.Y(n_219)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_125),
.Y(n_289)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_128),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_128),
.Y(n_353)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_128),
.Y(n_370)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_130),
.Y(n_306)
);

OAI22xp33_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_136),
.B1(n_139),
.B2(n_141),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_135),
.Y(n_272)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_139),
.Y(n_300)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_143),
.A2(n_151),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_148),
.Y(n_345)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_151),
.A2(n_228),
.B1(n_265),
.B2(n_273),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_152),
.B(n_189),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_178),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_153),
.B(n_178),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_159),
.B1(n_168),
.B2(n_170),
.Y(n_153)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_154),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_154),
.A2(n_170),
.B1(n_216),
.B2(n_225),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_154),
.A2(n_326),
.B1(n_334),
.B2(n_335),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_154),
.A2(n_351),
.B1(n_373),
.B2(n_377),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_157),
.Y(n_334)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_158),
.Y(n_161)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_158),
.Y(n_299)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI22x1_ASAP7_75t_SL g198 ( 
.A1(n_160),
.A2(n_199),
.B1(n_200),
.B2(n_206),
.Y(n_198)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_166),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_167),
.Y(n_224)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_173),
.Y(n_290)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_174),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_174),
.Y(n_328)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_185),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_187),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_198),
.C(n_210),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_190),
.B(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx2_ASAP7_75t_SL g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_196),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_198),
.B(n_210),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_199),
.A2(n_200),
.B1(n_226),
.B2(n_284),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_199),
.A2(n_350),
.B1(n_357),
.B2(n_358),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_201),
.Y(n_374)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_208),
.Y(n_226)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_236),
.B1(n_237),
.B2(n_253),
.Y(n_211)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_212),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

XOR2x2_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_227),
.Y(n_214)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_225),
.Y(n_357)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_245),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

AOI21x1_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_291),
.B(n_410),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_258),
.B(n_260),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_264),
.C(n_274),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_261),
.A2(n_262),
.B1(n_405),
.B2(n_406),
.Y(n_404)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_264),
.A2(n_274),
.B1(n_275),
.B2(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_264),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_268),
.Y(n_315)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_282),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_276),
.A2(n_282),
.B1(n_283),
.B2(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_276),
.Y(n_388)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_281),
.Y(n_302)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_284),
.Y(n_335)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI21x1_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_403),
.B(n_409),
.Y(n_291)
);

AOI21x1_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_384),
.B(n_402),
.Y(n_292)
);

OAI21x1_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_347),
.B(n_383),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_324),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_295),
.B(n_324),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_310),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_296),
.A2(n_310),
.B1(n_311),
.B2(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_296),
.Y(n_360)
);

OAI32xp33_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_299),
.A3(n_300),
.B1(n_301),
.B2(n_303),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_307),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_321),
.Y(n_323)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_321),
.Y(n_343)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_336),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_325),
.B(n_338),
.C(n_346),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_326),
.Y(n_358)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_338),
.B1(n_339),
.B2(n_346),
.Y(n_336)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_337),
.Y(n_346)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_361),
.B(n_382),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_359),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_349),
.B(n_359),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_SL g355 ( 
.A(n_356),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_375),
.B(n_381),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_372),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_371),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_380),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_376),
.B(n_380),
.Y(n_381)
);

INVx6_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

BUFx12f_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_386),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_385),
.B(n_386),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_389),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_387),
.B(n_390),
.C(n_401),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_390),
.A2(n_391),
.B1(n_400),
.B2(n_401),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

NOR2xp67_ASAP7_75t_SL g403 ( 
.A(n_404),
.B(n_408),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_404),
.B(n_408),
.Y(n_409)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);


endmodule