module fake_jpeg_184_n_130 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_130);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx6_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_33),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_50),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_0),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_51),
.B(n_52),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_1),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_54),
.B(n_47),
.Y(n_61)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_48),
.B(n_40),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_58),
.B(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_66),
.B(n_70),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_2),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_59),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_40),
.C(n_46),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_36),
.C(n_12),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_76),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_34),
.B1(n_37),
.B2(n_35),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_59),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_46),
.B1(n_37),
.B2(n_34),
.Y(n_76)
);

INVxp33_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_77),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_55),
.B(n_57),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_78),
.A2(n_85),
.B(n_8),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_81),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_1),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_2),
.Y(n_83)
);

NOR3xp33_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_36),
.C(n_4),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_90),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_3),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_89),
.B(n_8),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_4),
.Y(n_90)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_77),
.B1(n_71),
.B2(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_93),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_84),
.A2(n_71),
.B1(n_6),
.B2(n_7),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_92),
.A2(n_94),
.B1(n_103),
.B2(n_101),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_88),
.B(n_14),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_80),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_97),
.B(n_100),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_16),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_15),
.Y(n_115)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_85),
.B(n_17),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_103),
.B(n_9),
.Y(n_111)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_29),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_110),
.C(n_115),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_93),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_113),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_96),
.C(n_19),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_SL g121 ( 
.A1(n_118),
.A2(n_119),
.B(n_24),
.C(n_25),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_96),
.C(n_21),
.Y(n_119)
);

AOI21x1_ASAP7_75t_L g124 ( 
.A1(n_121),
.A2(n_122),
.B(n_123),
.Y(n_124)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_123),
.B(n_107),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_117),
.B1(n_105),
.B2(n_114),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_124),
.B1(n_106),
.B2(n_112),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_111),
.B(n_11),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_10),
.B(n_11),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_10),
.Y(n_130)
);


endmodule