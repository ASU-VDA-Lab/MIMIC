module fake_aes_8690_n_14 (n_1, n_2, n_0, n_14);
input n_1;
input n_2;
input n_0;
output n_14;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
NOR2xp33_ASAP7_75t_L g3 ( .A(n_0), .B(n_2), .Y(n_3) );
INVx5_ASAP7_75t_L g4 ( .A(n_1), .Y(n_4) );
HB1xp67_ASAP7_75t_L g5 ( .A(n_2), .Y(n_5) );
OAI22xp5_ASAP7_75t_L g6 ( .A1(n_5), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_6) );
BUFx3_ASAP7_75t_L g7 ( .A(n_4), .Y(n_7) );
AOI211xp5_ASAP7_75t_L g8 ( .A1(n_6), .A2(n_3), .B(n_1), .C(n_2), .Y(n_8) );
AOI33xp33_ASAP7_75t_L g9 ( .A1(n_7), .A2(n_0), .A3(n_1), .B1(n_2), .B2(n_4), .B3(n_6), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
NAND2xp5_ASAP7_75t_L g11 ( .A(n_8), .B(n_4), .Y(n_11) );
NAND3xp33_ASAP7_75t_L g12 ( .A(n_10), .B(n_8), .C(n_4), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
OR2x6_ASAP7_75t_L g14 ( .A(n_13), .B(n_11), .Y(n_14) );
endmodule