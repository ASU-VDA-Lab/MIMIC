module fake_netlist_1_702_n_657 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_657);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_657;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx2_ASAP7_75t_L g75 ( .A(n_30), .Y(n_75) );
INVxp67_ASAP7_75t_L g76 ( .A(n_66), .Y(n_76) );
CKINVDCx20_ASAP7_75t_R g77 ( .A(n_2), .Y(n_77) );
HB1xp67_ASAP7_75t_L g78 ( .A(n_41), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_15), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_38), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_10), .Y(n_81) );
INVxp33_ASAP7_75t_SL g82 ( .A(n_11), .Y(n_82) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_61), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_34), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_59), .Y(n_85) );
CKINVDCx16_ASAP7_75t_R g86 ( .A(n_40), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_14), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_71), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_50), .Y(n_89) );
OR2x2_ASAP7_75t_L g90 ( .A(n_46), .B(n_2), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_4), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_55), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_20), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_6), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_24), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_58), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_9), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_60), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_16), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_63), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_69), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_29), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_25), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_5), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_23), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_37), .Y(n_106) );
INVxp33_ASAP7_75t_L g107 ( .A(n_5), .Y(n_107) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_1), .Y(n_108) );
INVx1_ASAP7_75t_SL g109 ( .A(n_13), .Y(n_109) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_68), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_65), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_62), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_36), .B(n_33), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_44), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_0), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_49), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_8), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_18), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_57), .Y(n_119) );
INVxp67_ASAP7_75t_L g120 ( .A(n_28), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_84), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_85), .Y(n_122) );
AND2x4_ASAP7_75t_L g123 ( .A(n_75), .B(n_0), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_85), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_108), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_93), .Y(n_126) );
BUFx2_ASAP7_75t_L g127 ( .A(n_75), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_93), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_96), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_84), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_89), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_89), .Y(n_132) );
INVxp67_ASAP7_75t_L g133 ( .A(n_94), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_78), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_110), .B(n_1), .Y(n_135) );
OAI22xp5_ASAP7_75t_L g136 ( .A1(n_107), .A2(n_3), .B1(n_4), .B2(n_6), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_96), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_79), .B(n_3), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_103), .Y(n_139) );
AND2x6_ASAP7_75t_L g140 ( .A(n_103), .B(n_35), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_100), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_79), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_81), .B(n_7), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_114), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_100), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_81), .B(n_7), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_87), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_114), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_116), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_116), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_118), .B(n_8), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_97), .B(n_9), .Y(n_152) );
AND2x6_ASAP7_75t_L g153 ( .A(n_118), .B(n_42), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_119), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_119), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_80), .Y(n_156) );
OAI21x1_ASAP7_75t_L g157 ( .A1(n_95), .A2(n_43), .B(n_73), .Y(n_157) );
NAND2xp33_ASAP7_75t_SL g158 ( .A(n_90), .B(n_10), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_99), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_87), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_82), .B(n_11), .Y(n_161) );
INVxp67_ASAP7_75t_L g162 ( .A(n_91), .Y(n_162) );
BUFx4f_ASAP7_75t_L g163 ( .A(n_140), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_141), .Y(n_164) );
AND2x6_ASAP7_75t_L g165 ( .A(n_123), .B(n_102), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_134), .B(n_120), .Y(n_166) );
OR2x2_ASAP7_75t_L g167 ( .A(n_127), .B(n_125), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_127), .B(n_86), .Y(n_168) );
INVx1_ASAP7_75t_SL g169 ( .A(n_143), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_123), .B(n_117), .Y(n_170) );
INVx4_ASAP7_75t_L g171 ( .A(n_140), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_162), .B(n_117), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_133), .B(n_115), .Y(n_173) );
NOR2xp33_ASAP7_75t_SL g174 ( .A(n_140), .B(n_106), .Y(n_174) );
INVx1_ASAP7_75t_SL g175 ( .A(n_146), .Y(n_175) );
OAI22xp5_ASAP7_75t_SL g176 ( .A1(n_136), .A2(n_77), .B1(n_83), .B2(n_105), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_121), .B(n_92), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_123), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_138), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_141), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_147), .B(n_76), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_138), .Y(n_182) );
NOR3xp33_ASAP7_75t_SL g183 ( .A(n_158), .B(n_112), .C(n_92), .Y(n_183) );
OAI21xp33_ASAP7_75t_L g184 ( .A1(n_121), .A2(n_115), .B(n_91), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_141), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_160), .B(n_142), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_130), .B(n_101), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_138), .Y(n_188) );
OAI22xp5_ASAP7_75t_L g189 ( .A1(n_130), .A2(n_104), .B1(n_90), .B2(n_109), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_141), .Y(n_190) );
AND2x2_ASAP7_75t_SL g191 ( .A(n_135), .B(n_104), .Y(n_191) );
BUFx3_ASAP7_75t_L g192 ( .A(n_140), .Y(n_192) );
INVx3_ASAP7_75t_L g193 ( .A(n_142), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_141), .Y(n_194) );
NAND2x1p5_ASAP7_75t_L g195 ( .A(n_151), .B(n_113), .Y(n_195) );
AO22x2_ASAP7_75t_L g196 ( .A1(n_131), .A2(n_111), .B1(n_88), .B2(n_14), .Y(n_196) );
AND2x4_ASAP7_75t_L g197 ( .A(n_142), .B(n_112), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_158), .Y(n_198) );
AO21x2_ASAP7_75t_L g199 ( .A1(n_157), .A2(n_98), .B(n_47), .Y(n_199) );
AND2x4_ASAP7_75t_SL g200 ( .A(n_161), .B(n_98), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_131), .B(n_12), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_148), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_132), .B(n_12), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_132), .B(n_13), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_150), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_139), .B(n_15), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_148), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_139), .B(n_17), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_157), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_152), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_148), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_148), .Y(n_212) );
BUFx3_ASAP7_75t_L g213 ( .A(n_140), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_148), .Y(n_214) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_140), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_153), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_144), .B(n_19), .Y(n_217) );
BUFx4f_ASAP7_75t_L g218 ( .A(n_165), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_193), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_193), .Y(n_220) );
AND2x2_ASAP7_75t_SL g221 ( .A(n_174), .B(n_155), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_193), .Y(n_222) );
INVx3_ASAP7_75t_L g223 ( .A(n_204), .Y(n_223) );
AND2x6_ASAP7_75t_SL g224 ( .A(n_168), .B(n_155), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_204), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_186), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_202), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_210), .Y(n_228) );
BUFx3_ASAP7_75t_L g229 ( .A(n_192), .Y(n_229) );
BUFx3_ASAP7_75t_L g230 ( .A(n_192), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_167), .B(n_144), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_186), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_204), .Y(n_233) );
AOI22x1_ASAP7_75t_L g234 ( .A1(n_209), .A2(n_159), .B1(n_156), .B2(n_150), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_177), .B(n_154), .Y(n_235) );
INVx4_ASAP7_75t_L g236 ( .A(n_165), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_206), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_206), .Y(n_238) );
AND2x4_ASAP7_75t_L g239 ( .A(n_170), .B(n_159), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_206), .Y(n_240) );
AOI22xp5_ASAP7_75t_L g241 ( .A1(n_178), .A2(n_175), .B1(n_169), .B2(n_191), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_205), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_215), .Y(n_243) );
BUFx8_ASAP7_75t_L g244 ( .A(n_167), .Y(n_244) );
INVx3_ASAP7_75t_L g245 ( .A(n_165), .Y(n_245) );
AOI22xp5_ASAP7_75t_L g246 ( .A1(n_178), .A2(n_154), .B1(n_149), .B2(n_153), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_171), .B(n_149), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g248 ( .A1(n_191), .A2(n_153), .B1(n_156), .B2(n_145), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_179), .Y(n_249) );
BUFx8_ASAP7_75t_L g250 ( .A(n_165), .Y(n_250) );
INVx4_ASAP7_75t_L g251 ( .A(n_165), .Y(n_251) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_215), .Y(n_252) );
BUFx4f_ASAP7_75t_SL g253 ( .A(n_165), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_171), .B(n_128), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_182), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_172), .B(n_128), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_202), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_188), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_198), .A2(n_153), .B1(n_145), .B2(n_137), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g260 ( .A1(n_198), .A2(n_153), .B1(n_137), .B2(n_129), .Y(n_260) );
INVx5_ASAP7_75t_L g261 ( .A(n_185), .Y(n_261) );
AND2x4_ASAP7_75t_L g262 ( .A(n_170), .B(n_153), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_197), .B(n_129), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_197), .Y(n_264) );
BUFx4f_ASAP7_75t_L g265 ( .A(n_197), .Y(n_265) );
INVx1_ASAP7_75t_SL g266 ( .A(n_210), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_183), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_207), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_172), .B(n_126), .Y(n_269) );
NAND3xp33_ASAP7_75t_L g270 ( .A(n_166), .B(n_126), .C(n_124), .Y(n_270) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_173), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_170), .B(n_124), .Y(n_272) );
INVx1_ASAP7_75t_SL g273 ( .A(n_173), .Y(n_273) );
INVx3_ASAP7_75t_L g274 ( .A(n_171), .Y(n_274) );
INVx3_ASAP7_75t_L g275 ( .A(n_215), .Y(n_275) );
INVxp67_ASAP7_75t_SL g276 ( .A(n_215), .Y(n_276) );
INVx3_ASAP7_75t_L g277 ( .A(n_216), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_219), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_219), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_243), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_222), .Y(n_281) );
BUFx2_ASAP7_75t_L g282 ( .A(n_250), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_222), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_243), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_236), .B(n_213), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_244), .Y(n_286) );
INVx2_ASAP7_75t_SL g287 ( .A(n_265), .Y(n_287) );
AOI221xp5_ASAP7_75t_SL g288 ( .A1(n_264), .A2(n_189), .B1(n_184), .B2(n_181), .C(n_187), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_223), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_243), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_244), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_231), .B(n_196), .Y(n_292) );
BUFx12f_ASAP7_75t_L g293 ( .A(n_244), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_223), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_243), .Y(n_295) );
OAI22xp5_ASAP7_75t_L g296 ( .A1(n_233), .A2(n_163), .B1(n_196), .B2(n_216), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_252), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_252), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_228), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_223), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_225), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_236), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_252), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_225), .Y(n_304) );
INVx3_ASAP7_75t_L g305 ( .A(n_236), .Y(n_305) );
BUFx3_ASAP7_75t_L g306 ( .A(n_250), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_225), .A2(n_196), .B1(n_176), .B2(n_163), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_273), .B(n_200), .Y(n_308) );
BUFx2_ASAP7_75t_L g309 ( .A(n_250), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_242), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_252), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_247), .A2(n_163), .B(n_213), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_237), .A2(n_216), .B1(n_200), .B2(n_195), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_271), .B(n_195), .Y(n_314) );
NAND3xp33_ASAP7_75t_L g315 ( .A(n_246), .B(n_209), .C(n_216), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_228), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_220), .Y(n_317) );
BUFx4f_ASAP7_75t_L g318 ( .A(n_245), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_238), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_239), .B(n_201), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_240), .Y(n_321) );
INVx3_ASAP7_75t_L g322 ( .A(n_251), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_220), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_224), .Y(n_324) );
OR2x2_ASAP7_75t_L g325 ( .A(n_266), .B(n_203), .Y(n_325) );
BUFx4f_ASAP7_75t_SL g326 ( .A(n_293), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_303), .Y(n_327) );
CKINVDCx14_ASAP7_75t_R g328 ( .A(n_293), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_303), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_310), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_292), .B(n_256), .Y(n_331) );
AND2x4_ASAP7_75t_L g332 ( .A(n_306), .B(n_251), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_303), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_310), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_307), .A2(n_265), .B1(n_241), .B2(n_267), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_292), .A2(n_267), .B1(n_226), .B2(n_232), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_314), .A2(n_239), .B1(n_221), .B2(n_272), .Y(n_337) );
INVx4_ASAP7_75t_L g338 ( .A(n_306), .Y(n_338) );
INVx1_ASAP7_75t_SL g339 ( .A(n_314), .Y(n_339) );
CKINVDCx20_ASAP7_75t_R g340 ( .A(n_286), .Y(n_340) );
OAI21x1_ASAP7_75t_L g341 ( .A1(n_296), .A2(n_234), .B(n_248), .Y(n_341) );
NAND2x1p5_ASAP7_75t_L g342 ( .A(n_302), .B(n_251), .Y(n_342) );
A2O1A1Ixp33_ASAP7_75t_L g343 ( .A1(n_288), .A2(n_235), .B(n_259), .C(n_260), .Y(n_343) );
NOR2xp67_ASAP7_75t_L g344 ( .A(n_306), .B(n_262), .Y(n_344) );
INVx3_ASAP7_75t_L g345 ( .A(n_302), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_303), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_308), .A2(n_239), .B1(n_221), .B2(n_272), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_303), .Y(n_348) );
OAI221xp5_ASAP7_75t_L g349 ( .A1(n_325), .A2(n_269), .B1(n_263), .B2(n_270), .C(n_249), .Y(n_349) );
INVx3_ASAP7_75t_L g350 ( .A(n_302), .Y(n_350) );
NOR2xp67_ASAP7_75t_SL g351 ( .A(n_303), .B(n_230), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_320), .A2(n_218), .B1(n_253), .B2(n_255), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_325), .A2(n_272), .B1(n_262), .B2(n_258), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_278), .Y(n_354) );
AND2x4_ASAP7_75t_L g355 ( .A(n_282), .B(n_245), .Y(n_355) );
OAI21x1_ASAP7_75t_L g356 ( .A1(n_341), .A2(n_315), .B(n_298), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_354), .Y(n_357) );
AOI22xp33_ASAP7_75t_SL g358 ( .A1(n_326), .A2(n_291), .B1(n_324), .B2(n_309), .Y(n_358) );
INVx3_ASAP7_75t_L g359 ( .A(n_342), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_330), .B(n_319), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_354), .Y(n_361) );
OAI222xp33_ASAP7_75t_L g362 ( .A1(n_349), .A2(n_299), .B1(n_316), .B2(n_309), .C1(n_282), .C2(n_313), .Y(n_362) );
INVx1_ASAP7_75t_SL g363 ( .A(n_339), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_354), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_339), .Y(n_365) );
AOI22xp33_ASAP7_75t_SL g366 ( .A1(n_338), .A2(n_253), .B1(n_287), .B2(n_199), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_331), .A2(n_321), .B1(n_319), .B2(n_287), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_331), .A2(n_321), .B1(n_262), .B2(n_300), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_330), .Y(n_369) );
AOI222xp33_ASAP7_75t_L g370 ( .A1(n_334), .A2(n_304), .B1(n_289), .B2(n_300), .C1(n_301), .C2(n_294), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_328), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_337), .A2(n_218), .B1(n_279), .B2(n_281), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_334), .B(n_278), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_340), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_353), .B(n_279), .Y(n_375) );
OAI21x1_ASAP7_75t_L g376 ( .A1(n_341), .A2(n_290), .B(n_298), .Y(n_376) );
INVx3_ASAP7_75t_L g377 ( .A(n_342), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_343), .B(n_289), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_336), .B(n_294), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_338), .B(n_281), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g381 ( .A1(n_347), .A2(n_218), .B1(n_283), .B2(n_122), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_338), .B(n_283), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_361), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_357), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_357), .B(n_349), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_364), .B(n_338), .Y(n_386) );
AOI21xp5_ASAP7_75t_L g387 ( .A1(n_361), .A2(n_352), .B(n_341), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_364), .B(n_361), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_362), .A2(n_335), .B1(n_122), .B2(n_355), .C(n_217), .Y(n_389) );
OAI221xp5_ASAP7_75t_L g390 ( .A1(n_367), .A2(n_344), .B1(n_352), .B2(n_301), .C(n_304), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_369), .Y(n_391) );
BUFx12f_ASAP7_75t_L g392 ( .A(n_371), .Y(n_392) );
OAI22xp33_ASAP7_75t_L g393 ( .A1(n_363), .A2(n_344), .B1(n_350), .B2(n_345), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_376), .Y(n_394) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_375), .A2(n_332), .B1(n_355), .B2(n_199), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_380), .B(n_199), .Y(n_396) );
OA222x2_ASAP7_75t_L g397 ( .A1(n_373), .A2(n_345), .B1(n_350), .B2(n_346), .C1(n_348), .C2(n_329), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_369), .Y(n_398) );
OAI211xp5_ASAP7_75t_L g399 ( .A1(n_358), .A2(n_208), .B(n_220), .C(n_345), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_380), .B(n_345), .Y(n_400) );
OA21x2_ASAP7_75t_L g401 ( .A1(n_356), .A2(n_327), .B(n_348), .Y(n_401) );
AOI22xp33_ASAP7_75t_SL g402 ( .A1(n_372), .A2(n_332), .B1(n_355), .B2(n_350), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_382), .B(n_350), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_373), .A2(n_332), .B1(n_333), .B2(n_346), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_365), .B(n_355), .Y(n_405) );
OAI211xp5_ASAP7_75t_L g406 ( .A1(n_366), .A2(n_208), .B(n_317), .C(n_323), .Y(n_406) );
INVx2_ASAP7_75t_SL g407 ( .A(n_382), .Y(n_407) );
AOI22xp33_ASAP7_75t_SL g408 ( .A1(n_372), .A2(n_332), .B1(n_333), .B2(n_346), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_375), .A2(n_317), .B1(n_323), .B2(n_209), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_363), .B(n_317), .Y(n_410) );
INVxp67_ASAP7_75t_SL g411 ( .A(n_360), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_360), .B(n_323), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_379), .A2(n_209), .B1(n_305), .B2(n_322), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_366), .A2(n_381), .B1(n_378), .B2(n_379), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_368), .B(n_342), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_383), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_391), .Y(n_417) );
NAND2x1_ASAP7_75t_L g418 ( .A(n_383), .B(n_359), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_388), .B(n_359), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_388), .B(n_359), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_391), .Y(n_421) );
AO21x2_ASAP7_75t_L g422 ( .A1(n_387), .A2(n_356), .B(n_376), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_383), .B(n_359), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_384), .B(n_377), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_384), .B(n_377), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_398), .Y(n_426) );
NAND3xp33_ASAP7_75t_L g427 ( .A(n_389), .B(n_370), .C(n_378), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_411), .B(n_370), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_407), .B(n_377), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_398), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_407), .A2(n_381), .B1(n_374), .B2(n_377), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_392), .B(n_362), .Y(n_432) );
OAI31xp33_ASAP7_75t_L g433 ( .A1(n_399), .A2(n_414), .A3(n_393), .B(n_386), .Y(n_433) );
INVx2_ASAP7_75t_SL g434 ( .A(n_386), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_412), .Y(n_435) );
NOR2xp67_ASAP7_75t_L g436 ( .A(n_395), .B(n_21), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_385), .B(n_376), .Y(n_437) );
AND2x2_ASAP7_75t_SL g438 ( .A(n_397), .B(n_333), .Y(n_438) );
AND2x4_ASAP7_75t_L g439 ( .A(n_400), .B(n_356), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_394), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_412), .B(n_348), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_415), .A2(n_322), .B1(n_302), .B2(n_305), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_410), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_405), .Y(n_444) );
AOI33xp33_ASAP7_75t_L g445 ( .A1(n_402), .A2(n_214), .A3(n_207), .B1(n_211), .B2(n_212), .B3(n_190), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_396), .B(n_329), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_396), .B(n_329), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_385), .B(n_327), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_404), .B(n_327), .Y(n_449) );
OR2x2_ASAP7_75t_SL g450 ( .A(n_397), .B(n_333), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_394), .Y(n_451) );
NAND3xp33_ASAP7_75t_L g452 ( .A(n_395), .B(n_185), .C(n_164), .Y(n_452) );
AND2x4_ASAP7_75t_L g453 ( .A(n_400), .B(n_333), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_394), .Y(n_454) );
INVx2_ASAP7_75t_SL g455 ( .A(n_410), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_401), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_403), .B(n_333), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_403), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_404), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_390), .Y(n_460) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_401), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_414), .B(n_401), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_417), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_444), .B(n_409), .Y(n_464) );
AND4x1_ASAP7_75t_L g465 ( .A(n_432), .B(n_392), .C(n_413), .D(n_351), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_435), .B(n_408), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_458), .B(n_22), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_421), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_440), .Y(n_469) );
BUFx3_ASAP7_75t_L g470 ( .A(n_418), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_443), .B(n_401), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_426), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_434), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_462), .B(n_406), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_430), .Y(n_475) );
NAND3xp33_ASAP7_75t_L g476 ( .A(n_433), .B(n_185), .C(n_190), .Y(n_476) );
INVx4_ASAP7_75t_L g477 ( .A(n_429), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_434), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_440), .Y(n_479) );
INVxp67_ASAP7_75t_L g480 ( .A(n_455), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_462), .B(n_194), .Y(n_481) );
AND2x4_ASAP7_75t_L g482 ( .A(n_439), .B(n_26), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_446), .B(n_194), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_455), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_428), .B(n_185), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_451), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_446), .B(n_180), .Y(n_487) );
INVx2_ASAP7_75t_SL g488 ( .A(n_418), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_424), .Y(n_489) );
NAND4xp25_ASAP7_75t_SL g490 ( .A(n_431), .B(n_27), .C(n_31), .D(n_32), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_447), .B(n_180), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_447), .B(n_164), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_437), .B(n_214), .Y(n_493) );
INVx1_ASAP7_75t_SL g494 ( .A(n_419), .Y(n_494) );
OAI31xp33_ASAP7_75t_L g495 ( .A1(n_427), .A2(n_322), .A3(n_305), .B(n_245), .Y(n_495) );
OAI322xp33_ASAP7_75t_L g496 ( .A1(n_460), .A2(n_211), .A3(n_212), .B1(n_254), .B2(n_257), .C1(n_227), .C2(n_268), .Y(n_496) );
AOI21xp33_ASAP7_75t_L g497 ( .A1(n_437), .A2(n_351), .B(n_295), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_424), .Y(n_498) );
INVx3_ASAP7_75t_L g499 ( .A(n_461), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_439), .B(n_39), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_439), .B(n_45), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_419), .B(n_48), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_425), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_459), .B(n_51), .Y(n_504) );
NOR2x1_ASAP7_75t_SL g505 ( .A(n_429), .B(n_280), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_425), .B(n_52), .Y(n_506) );
INVx1_ASAP7_75t_SL g507 ( .A(n_420), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_420), .B(n_53), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_416), .B(n_54), .Y(n_509) );
OAI21xp5_ASAP7_75t_SL g510 ( .A1(n_450), .A2(n_322), .B(n_305), .Y(n_510) );
AND2x4_ASAP7_75t_L g511 ( .A(n_456), .B(n_56), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_451), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_457), .B(n_64), .Y(n_513) );
INVxp67_ASAP7_75t_L g514 ( .A(n_423), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_416), .B(n_67), .Y(n_515) );
INVx1_ASAP7_75t_SL g516 ( .A(n_423), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_454), .Y(n_517) );
NAND2x1_ASAP7_75t_L g518 ( .A(n_477), .B(n_456), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_494), .B(n_457), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_473), .B(n_448), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_478), .B(n_441), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_507), .B(n_449), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_474), .B(n_456), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_474), .B(n_461), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_489), .B(n_461), .Y(n_525) );
OAI31xp33_ASAP7_75t_L g526 ( .A1(n_510), .A2(n_452), .A3(n_450), .B(n_449), .Y(n_526) );
NOR3xp33_ASAP7_75t_L g527 ( .A(n_490), .B(n_445), .C(n_436), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_468), .Y(n_528) );
AOI21x1_ASAP7_75t_SL g529 ( .A1(n_485), .A2(n_453), .B(n_438), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_498), .B(n_461), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_503), .B(n_461), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_481), .B(n_454), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_484), .B(n_453), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_466), .A2(n_438), .B1(n_453), .B2(n_442), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_516), .B(n_422), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_469), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_514), .B(n_422), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_480), .B(n_422), .Y(n_538) );
HB1xp67_ASAP7_75t_SL g539 ( .A(n_477), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_468), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_481), .B(n_445), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_513), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_477), .B(n_70), .Y(n_543) );
AND4x1_ASAP7_75t_L g544 ( .A(n_495), .B(n_72), .C(n_74), .D(n_312), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_472), .Y(n_545) );
NAND2x1p5_ASAP7_75t_L g546 ( .A(n_482), .B(n_285), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_472), .B(n_280), .Y(n_547) );
OR2x6_ASAP7_75t_L g548 ( .A(n_482), .B(n_285), .Y(n_548) );
AND3x2_ASAP7_75t_L g549 ( .A(n_500), .B(n_285), .C(n_280), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_463), .B(n_297), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_471), .B(n_290), .Y(n_551) );
AOI211x1_ASAP7_75t_SL g552 ( .A1(n_476), .A2(n_298), .B(n_290), .C(n_295), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_517), .B(n_297), .Y(n_553) );
INVx3_ASAP7_75t_L g554 ( .A(n_470), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_475), .B(n_297), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_471), .Y(n_556) );
AND2x2_ASAP7_75t_SL g557 ( .A(n_482), .B(n_318), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_500), .B(n_295), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_464), .B(n_311), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_517), .Y(n_560) );
NAND3xp33_ASAP7_75t_L g561 ( .A(n_465), .B(n_261), .C(n_311), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_493), .B(n_284), .Y(n_562) );
NAND2x1p5_ASAP7_75t_L g563 ( .A(n_511), .B(n_285), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_493), .B(n_284), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_501), .B(n_261), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_483), .B(n_261), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_483), .B(n_261), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_539), .A2(n_504), .B1(n_501), .B2(n_506), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_528), .Y(n_569) );
OAI32xp33_ASAP7_75t_L g570 ( .A1(n_527), .A2(n_504), .A3(n_470), .B1(n_502), .B2(n_508), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_556), .B(n_486), .Y(n_571) );
AOI322xp5_ASAP7_75t_L g572 ( .A1(n_523), .A2(n_467), .A3(n_502), .B1(n_508), .B2(n_513), .C1(n_511), .C2(n_488), .Y(n_572) );
INVx1_ASAP7_75t_SL g573 ( .A(n_519), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_523), .B(n_499), .Y(n_574) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_526), .B(n_488), .Y(n_575) );
INVxp67_ASAP7_75t_L g576 ( .A(n_538), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_540), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_537), .B(n_479), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_524), .B(n_499), .Y(n_579) );
OAI22xp33_ASAP7_75t_L g580 ( .A1(n_548), .A2(n_515), .B1(n_509), .B2(n_511), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_524), .B(n_469), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_545), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_522), .B(n_520), .Y(n_583) );
OAI221xp5_ASAP7_75t_L g584 ( .A1(n_534), .A2(n_499), .B1(n_515), .B2(n_509), .C(n_479), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_521), .B(n_512), .Y(n_585) );
OAI22xp33_ASAP7_75t_L g586 ( .A1(n_548), .A2(n_512), .B1(n_486), .B2(n_505), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_538), .B(n_492), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_542), .B(n_505), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_536), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_560), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_525), .B(n_492), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_536), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_525), .Y(n_593) );
OR2x6_ASAP7_75t_L g594 ( .A(n_518), .B(n_491), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_530), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_530), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_533), .B(n_491), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_531), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_531), .B(n_487), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_532), .B(n_487), .Y(n_600) );
NAND2x1_ASAP7_75t_L g601 ( .A(n_554), .B(n_497), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_541), .B(n_496), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_532), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_548), .A2(n_318), .B1(n_254), .B2(n_274), .Y(n_604) );
NOR3xp33_ASAP7_75t_L g605 ( .A(n_527), .B(n_247), .C(n_277), .Y(n_605) );
OAI21xp5_ASAP7_75t_SL g606 ( .A1(n_549), .A2(n_274), .B(n_277), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_535), .Y(n_607) );
OAI22xp33_ASAP7_75t_SL g608 ( .A1(n_554), .A2(n_318), .B1(n_274), .B2(n_275), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_554), .B(n_227), .Y(n_609) );
OAI22xp33_ASAP7_75t_L g610 ( .A1(n_546), .A2(n_318), .B1(n_230), .B2(n_229), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_551), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_547), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_541), .A2(n_276), .B1(n_257), .B2(n_268), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_558), .B(n_275), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_547), .Y(n_615) );
XOR2x2_ASAP7_75t_L g616 ( .A(n_557), .B(n_229), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_555), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_550), .Y(n_618) );
OAI22xp33_ASAP7_75t_L g619 ( .A1(n_546), .A2(n_275), .B1(n_277), .B2(n_563), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_557), .A2(n_549), .B1(n_550), .B2(n_566), .Y(n_620) );
NOR3xp33_ASAP7_75t_L g621 ( .A(n_561), .B(n_567), .C(n_543), .Y(n_621) );
AOI211xp5_ASAP7_75t_L g622 ( .A1(n_565), .A2(n_559), .B(n_529), .C(n_562), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_553), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_553), .B(n_564), .Y(n_624) );
O2A1O1Ixp5_ASAP7_75t_L g625 ( .A1(n_575), .A2(n_570), .B(n_601), .C(n_602), .Y(n_625) );
OAI21xp5_ASAP7_75t_L g626 ( .A1(n_575), .A2(n_605), .B(n_621), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_576), .B(n_587), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_583), .Y(n_628) );
OAI22xp5_ASAP7_75t_SL g629 ( .A1(n_594), .A2(n_620), .B1(n_568), .B2(n_588), .Y(n_629) );
XNOR2xp5_ASAP7_75t_L g630 ( .A(n_600), .B(n_573), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g631 ( .A1(n_576), .A2(n_618), .B1(n_605), .B2(n_584), .C(n_598), .Y(n_631) );
OAI22xp33_ASAP7_75t_L g632 ( .A1(n_594), .A2(n_586), .B1(n_606), .B2(n_588), .Y(n_632) );
XNOR2xp5_ASAP7_75t_L g633 ( .A(n_591), .B(n_616), .Y(n_633) );
AOI211xp5_ASAP7_75t_SL g634 ( .A1(n_621), .A2(n_608), .B(n_619), .C(n_586), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_585), .Y(n_635) );
O2A1O1Ixp33_ASAP7_75t_L g636 ( .A1(n_619), .A2(n_580), .B(n_594), .C(n_622), .Y(n_636) );
XNOR2xp5_ASAP7_75t_L g637 ( .A(n_597), .B(n_620), .Y(n_637) );
OAI221xp5_ASAP7_75t_L g638 ( .A1(n_629), .A2(n_572), .B1(n_607), .B2(n_613), .C(n_578), .Y(n_638) );
NAND4xp25_ASAP7_75t_L g639 ( .A(n_634), .B(n_636), .C(n_625), .D(n_626), .Y(n_639) );
A2O1A1Ixp33_ASAP7_75t_L g640 ( .A1(n_634), .A2(n_599), .B(n_603), .C(n_596), .Y(n_640) );
AOI221x1_ASAP7_75t_L g641 ( .A1(n_627), .A2(n_577), .B1(n_582), .B2(n_569), .C(n_590), .Y(n_641) );
OAI311xp33_ASAP7_75t_L g642 ( .A1(n_631), .A2(n_624), .A3(n_617), .B1(n_571), .C1(n_581), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_632), .A2(n_593), .B1(n_599), .B2(n_580), .C(n_595), .Y(n_643) );
AOI22xp33_ASAP7_75t_SL g644 ( .A1(n_628), .A2(n_574), .B1(n_563), .B2(n_579), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_638), .A2(n_637), .B1(n_630), .B2(n_633), .Y(n_645) );
OA22x2_ASAP7_75t_L g646 ( .A1(n_639), .A2(n_635), .B1(n_595), .B2(n_611), .Y(n_646) );
OAI211xp5_ASAP7_75t_SL g647 ( .A1(n_640), .A2(n_552), .B(n_610), .C(n_604), .Y(n_647) );
AND4x1_ASAP7_75t_L g648 ( .A(n_643), .B(n_609), .C(n_614), .D(n_615), .Y(n_648) );
AOI22xp33_ASAP7_75t_SL g649 ( .A1(n_645), .A2(n_642), .B1(n_641), .B2(n_644), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_646), .B(n_610), .Y(n_650) );
NOR3xp33_ASAP7_75t_L g651 ( .A(n_647), .B(n_589), .C(n_592), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_650), .Y(n_652) );
XOR2xp5_ASAP7_75t_L g653 ( .A(n_649), .B(n_648), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_652), .Y(n_654) );
BUFx2_ASAP7_75t_L g655 ( .A(n_654), .Y(n_655) );
OAI22xp33_ASAP7_75t_L g656 ( .A1(n_655), .A2(n_653), .B1(n_651), .B2(n_612), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g657 ( .A1(n_656), .A2(n_623), .B(n_544), .Y(n_657) );
endmodule