module real_aes_5392_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_693;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_298;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_602;
wire n_402;
wire n_552;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_898;
wire n_115;
wire n_604;
wire n_110;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_756;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_899;
wire n_526;
wire n_637;
wire n_155;
wire n_653;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_922;
wire n_679;
wire n_520;
wire n_482;
wire n_633;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_639;
wire n_151;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_237;
wire n_797;
wire n_862;
NAND2xp5_ASAP7_75t_L g570 ( .A(n_0), .B(n_162), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_1), .Y(n_583) );
O2A1O1Ixp33_ASAP7_75t_SL g637 ( .A1(n_2), .A2(n_139), .B(n_638), .C(n_639), .Y(n_637) );
OAI22xp33_ASAP7_75t_L g575 ( .A1(n_3), .A2(n_78), .B1(n_133), .B2(n_136), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g227 ( .A1(n_4), .A2(n_28), .B1(n_142), .B2(n_228), .Y(n_227) );
INVxp67_ASAP7_75t_L g108 ( .A(n_5), .Y(n_108) );
INVx1_ASAP7_75t_L g548 ( .A(n_5), .Y(n_548) );
INVx1_ASAP7_75t_L g897 ( .A(n_5), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g215 ( .A1(n_6), .A2(n_86), .B1(n_216), .B2(n_217), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g600 ( .A(n_7), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_8), .A2(n_65), .B1(n_136), .B2(n_144), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g246 ( .A1(n_9), .A2(n_29), .B1(n_247), .B2(n_248), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g666 ( .A(n_10), .Y(n_666) );
INVx2_ASAP7_75t_L g183 ( .A(n_11), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_12), .A2(n_59), .B1(n_133), .B2(n_176), .Y(n_628) );
OA21x2_ASAP7_75t_L g127 ( .A1(n_13), .A2(n_64), .B(n_128), .Y(n_127) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_13), .A2(n_64), .B(n_128), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_14), .B(n_105), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g314 ( .A(n_15), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_SL g180 ( .A(n_16), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_17), .B(n_318), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g596 ( .A(n_18), .Y(n_596) );
BUFx3_ASAP7_75t_L g103 ( .A(n_19), .Y(n_103) );
O2A1O1Ixp33_ASAP7_75t_L g642 ( .A1(n_20), .A2(n_148), .B(n_202), .C(n_643), .Y(n_642) );
OAI22xp33_ASAP7_75t_SL g573 ( .A1(n_21), .A2(n_44), .B1(n_133), .B2(n_179), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_22), .A2(n_27), .B1(n_179), .B2(n_220), .Y(n_562) );
O2A1O1Ixp5_ASAP7_75t_L g188 ( .A1(n_23), .A2(n_189), .B(n_192), .C(n_194), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_24), .B(n_233), .Y(n_311) );
O2A1O1Ixp5_ASAP7_75t_L g611 ( .A1(n_25), .A2(n_139), .B(n_170), .C(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g113 ( .A(n_26), .Y(n_113) );
AND2x2_ASAP7_75t_L g921 ( .A(n_30), .B(n_922), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_31), .B(n_212), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g613 ( .A(n_32), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g231 ( .A1(n_33), .A2(n_37), .B1(n_219), .B2(n_232), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g218 ( .A1(n_34), .A2(n_63), .B1(n_135), .B2(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g310 ( .A(n_35), .B(n_229), .Y(n_310) );
INVx2_ASAP7_75t_L g125 ( .A(n_36), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g640 ( .A(n_38), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_39), .B(n_205), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_40), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_L g174 ( .A1(n_41), .A2(n_148), .B(n_175), .C(n_177), .Y(n_174) );
INVx1_ASAP7_75t_L g277 ( .A(n_42), .Y(n_277) );
INVx2_ASAP7_75t_L g203 ( .A(n_43), .Y(n_203) );
INVx1_ASAP7_75t_L g128 ( .A(n_45), .Y(n_128) );
AND2x4_ASAP7_75t_L g150 ( .A(n_46), .B(n_151), .Y(n_150) );
AND2x4_ASAP7_75t_L g207 ( .A(n_46), .B(n_151), .Y(n_207) );
INVx2_ASAP7_75t_L g138 ( .A(n_47), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_48), .B(n_212), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_48), .A2(n_62), .B1(n_212), .B2(n_679), .Y(n_678) );
INVxp67_ASAP7_75t_SL g693 ( .A(n_48), .Y(n_693) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_49), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g581 ( .A(n_50), .Y(n_581) );
O2A1O1Ixp33_ASAP7_75t_L g597 ( .A1(n_51), .A2(n_139), .B(n_598), .C(n_599), .Y(n_597) );
CKINVDCx5p33_ASAP7_75t_R g619 ( .A(n_52), .Y(n_619) );
INVx2_ASAP7_75t_L g671 ( .A(n_53), .Y(n_671) );
CKINVDCx5p33_ASAP7_75t_R g580 ( .A(n_54), .Y(n_580) );
INVx1_ASAP7_75t_SL g193 ( .A(n_55), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g99 ( .A1(n_56), .A2(n_100), .B1(n_916), .B2(n_923), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_57), .B(n_318), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_58), .A2(n_75), .B1(n_143), .B2(n_564), .Y(n_563) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_60), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g584 ( .A(n_61), .Y(n_584) );
NAND2xp33_ASAP7_75t_R g631 ( .A(n_62), .B(n_127), .Y(n_631) );
INVx1_ASAP7_75t_L g911 ( .A(n_66), .Y(n_911) );
O2A1O1Ixp33_ASAP7_75t_L g141 ( .A1(n_67), .A2(n_142), .B(n_146), .C(n_148), .Y(n_141) );
OR2x6_ASAP7_75t_L g110 ( .A(n_68), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g273 ( .A(n_69), .Y(n_273) );
CKINVDCx16_ASAP7_75t_R g281 ( .A(n_70), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g670 ( .A(n_71), .Y(n_670) );
CKINVDCx5p33_ASAP7_75t_R g667 ( .A(n_72), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_73), .B(n_247), .Y(n_316) );
NOR2xp67_ASAP7_75t_L g169 ( .A(n_74), .B(n_170), .Y(n_169) );
O2A1O1Ixp33_ASAP7_75t_L g130 ( .A1(n_76), .A2(n_131), .B(n_134), .C(n_139), .Y(n_130) );
O2A1O1Ixp33_ASAP7_75t_L g328 ( .A1(n_76), .A2(n_131), .B(n_134), .C(n_139), .Y(n_328) );
INVx1_ASAP7_75t_L g112 ( .A(n_77), .Y(n_112) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_79), .A2(n_90), .B1(n_251), .B2(n_253), .Y(n_250) );
INVx1_ASAP7_75t_L g922 ( .A(n_80), .Y(n_922) );
BUFx5_ASAP7_75t_L g133 ( .A(n_81), .Y(n_133) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_81), .Y(n_137) );
INVx1_ASAP7_75t_L g145 ( .A(n_81), .Y(n_145) );
INVx2_ASAP7_75t_L g647 ( .A(n_82), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_83), .B(n_284), .Y(n_283) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_84), .Y(n_115) );
INVx2_ASAP7_75t_L g602 ( .A(n_85), .Y(n_602) );
CKINVDCx5p33_ASAP7_75t_R g644 ( .A(n_87), .Y(n_644) );
INVx2_ASAP7_75t_SL g151 ( .A(n_88), .Y(n_151) );
INVx1_ASAP7_75t_L g617 ( .A(n_89), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_91), .B(n_127), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g903 ( .A(n_92), .Y(n_903) );
INVx1_ASAP7_75t_SL g239 ( .A(n_93), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_94), .B(n_152), .Y(n_208) );
INVx2_ASAP7_75t_L g621 ( .A(n_95), .Y(n_621) );
AND2x2_ASAP7_75t_L g256 ( .A(n_96), .B(n_257), .Y(n_256) );
OAI21xp33_ASAP7_75t_SL g594 ( .A1(n_97), .A2(n_133), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_SL g201 ( .A(n_98), .Y(n_201) );
OA22x2_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_114), .B1(n_907), .B2(n_913), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_102), .B(n_104), .Y(n_101) );
BUFx3_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
CKINVDCx6p67_ASAP7_75t_R g915 ( .A(n_103), .Y(n_915) );
OAI21xp5_ASAP7_75t_L g907 ( .A1(n_104), .A2(n_908), .B(n_909), .Y(n_907) );
INVx2_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx3_ASAP7_75t_L g908 ( .A(n_106), .Y(n_908) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
OR2x6_ASAP7_75t_L g547 ( .A(n_109), .B(n_548), .Y(n_547) );
INVx8_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g896 ( .A(n_110), .B(n_897), .Y(n_896) );
OR2x6_ASAP7_75t_L g906 ( .A(n_110), .B(n_897), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
OAI21x1_ASAP7_75t_SL g114 ( .A1(n_115), .A2(n_116), .B(n_898), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g898 ( .A1(n_115), .A2(n_899), .B(n_902), .Y(n_898) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI22x1_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_546), .B1(n_549), .B2(n_893), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI22x1_ASAP7_75t_L g899 ( .A1(n_119), .A2(n_546), .B1(n_550), .B2(n_900), .Y(n_899) );
AND2x4_ASAP7_75t_L g119 ( .A(n_120), .B(n_419), .Y(n_119) );
NOR3xp33_ASAP7_75t_SL g120 ( .A(n_121), .B(n_350), .C(n_389), .Y(n_120) );
OAI211xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_154), .B(n_240), .C(n_333), .Y(n_121) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_122), .A2(n_425), .B1(n_426), .B2(n_428), .Y(n_424) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
NOR2x1_ASAP7_75t_L g258 ( .A(n_123), .B(n_259), .Y(n_258) );
AND2x4_ASAP7_75t_L g295 ( .A(n_123), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_123), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g412 ( .A(n_123), .Y(n_412) );
AND2x2_ASAP7_75t_L g454 ( .A(n_123), .B(n_243), .Y(n_454) );
OR2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_129), .Y(n_123) );
INVxp67_ASAP7_75t_SL g330 ( .A(n_124), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_125), .B(n_126), .Y(n_124) );
INVx1_ASAP7_75t_L g261 ( .A(n_126), .Y(n_261) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g153 ( .A(n_127), .Y(n_153) );
BUFx3_ASAP7_75t_L g257 ( .A(n_127), .Y(n_257) );
INVx1_ASAP7_75t_L g592 ( .A(n_127), .Y(n_592) );
INVx1_ASAP7_75t_L g622 ( .A(n_127), .Y(n_622) );
NOR4xp25_ASAP7_75t_L g129 ( .A(n_130), .B(n_141), .C(n_149), .D(n_152), .Y(n_129) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NAND2xp33_ASAP7_75t_L g167 ( .A(n_133), .B(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g216 ( .A(n_133), .Y(n_216) );
INVx2_ASAP7_75t_L g233 ( .A(n_133), .Y(n_233) );
INVx2_ASAP7_75t_L g247 ( .A(n_133), .Y(n_247) );
INVx2_ASAP7_75t_L g253 ( .A(n_133), .Y(n_253) );
AOI22xp33_ASAP7_75t_SL g579 ( .A1(n_133), .A2(n_179), .B1(n_580), .B2(n_581), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_133), .A2(n_176), .B1(n_583), .B2(n_584), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_133), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_133), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_133), .B(n_619), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g665 ( .A1(n_133), .A2(n_179), .B1(n_666), .B2(n_667), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_138), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_135), .B(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g200 ( .A(n_135), .Y(n_200) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g284 ( .A(n_136), .Y(n_284) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx3_ASAP7_75t_L g171 ( .A(n_137), .Y(n_171) );
INVx2_ASAP7_75t_L g176 ( .A(n_137), .Y(n_176) );
INVx6_ASAP7_75t_L g179 ( .A(n_137), .Y(n_179) );
INVx1_ASAP7_75t_L g172 ( .A(n_139), .Y(n_172) );
INVx2_ASAP7_75t_SL g221 ( .A(n_139), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_139), .B(n_273), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_139), .B(n_277), .Y(n_276) );
OAI221xp5_ASAP7_75t_L g578 ( .A1(n_139), .A2(n_148), .B1(n_207), .B2(n_579), .C(n_582), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_139), .A2(n_285), .B1(n_628), .B2(n_629), .Y(n_627) );
INVx1_ASAP7_75t_L g672 ( .A(n_139), .Y(n_672) );
OAI22xp33_ASAP7_75t_L g691 ( .A1(n_139), .A2(n_285), .B1(n_665), .B2(n_669), .Y(n_691) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx3_ASAP7_75t_L g148 ( .A(n_140), .Y(n_148) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_140), .Y(n_195) );
INVxp67_ASAP7_75t_L g198 ( .A(n_140), .Y(n_198) );
INVx4_ASAP7_75t_L g285 ( .A(n_140), .Y(n_285) );
INVx1_ASAP7_75t_L g565 ( .A(n_140), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_140), .B(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_140), .B(n_617), .Y(n_616) );
INVxp67_ASAP7_75t_SL g329 ( .A(n_141), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_142), .B(n_193), .Y(n_192) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g638 ( .A(n_143), .Y(n_638) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g220 ( .A(n_145), .Y(n_220) );
INVx3_ASAP7_75t_L g234 ( .A(n_148), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_148), .A2(n_575), .B(n_576), .Y(n_574) );
NOR2x1_ASAP7_75t_SL g159 ( .A(n_149), .B(n_160), .Y(n_159) );
NOR3xp33_ASAP7_75t_L g610 ( .A(n_149), .B(n_611), .C(n_614), .Y(n_610) );
NOR2xp33_ASAP7_75t_SL g645 ( .A(n_149), .B(n_162), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g663 ( .A1(n_149), .A2(n_312), .B1(n_664), .B2(n_668), .C(n_672), .Y(n_663) );
INVx4_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_150), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g591 ( .A(n_150), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_153), .B(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g679 ( .A(n_153), .Y(n_679) );
NAND2x1_ASAP7_75t_L g154 ( .A(n_155), .B(n_184), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g355 ( .A(n_157), .Y(n_355) );
AND2x2_ASAP7_75t_L g388 ( .A(n_157), .B(n_347), .Y(n_388) );
AND2x2_ASAP7_75t_L g416 ( .A(n_157), .B(n_305), .Y(n_416) );
AND2x2_ASAP7_75t_L g448 ( .A(n_157), .B(n_434), .Y(n_448) );
INVx1_ASAP7_75t_L g536 ( .A(n_157), .Y(n_536) );
OR2x2_ASAP7_75t_L g541 ( .A(n_157), .B(n_534), .Y(n_541) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
OR2x2_ASAP7_75t_L g332 ( .A(n_158), .B(n_268), .Y(n_332) );
OR2x2_ASAP7_75t_L g343 ( .A(n_158), .B(n_303), .Y(n_343) );
AND2x4_ASAP7_75t_L g363 ( .A(n_158), .B(n_303), .Y(n_363) );
INVx1_ASAP7_75t_L g371 ( .A(n_158), .Y(n_371) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_158), .Y(n_458) );
AND2x2_ASAP7_75t_L g473 ( .A(n_158), .B(n_268), .Y(n_473) );
AO31x2_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_165), .A3(n_173), .B(n_181), .Y(n_158) );
OA21x2_ASAP7_75t_L g577 ( .A1(n_160), .A2(n_578), .B(n_585), .Y(n_577) );
OA21x2_ASAP7_75t_L g654 ( .A1(n_160), .A2(n_578), .B(n_585), .Y(n_654) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
OR2x2_ASAP7_75t_L g692 ( .A(n_161), .B(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g212 ( .A(n_163), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_163), .B(n_207), .Y(n_576) );
NOR2xp33_ASAP7_75t_SL g646 ( .A(n_163), .B(n_647), .Y(n_646) );
INVx4_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g182 ( .A(n_164), .Y(n_182) );
BUFx3_ASAP7_75t_L g205 ( .A(n_164), .Y(n_205) );
OAI21xp5_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_169), .B(n_172), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g217 ( .A(n_171), .Y(n_217) );
INVx2_ASAP7_75t_L g229 ( .A(n_171), .Y(n_229) );
INVx1_ASAP7_75t_L g598 ( .A(n_171), .Y(n_598) );
INVx1_ASAP7_75t_L g615 ( .A(n_171), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g313 ( .A1(n_172), .A2(n_314), .B(n_316), .Y(n_313) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVxp67_ASAP7_75t_SL g175 ( .A(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g202 ( .A(n_176), .Y(n_202) );
INVx2_ASAP7_75t_L g248 ( .A(n_176), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_176), .A2(n_220), .B1(n_670), .B2(n_671), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_178), .B(n_180), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_178), .B(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g191 ( .A(n_179), .Y(n_191) );
INVx1_ASAP7_75t_L g279 ( .A(n_179), .Y(n_279) );
INVx1_ASAP7_75t_L g315 ( .A(n_179), .Y(n_315) );
INVx2_ASAP7_75t_SL g564 ( .A(n_179), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
BUFx3_ASAP7_75t_L g288 ( .A(n_182), .Y(n_288) );
INVx3_ASAP7_75t_L g318 ( .A(n_182), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_182), .B(n_602), .Y(n_601) );
AOI322xp5_ASAP7_75t_L g403 ( .A1(n_184), .A2(n_391), .A3(n_404), .B1(n_405), .B2(n_407), .C1(n_409), .C2(n_414), .Y(n_403) );
AND2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_209), .Y(n_184) );
INVx1_ASAP7_75t_L g289 ( .A(n_185), .Y(n_289) );
BUFx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g341 ( .A(n_186), .B(n_306), .Y(n_341) );
INVx2_ASAP7_75t_SL g348 ( .A(n_186), .Y(n_348) );
AND2x2_ASAP7_75t_L g418 ( .A(n_186), .B(n_303), .Y(n_418) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g300 ( .A(n_187), .Y(n_300) );
INVx3_ASAP7_75t_L g435 ( .A(n_187), .Y(n_435) );
OA21x2_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_196), .B(n_208), .Y(n_187) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_194), .B(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_194), .B(n_250), .Y(n_249) );
INVx4_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
OA22x2_ASAP7_75t_L g561 ( .A1(n_195), .A2(n_562), .B1(n_563), .B2(n_565), .Y(n_561) );
OAI21xp5_ASAP7_75t_SL g196 ( .A1(n_197), .A2(n_199), .B(n_204), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g214 ( .A1(n_197), .A2(n_215), .B1(n_218), .B2(n_221), .Y(n_214) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B1(n_202), .B2(n_203), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
INVx3_ASAP7_75t_L g255 ( .A(n_205), .Y(n_255) );
NOR2xp67_ASAP7_75t_L g630 ( .A(n_206), .B(n_318), .Y(n_630) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx3_ASAP7_75t_L g237 ( .A(n_207), .Y(n_237) );
AND2x2_ASAP7_75t_L g254 ( .A(n_207), .B(n_255), .Y(n_254) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_207), .Y(n_263) );
AND2x6_ASAP7_75t_SL g349 ( .A(n_209), .B(n_242), .Y(n_349) );
AND2x2_ASAP7_75t_L g480 ( .A(n_209), .B(n_443), .Y(n_480) );
AND2x2_ASAP7_75t_L g491 ( .A(n_209), .B(n_461), .Y(n_491) );
AND2x4_ASAP7_75t_L g538 ( .A(n_209), .B(n_295), .Y(n_538) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_224), .Y(n_209) );
OR2x2_ASAP7_75t_L g292 ( .A(n_210), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g322 ( .A(n_210), .Y(n_322) );
AOI21x1_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_213), .B(n_222), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_211), .B(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_214), .B(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g252 ( .A(n_220), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_220), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_220), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
OA21x2_ASAP7_75t_L g260 ( .A1(n_223), .A2(n_261), .B(n_262), .Y(n_260) );
NOR2x1_ASAP7_75t_L g323 ( .A(n_224), .B(n_324), .Y(n_323) );
NAND2x1_ASAP7_75t_L g366 ( .A(n_224), .B(n_297), .Y(n_366) );
INVx1_ASAP7_75t_L g487 ( .A(n_224), .Y(n_487) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g294 ( .A(n_225), .Y(n_294) );
AOI21x1_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_230), .B(n_238), .Y(n_225) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_234), .B(n_235), .Y(n_230) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_234), .B(n_246), .Y(n_245) );
OAI21x1_ASAP7_75t_L g308 ( .A1(n_236), .A2(n_309), .B(n_313), .Y(n_308) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
OAI21x1_ASAP7_75t_L g286 ( .A1(n_237), .A2(n_274), .B(n_287), .Y(n_286) );
AOI222xp33_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_264), .B1(n_290), .B2(n_298), .C1(n_319), .C2(n_331), .Y(n_240) );
AND2x2_ASAP7_75t_L g486 ( .A(n_241), .B(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_258), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_242), .B(n_323), .Y(n_379) );
INVx1_ASAP7_75t_L g522 ( .A(n_242), .Y(n_522) );
BUFx3_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_SL g297 ( .A(n_244), .Y(n_297) );
AO31x2_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_249), .A3(n_254), .B(n_256), .Y(n_244) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g271 ( .A(n_253), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_255), .B(n_263), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g699 ( .A1(n_255), .A2(n_700), .B(n_701), .Y(n_699) );
INVx1_ASAP7_75t_L g560 ( .A(n_257), .Y(n_560) );
INVx1_ASAP7_75t_L g367 ( .A(n_258), .Y(n_367) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_260), .Y(n_387) );
AND2x2_ASAP7_75t_L g438 ( .A(n_260), .B(n_293), .Y(n_438) );
OAI21x1_ASAP7_75t_L g357 ( .A1(n_261), .A2(n_308), .B(n_317), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_263), .B(n_560), .Y(n_690) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_289), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g440 ( .A(n_267), .B(n_441), .Y(n_440) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OAI21xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_280), .B(n_286), .Y(n_268) );
OAI21x1_ASAP7_75t_L g304 ( .A1(n_269), .A2(n_280), .B(n_286), .Y(n_304) );
NAND3x1_ASAP7_75t_L g269 ( .A(n_270), .B(n_274), .C(n_275), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
INVx1_ASAP7_75t_L g282 ( .A(n_278), .Y(n_282) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
O2A1O1Ixp5_ASAP7_75t_SL g280 ( .A1(n_281), .A2(n_282), .B(n_283), .C(n_285), .Y(n_280) );
INVx2_ASAP7_75t_L g312 ( .A(n_285), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_285), .A2(n_615), .B1(n_616), .B2(n_618), .Y(n_614) );
OAI21x1_ASAP7_75t_L g307 ( .A1(n_287), .A2(n_308), .B(n_317), .Y(n_307) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AO21x2_ASAP7_75t_L g609 ( .A1(n_288), .A2(n_610), .B(n_620), .Y(n_609) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_288), .B(n_663), .Y(n_662) );
AND2x4_ASAP7_75t_L g290 ( .A(n_291), .B(n_295), .Y(n_290) );
AND2x4_ASAP7_75t_L g460 ( .A(n_291), .B(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_292), .A2(n_516), .B1(n_519), .B2(n_520), .Y(n_515) );
AND2x4_ASAP7_75t_L g376 ( .A(n_293), .B(n_324), .Y(n_376) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g337 ( .A(n_294), .Y(n_337) );
AND2x2_ASAP7_75t_L g405 ( .A(n_295), .B(n_406), .Y(n_405) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_295), .Y(n_427) );
INVx2_ASAP7_75t_SL g439 ( .A(n_295), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_295), .B(n_466), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_296), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g361 ( .A(n_296), .Y(n_361) );
BUFx2_ASAP7_75t_SL g443 ( .A(n_296), .Y(n_443) );
AND2x2_ASAP7_75t_L g461 ( .A(n_296), .B(n_324), .Y(n_461) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_299), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g478 ( .A(n_299), .B(n_356), .Y(n_478) );
AND2x2_ASAP7_75t_L g500 ( .A(n_299), .B(n_363), .Y(n_500) );
INVx2_ASAP7_75t_R g299 ( .A(n_300), .Y(n_299) );
BUFx2_ASAP7_75t_L g429 ( .A(n_300), .Y(n_429) );
INVx1_ASAP7_75t_L g485 ( .A(n_301), .Y(n_485) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g503 ( .A(n_302), .B(n_370), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g347 ( .A(n_304), .B(n_306), .Y(n_347) );
AND2x2_ASAP7_75t_L g356 ( .A(n_304), .B(n_357), .Y(n_356) );
BUFx2_ASAP7_75t_SL g372 ( .A(n_305), .Y(n_372) );
INVx1_ASAP7_75t_L g396 ( .A(n_305), .Y(n_396) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_305), .Y(n_450) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g433 ( .A(n_306), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_311), .B(n_312), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g593 ( .A1(n_312), .A2(n_594), .B(n_597), .Y(n_593) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_323), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g374 ( .A(n_321), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g358 ( .A(n_322), .B(n_337), .Y(n_358) );
OA21x2_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_326), .B(n_330), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_331), .B(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g475 ( .A(n_332), .B(n_476), .Y(n_475) );
OR2x2_ASAP7_75t_L g498 ( .A(n_332), .B(n_348), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_338), .B1(n_344), .B2(n_349), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_337), .Y(n_406) );
INVx1_ASAP7_75t_L g466 ( .A(n_337), .Y(n_466) );
INVxp67_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
NAND2x1p5_ASAP7_75t_L g339 ( .A(n_340), .B(n_342), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_340), .B(n_382), .Y(n_381) );
BUFx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2x1_ASAP7_75t_SL g457 ( .A(n_341), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g476 ( .A(n_341), .Y(n_476) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVxp67_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_345), .A2(n_456), .B(n_459), .Y(n_455) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
AND2x2_ASAP7_75t_L g514 ( .A(n_347), .B(n_472), .Y(n_514) );
INVx2_ASAP7_75t_L g534 ( .A(n_347), .Y(n_534) );
AND2x2_ASAP7_75t_L g393 ( .A(n_348), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g408 ( .A(n_348), .Y(n_408) );
INVx2_ASAP7_75t_L g472 ( .A(n_348), .Y(n_472) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_348), .Y(n_543) );
OAI311xp33_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_358), .A3(n_359), .B1(n_362), .C1(n_377), .Y(n_350) );
INVxp67_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x4_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
AND2x4_ASAP7_75t_L g391 ( .A(n_356), .B(n_371), .Y(n_391) );
NAND2xp5_ASAP7_75t_SL g428 ( .A(n_356), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g447 ( .A(n_356), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g508 ( .A(n_356), .Y(n_508) );
AND2x2_ASAP7_75t_L g495 ( .A(n_357), .B(n_435), .Y(n_495) );
AND2x2_ASAP7_75t_L g513 ( .A(n_358), .B(n_361), .Y(n_513) );
INVx1_ASAP7_75t_L g523 ( .A(n_358), .Y(n_523) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g404 ( .A(n_360), .Y(n_404) );
NAND2x1p5_ASAP7_75t_L g468 ( .A(n_360), .B(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B1(n_368), .B2(n_373), .Y(n_362) );
INVx2_ASAP7_75t_L g382 ( .A(n_363), .Y(n_382) );
AND2x2_ASAP7_75t_L g394 ( .A(n_363), .B(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_363), .B(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g530 ( .A(n_363), .B(n_433), .Y(n_530) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
NOR2x1p5_ASAP7_75t_L g386 ( .A(n_366), .B(n_387), .Y(n_386) );
INVxp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NOR2x2_ASAP7_75t_L g407 ( .A(n_369), .B(n_408), .Y(n_407) );
OR2x6_ASAP7_75t_L g369 ( .A(n_370), .B(n_372), .Y(n_369) );
INVx2_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
OR2x2_ASAP7_75t_L g493 ( .A(n_371), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_374), .B(n_508), .Y(n_507) );
OR2x2_ASAP7_75t_L g506 ( .A(n_375), .B(n_443), .Y(n_506) );
INVx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x4_ASAP7_75t_L g446 ( .A(n_376), .B(n_443), .Y(n_446) );
NAND2x1p5_ASAP7_75t_L g470 ( .A(n_376), .B(n_387), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_380), .B1(n_383), .B2(n_388), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g402 ( .A(n_379), .Y(n_402) );
INVxp67_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g413 ( .A(n_386), .Y(n_413) );
AND2x2_ASAP7_75t_L g545 ( .A(n_386), .B(n_411), .Y(n_545) );
INVx2_ASAP7_75t_L g401 ( .A(n_387), .Y(n_401) );
INVx2_ASAP7_75t_L g453 ( .A(n_387), .Y(n_453) );
INVx1_ASAP7_75t_L g512 ( .A(n_387), .Y(n_512) );
INVx1_ASAP7_75t_L g425 ( .A(n_388), .Y(n_425) );
A2O1A1Ixp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_392), .B(n_397), .C(n_403), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVxp67_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI221xp5_ASAP7_75t_L g462 ( .A1(n_394), .A2(n_463), .B1(n_467), .B2(n_471), .C(n_474), .Y(n_462) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AND2x4_ASAP7_75t_L g398 ( .A(n_399), .B(n_402), .Y(n_398) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_399), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_399), .B(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g489 ( .A(n_405), .Y(n_489) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_413), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g465 ( .A(n_412), .B(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_415), .B(n_417), .Y(n_414) );
AOI21xp33_ASAP7_75t_L g531 ( .A1(n_415), .A2(n_532), .B(n_537), .Y(n_531) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g449 ( .A(n_418), .B(n_450), .Y(n_449) );
NOR3xp33_ASAP7_75t_L g419 ( .A(n_420), .B(n_481), .C(n_509), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_421), .B(n_462), .Y(n_420) );
AOI211xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_424), .B(n_430), .C(n_455), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OAI221xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_436), .B1(n_440), .B2(n_442), .C(n_445), .Y(n_430) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVxp67_ASAP7_75t_L g441 ( .A(n_433), .Y(n_441) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_435), .B(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_439), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g444 ( .A(n_438), .Y(n_444) );
INVx1_ASAP7_75t_L g544 ( .A(n_440), .Y(n_544) );
OR2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_447), .B1(n_449), .B2(n_451), .Y(n_445) );
INVx2_ASAP7_75t_L g519 ( .A(n_448), .Y(n_519) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_454), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g511 ( .A(n_454), .B(n_512), .Y(n_511) );
BUFx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVxp67_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g501 ( .A(n_470), .Y(n_501) );
AND2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
AOI21xp33_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_477), .B(n_479), .Y(n_474) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_482), .B(n_496), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_486), .B1(n_488), .B2(n_492), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_486), .A2(n_540), .B1(n_544), .B2(n_545), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g518 ( .A(n_495), .Y(n_518) );
AOI221xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_501), .B1(n_502), .B2(n_504), .C(n_507), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
BUFx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g529 ( .A(n_506), .Y(n_529) );
NAND3xp33_ASAP7_75t_SL g509 ( .A(n_510), .B(n_524), .C(n_539), .Y(n_509) );
O2A1O1Ixp33_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_513), .B(n_514), .C(n_515), .Y(n_510) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
OR2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_523), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_527), .B(n_530), .C(n_531), .Y(n_524) );
INVxp67_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
INVxp67_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
NOR2x1_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp33_ASAP7_75t_SL g540 ( .A(n_541), .B(n_542), .Y(n_540) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
BUFx4_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g912 ( .A(n_550), .Y(n_912) );
AND2x4_ASAP7_75t_L g550 ( .A(n_551), .B(n_763), .Y(n_550) );
AND4x1_ASAP7_75t_L g551 ( .A(n_552), .B(n_711), .C(n_731), .D(n_743), .Y(n_551) );
AOI311xp33_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_603), .A3(n_632), .B(n_648), .C(n_684), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_586), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_556), .B(n_567), .Y(n_555) );
INVx3_ASAP7_75t_L g683 ( .A(n_556), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_556), .B(n_704), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_556), .B(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g833 ( .A(n_556), .B(n_817), .Y(n_833) );
INVx3_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g722 ( .A(n_557), .B(n_652), .Y(n_722) );
INVx1_ASAP7_75t_L g785 ( .A(n_557), .Y(n_785) );
AND2x2_ASAP7_75t_L g827 ( .A(n_557), .B(n_577), .Y(n_827) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g803 ( .A(n_558), .Y(n_803) );
OAI21x1_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_561), .B(n_566), .Y(n_558) );
INVx1_ASAP7_75t_L g700 ( .A(n_561), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_566), .Y(n_701) );
AND2x2_ASAP7_75t_L g814 ( .A(n_567), .B(n_683), .Y(n_814) );
INVx1_ASAP7_75t_SL g838 ( .A(n_567), .Y(n_838) );
AND2x2_ASAP7_75t_L g851 ( .A(n_567), .B(n_802), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_567), .B(n_650), .Y(n_852) );
AND2x4_ASAP7_75t_L g567 ( .A(n_568), .B(n_577), .Y(n_567) );
AND2x2_ASAP7_75t_L g735 ( .A(n_568), .B(n_589), .Y(n_735) );
INVx3_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g652 ( .A(n_569), .Y(n_652) );
NAND2xp33_ASAP7_75t_R g696 ( .A(n_569), .B(n_589), .Y(n_696) );
AND2x2_ASAP7_75t_L g704 ( .A(n_569), .B(n_577), .Y(n_704) );
INVx1_ASAP7_75t_L g775 ( .A(n_569), .Y(n_775) );
AND2x2_ASAP7_75t_L g817 ( .A(n_569), .B(n_589), .Y(n_817) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_569), .Y(n_844) );
AND2x4_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
OR2x2_ASAP7_75t_L g698 ( .A(n_577), .B(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g784 ( .A(n_577), .B(n_785), .Y(n_784) );
AND2x2_ASAP7_75t_L g847 ( .A(n_586), .B(n_828), .Y(n_847) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g856 ( .A(n_587), .B(n_794), .Y(n_856) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g703 ( .A(n_588), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g797 ( .A(n_588), .Y(n_797) );
AND2x2_ASAP7_75t_L g802 ( .A(n_588), .B(n_803), .Y(n_802) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
BUFx2_ASAP7_75t_L g650 ( .A(n_589), .Y(n_650) );
INVx2_ASAP7_75t_L g717 ( .A(n_589), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_589), .B(n_654), .Y(n_720) );
INVx1_ASAP7_75t_L g747 ( .A(n_589), .Y(n_747) );
OR2x2_ASAP7_75t_L g754 ( .A(n_589), .B(n_652), .Y(n_754) );
AND2x2_ASAP7_75t_L g788 ( .A(n_589), .B(n_789), .Y(n_788) );
INVx3_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AOI21x1_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_593), .B(n_601), .Y(n_590) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
BUFx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_605), .B(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g771 ( .A(n_606), .B(n_708), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_623), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g879 ( .A(n_607), .B(n_660), .Y(n_879) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g758 ( .A(n_608), .B(n_625), .Y(n_758) );
AND2x2_ASAP7_75t_L g779 ( .A(n_608), .B(n_676), .Y(n_779) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
BUFx2_ASAP7_75t_R g657 ( .A(n_609), .Y(n_657) );
INVx2_ASAP7_75t_L g710 ( .A(n_609), .Y(n_710) );
AND2x2_ASAP7_75t_L g760 ( .A(n_609), .B(n_761), .Y(n_760) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_609), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_609), .B(n_635), .Y(n_808) );
AND2x2_ASAP7_75t_L g813 ( .A(n_609), .B(n_729), .Y(n_813) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AND2x4_ASAP7_75t_L g709 ( .A(n_624), .B(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g882 ( .A(n_624), .B(n_729), .Y(n_882) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g688 ( .A(n_625), .B(n_689), .Y(n_688) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_625), .Y(n_726) );
INVx1_ASAP7_75t_L g761 ( .A(n_625), .Y(n_761) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_631), .Y(n_625) );
AND2x2_ASAP7_75t_L g677 ( .A(n_626), .B(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_630), .Y(n_626) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx2_ASAP7_75t_SL g778 ( .A(n_634), .Y(n_778) );
INVx1_ASAP7_75t_L g800 ( .A(n_634), .Y(n_800) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g659 ( .A(n_635), .B(n_660), .Y(n_659) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_635), .Y(n_680) );
INVx1_ASAP7_75t_L g687 ( .A(n_635), .Y(n_687) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_635), .Y(n_708) );
AND2x4_ASAP7_75t_L g713 ( .A(n_635), .B(n_689), .Y(n_713) );
INVx2_ASAP7_75t_L g729 ( .A(n_635), .Y(n_729) );
AND2x2_ASAP7_75t_L g739 ( .A(n_635), .B(n_660), .Y(n_739) );
AO31x2_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_641), .A3(n_645), .B(n_646), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OAI22xp33_ASAP7_75t_SL g648 ( .A1(n_649), .A2(n_655), .B1(n_673), .B2(n_681), .Y(n_648) );
NAND2x1p5_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
AND2x2_ASAP7_75t_L g682 ( .A(n_651), .B(n_683), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_651), .A2(n_732), .B1(n_736), .B2(n_742), .Y(n_731) );
AND2x4_ASAP7_75t_L g828 ( .A(n_651), .B(n_829), .Y(n_828) );
NAND2x1p5_ASAP7_75t_L g873 ( .A(n_651), .B(n_796), .Y(n_873) );
AND2x4_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
AND2x4_ASAP7_75t_L g794 ( .A(n_653), .B(n_699), .Y(n_794) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g789 ( .A(n_654), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_658), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND2x4_ASAP7_75t_L g863 ( .A(n_658), .B(n_760), .Y(n_863) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OR2x2_ASAP7_75t_L g767 ( .A(n_659), .B(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_660), .B(n_710), .Y(n_730) );
AND2x2_ASAP7_75t_L g762 ( .A(n_660), .B(n_687), .Y(n_762) );
AND2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
AND2x2_ASAP7_75t_L g676 ( .A(n_662), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI21xp33_ASAP7_75t_L g886 ( .A1(n_673), .A2(n_887), .B(n_890), .Y(n_886) );
HB1xp67_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
OR2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_680), .Y(n_674) );
OR2x2_ASAP7_75t_L g849 ( .A(n_675), .B(n_687), .Y(n_849) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g870 ( .A(n_676), .Y(n_870) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g744 ( .A(n_683), .B(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_L g821 ( .A(n_683), .B(n_704), .Y(n_821) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_694), .B1(n_702), .B2(n_705), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
AND2x4_ASAP7_75t_L g806 ( .A(n_688), .B(n_807), .Y(n_806) );
AND2x2_ASAP7_75t_L g812 ( .A(n_688), .B(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g750 ( .A(n_689), .Y(n_750) );
OAI21x1_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_691), .B(n_692), .Y(n_689) );
INVxp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_697), .B(n_796), .Y(n_795) );
AND2x2_ASAP7_75t_L g891 ( .A(n_697), .B(n_892), .Y(n_891) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g755 ( .A(n_698), .Y(n_755) );
NAND2xp33_ASAP7_75t_L g831 ( .A(n_702), .B(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
BUFx3_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_707), .B(n_709), .Y(n_706) );
INVxp67_ASAP7_75t_L g823 ( .A(n_707), .Y(n_823) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g712 ( .A(n_709), .B(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g738 ( .A(n_709), .B(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g745 ( .A(n_709), .B(n_746), .Y(n_745) );
AND2x2_ASAP7_75t_L g819 ( .A(n_709), .B(n_778), .Y(n_819) );
OAI31xp33_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_714), .A3(n_716), .B(n_718), .Y(n_711) );
INVx2_ASAP7_75t_L g723 ( .A(n_712), .Y(n_723) );
INVx2_ASAP7_75t_SL g741 ( .A(n_713), .Y(n_741) );
AND2x2_ASAP7_75t_L g757 ( .A(n_713), .B(n_758), .Y(n_757) );
AND2x2_ASAP7_75t_L g854 ( .A(n_713), .B(n_768), .Y(n_854) );
AND2x4_ASAP7_75t_L g874 ( .A(n_713), .B(n_760), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_713), .B(n_725), .Y(n_889) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
BUFx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
A2O1A1Ixp33_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_721), .B(n_723), .C(n_724), .Y(n_718) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NOR2xp67_ASAP7_75t_L g774 ( .A(n_720), .B(n_775), .Y(n_774) );
OAI22xp33_ASAP7_75t_L g751 ( .A1(n_721), .A2(n_752), .B1(n_756), .B2(n_759), .Y(n_751) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g742 ( .A(n_724), .Y(n_742) );
OR2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_727), .Y(n_724) );
OR2x2_ASAP7_75t_L g740 ( .A(n_725), .B(n_741), .Y(n_740) );
AOI322xp5_ASAP7_75t_L g824 ( .A1(n_725), .A2(n_748), .A3(n_825), .B1(n_828), .B2(n_830), .C1(n_831), .C2(n_834), .Y(n_824) );
INVx2_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g885 ( .A(n_727), .Y(n_885) );
OR2x2_ASAP7_75t_L g727 ( .A(n_728), .B(n_730), .Y(n_727) );
INVx1_ASAP7_75t_L g861 ( .A(n_728), .Y(n_861) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g883 ( .A(n_730), .Y(n_883) );
INVxp67_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
BUFx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g792 ( .A(n_735), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_737), .B(n_740), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
AND2x2_ASAP7_75t_L g834 ( .A(n_739), .B(n_760), .Y(n_834) );
INVx2_ASAP7_75t_L g840 ( .A(n_740), .Y(n_840) );
AOI21xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_748), .B(n_751), .Y(n_743) );
INVx1_ASAP7_75t_L g810 ( .A(n_745), .Y(n_810) );
INVx1_ASAP7_75t_L g782 ( .A(n_746), .Y(n_782) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_747), .B(n_789), .Y(n_867) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g830 ( .A(n_749), .B(n_791), .Y(n_830) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_753), .B(n_755), .Y(n_752) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g892 ( .A(n_754), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_755), .A2(n_881), .B1(n_884), .B2(n_885), .Y(n_880) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
AND2x2_ASAP7_75t_L g860 ( .A(n_758), .B(n_861), .Y(n_860) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_759), .A2(n_777), .B1(n_780), .B2(n_786), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_760), .B(n_762), .Y(n_759) );
INVx2_ASAP7_75t_SL g791 ( .A(n_760), .Y(n_791) );
NOR2xp67_ASAP7_75t_L g763 ( .A(n_764), .B(n_845), .Y(n_763) );
NAND4xp25_ASAP7_75t_L g764 ( .A(n_765), .B(n_804), .C(n_824), .D(n_835), .Y(n_764) );
NOR3xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_776), .C(n_790), .Y(n_765) );
AOI21xp33_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_770), .B(n_772), .Y(n_766) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
BUFx2_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
NAND2x1p5_ASAP7_75t_SL g777 ( .A(n_778), .B(n_779), .Y(n_777) );
INVx1_ASAP7_75t_L g798 ( .A(n_779), .Y(n_798) );
HB1xp67_ASAP7_75t_L g857 ( .A(n_779), .Y(n_857) );
INVxp33_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
NOR2x1_ASAP7_75t_L g781 ( .A(n_782), .B(n_783), .Y(n_781) );
INVx3_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
OAI322xp33_ASAP7_75t_L g790 ( .A1(n_791), .A2(n_792), .A3(n_793), .B1(n_795), .B2(n_798), .C1(n_799), .C2(n_801), .Y(n_790) );
OR2x2_ASAP7_75t_L g822 ( .A(n_791), .B(n_823), .Y(n_822) );
INVx2_ASAP7_75t_L g805 ( .A(n_793), .Y(n_805) );
INVx2_ASAP7_75t_SL g793 ( .A(n_794), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_794), .B(n_817), .Y(n_816) );
INVx2_ASAP7_75t_L g839 ( .A(n_796), .Y(n_839) );
INVx2_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
OAI21xp33_ASAP7_75t_L g809 ( .A1(n_800), .A2(n_810), .B(n_811), .Y(n_809) );
INVx2_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx2_ASAP7_75t_L g829 ( .A(n_803), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_803), .B(n_844), .Y(n_843) );
AOI221x1_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_806), .B1(n_809), .B2(n_814), .C(n_815), .Y(n_804) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
OR2x2_ASAP7_75t_L g869 ( .A(n_808), .B(n_870), .Y(n_869) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
AOI21xp5_ASAP7_75t_L g846 ( .A1(n_812), .A2(n_847), .B(n_848), .Y(n_846) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_816), .A2(n_818), .B1(n_820), .B2(n_822), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_817), .B(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_819), .A2(n_836), .B1(n_840), .B2(n_841), .Y(n_835) );
OAI221xp5_ASAP7_75t_SL g875 ( .A1(n_820), .A2(n_869), .B1(n_876), .B2(n_877), .C(n_880), .Y(n_875) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx2_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
OR2x2_ASAP7_75t_L g837 ( .A(n_838), .B(n_839), .Y(n_837) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_838), .B(n_869), .Y(n_868) );
OR2x2_ASAP7_75t_L g842 ( .A(n_839), .B(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
HB1xp67_ASAP7_75t_L g876 ( .A(n_843), .Y(n_876) );
INVxp67_ASAP7_75t_L g866 ( .A(n_844), .Y(n_866) );
NAND3xp33_ASAP7_75t_L g845 ( .A(n_846), .B(n_855), .C(n_871), .Y(n_845) );
OAI22xp5_ASAP7_75t_L g848 ( .A1(n_849), .A2(n_850), .B1(n_852), .B2(n_853), .Y(n_848) );
INVxp67_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
AOI221xp5_ASAP7_75t_L g855 ( .A1(n_856), .A2(n_857), .B1(n_858), .B2(n_864), .C(n_868), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_859), .B(n_862), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
OR2x2_ASAP7_75t_L g865 ( .A(n_866), .B(n_867), .Y(n_865) );
INVx1_ASAP7_75t_L g884 ( .A(n_867), .Y(n_884) );
AOI211xp5_ASAP7_75t_L g871 ( .A1(n_872), .A2(n_874), .B(n_875), .C(n_886), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
HB1xp67_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
AND2x2_ASAP7_75t_L g881 ( .A(n_882), .B(n_883), .Y(n_881) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx2_ASAP7_75t_SL g890 ( .A(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
BUFx2_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
HB1xp67_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
BUFx8_ASAP7_75t_L g901 ( .A(n_896), .Y(n_901) );
INVx2_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
NOR2xp33_ASAP7_75t_L g902 ( .A(n_903), .B(n_904), .Y(n_902) );
BUFx3_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
BUFx2_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
NOR2xp33_ASAP7_75t_L g919 ( .A(n_906), .B(n_920), .Y(n_919) );
XNOR2xp5_ASAP7_75t_L g909 ( .A(n_910), .B(n_912), .Y(n_909) );
CKINVDCx20_ASAP7_75t_R g910 ( .A(n_911), .Y(n_910) );
BUFx4_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
BUFx3_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
CKINVDCx5p33_ASAP7_75t_R g917 ( .A(n_918), .Y(n_917) );
BUFx4_ASAP7_75t_R g923 ( .A(n_918), .Y(n_923) );
INVx2_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
CKINVDCx16_ASAP7_75t_R g920 ( .A(n_921), .Y(n_920) );
endmodule