module real_jpeg_2051_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_215;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_191;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

INVx2_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_1),
.A2(n_61),
.B1(n_66),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_1),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_1),
.A2(n_56),
.B1(n_58),
.B2(n_80),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_1),
.A2(n_27),
.B1(n_29),
.B2(n_80),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_1),
.A2(n_35),
.B1(n_38),
.B2(n_80),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_3),
.A2(n_35),
.B1(n_38),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_3),
.A2(n_27),
.B1(n_29),
.B2(n_48),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_4),
.A2(n_35),
.B1(n_38),
.B2(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_4),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_5),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_6),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_6),
.A2(n_55),
.B1(n_61),
.B2(n_66),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_6),
.A2(n_27),
.B1(n_29),
.B2(n_55),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_6),
.A2(n_35),
.B1(n_38),
.B2(n_55),
.Y(n_215)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_11),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_11),
.B(n_70),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_11),
.B(n_27),
.C(n_76),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_11),
.B(n_75),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_11),
.B(n_32),
.C(n_35),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_11),
.A2(n_27),
.B1(n_29),
.B2(n_112),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_11),
.B(n_46),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_11),
.B(n_41),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_11),
.A2(n_61),
.B1(n_66),
.B2(n_112),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_12),
.A2(n_35),
.B1(n_38),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_12),
.A2(n_27),
.B1(n_29),
.B2(n_50),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_13),
.A2(n_56),
.B1(n_58),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_13),
.A2(n_61),
.B1(n_66),
.B2(n_69),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_13),
.A2(n_27),
.B1(n_29),
.B2(n_69),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_13),
.A2(n_35),
.B1(n_38),
.B2(n_69),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_14),
.A2(n_27),
.B1(n_29),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_14),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_14),
.A2(n_35),
.B1(n_38),
.B2(n_40),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_14),
.A2(n_40),
.B1(n_61),
.B2(n_66),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_15),
.A2(n_26),
.B1(n_61),
.B2(n_66),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_15),
.A2(n_26),
.B1(n_35),
.B2(n_38),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_142),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_141),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_117),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_21),
.B(n_117),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_85),
.C(n_94),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_22),
.B(n_85),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_51),
.B1(n_83),
.B2(n_84),
.Y(n_22)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_42),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_24),
.B(n_42),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_39),
.B2(n_41),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_25),
.Y(n_177)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

AO22x1_ASAP7_75t_SL g75 ( 
.A1(n_27),
.A2(n_29),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_27),
.B(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_30),
.A2(n_39),
.B1(n_41),
.B2(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_30),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_30),
.A2(n_156),
.B(n_158),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_30),
.B(n_160),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_33),
.B1(n_35),
.B2(n_38),
.Y(n_34)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_34),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_34),
.A2(n_177),
.B(n_178),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_34),
.A2(n_178),
.B(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_34),
.A2(n_121),
.B1(n_157),
.B2(n_198),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_35),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_35),
.B(n_211),
.Y(n_210)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_41),
.B(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_43),
.A2(n_46),
.B(n_125),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_43),
.A2(n_112),
.B(n_192),
.Y(n_212)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_44),
.A2(n_45),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_44),
.A2(n_45),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_44),
.A2(n_45),
.B1(n_115),
.B2(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_44),
.B(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_44),
.A2(n_190),
.B(n_191),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_44),
.A2(n_45),
.B1(n_190),
.B2(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_45),
.A2(n_154),
.B(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_45),
.B(n_168),
.Y(n_192)
);

INVx3_ASAP7_75t_SL g45 ( 
.A(n_46),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_46),
.A2(n_167),
.B(n_215),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_71),
.B2(n_72),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_53),
.B(n_71),
.C(n_83),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_59),
.B1(n_68),
.B2(n_70),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_58),
.B1(n_63),
.B2(n_64),
.Y(n_67)
);

AOI32xp33_ASAP7_75t_L g109 ( 
.A1(n_56),
.A2(n_63),
.A3(n_66),
.B1(n_110),
.B2(n_113),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_56),
.B(n_112),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_56),
.A2(n_111),
.B(n_112),
.C(n_136),
.Y(n_173)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_59),
.Y(n_136)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_67),
.Y(n_59)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_60),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_60),
.B(n_101),
.Y(n_138)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_61),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_66),
.B1(n_76),
.B2(n_77),
.Y(n_82)
);

NAND2xp33_ASAP7_75t_SL g113 ( 
.A(n_61),
.B(n_64),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_61),
.B(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B(n_78),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_73),
.A2(n_74),
.B1(n_105),
.B2(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_74),
.A2(n_78),
.B(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_74),
.A2(n_104),
.B1(n_105),
.B2(n_148),
.Y(n_175)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_75),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_79),
.Y(n_106)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_90),
.B1(n_92),
.B2(n_93),
.Y(n_85)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_93),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_94),
.A2(n_95),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_102),
.C(n_107),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_96),
.A2(n_97),
.B1(n_102),
.B2(n_103),
.Y(n_245)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B(n_106),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_105),
.A2(n_106),
.B(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_107),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_114),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_108),
.A2(n_109),
.B1(n_114),
.B2(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_114),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_140),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_128),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_124),
.B1(n_126),
.B2(n_127),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_120),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_121),
.A2(n_159),
.B(n_206),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_124),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_139),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_129),
.Y(n_139)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_136),
.B(n_137),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_138),
.B(n_173),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_241),
.B(n_255),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_184),
.B(n_240),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_169),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_145),
.B(n_169),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_155),
.C(n_161),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_146),
.B(n_237),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_150),
.C(n_153),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_155),
.B(n_161),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_162),
.A2(n_163),
.B1(n_165),
.B2(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_165),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_180),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_170),
.B(n_181),
.C(n_183),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_174),
.B2(n_179),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_171),
.B(n_175),
.C(n_176),
.Y(n_248)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_174),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_235),
.B(n_239),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_225),
.B(n_234),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_207),
.B(n_224),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_201),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_201),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_193),
.B1(n_199),
.B2(n_200),
.Y(n_188)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_193),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_196),
.C(n_199),
.Y(n_226)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_202),
.A2(n_203),
.B1(n_205),
.B2(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_218),
.B(n_223),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_213),
.B(n_217),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_216),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_215),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_221),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_227),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_232),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_231),
.C(n_232),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_238),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_250),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_249),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_249),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_247),
.C(n_248),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_250),
.A2(n_256),
.B(n_257),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_254),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_254),
.Y(n_257)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);


endmodule