module fake_jpeg_29420_n_215 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_215);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_215;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx16_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_37),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_25),
.Y(n_36)
);

CKINVDCx9p33_ASAP7_75t_R g63 ( 
.A(n_36),
.Y(n_63)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_41),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_43),
.B(n_26),
.Y(n_51)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_13),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_30),
.A2(n_25),
.B1(n_17),
.B2(n_16),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_46),
.A2(n_47),
.B1(n_48),
.B2(n_60),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_20),
.B1(n_29),
.B2(n_17),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_29),
.B1(n_20),
.B2(n_14),
.Y(n_48)
);

NAND3xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_26),
.C(n_13),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_22),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_53),
.B(n_62),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_21),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_21),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_38),
.A2(n_25),
.B1(n_19),
.B2(n_22),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_61),
.B(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_15),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_38),
.B(n_15),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g99 ( 
.A(n_67),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_33),
.A2(n_28),
.B1(n_21),
.B2(n_18),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_70),
.B(n_31),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_40),
.A2(n_21),
.B1(n_18),
.B2(n_28),
.Y(n_70)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_18),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_73),
.B(n_79),
.Y(n_121)
);

AOI32xp33_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_63),
.A3(n_57),
.B1(n_59),
.B2(n_56),
.Y(n_74)
);

AOI32xp33_ASAP7_75t_L g109 ( 
.A1(n_74),
.A2(n_67),
.A3(n_49),
.B1(n_3),
.B2(n_6),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_44),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_88),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_52),
.A2(n_43),
.B1(n_42),
.B2(n_37),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_77),
.B(n_83),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_18),
.Y(n_79)
);

OR2x4_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_40),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g120 ( 
.A1(n_80),
.A2(n_49),
.B(n_2),
.Y(n_120)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_65),
.Y(n_82)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_58),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_56),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_84),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_86),
.A2(n_2),
.B(n_3),
.Y(n_126)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_0),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_94),
.Y(n_112)
);

NAND3xp33_ASAP7_75t_SL g91 ( 
.A(n_56),
.B(n_12),
.C(n_11),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_92),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_58),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_58),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_96),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_1),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_67),
.B(n_11),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx4_ASAP7_75t_SL g100 ( 
.A(n_65),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_58),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_104),
.Y(n_130)
);

XOR2x1_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_10),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_67),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_128),
.C(n_129),
.Y(n_148)
);

OR2x2_ASAP7_75t_SL g142 ( 
.A(n_120),
.B(n_89),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_71),
.B(n_1),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_122),
.B(n_123),
.Y(n_144)
);

NOR2x1_ASAP7_75t_L g123 ( 
.A(n_78),
.B(n_10),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_2),
.B(n_6),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_95),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_94),
.Y(n_129)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_136),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_84),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_134),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_130),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_84),
.B(n_86),
.Y(n_135)
);

FAx1_ASAP7_75t_SL g152 ( 
.A(n_135),
.B(n_114),
.CI(n_124),
.CON(n_152),
.SN(n_152)
);

BUFx12_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

OAI32xp33_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_103),
.A3(n_76),
.B1(n_102),
.B2(n_80),
.Y(n_137)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_97),
.B1(n_76),
.B2(n_98),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_138),
.A2(n_147),
.B1(n_116),
.B2(n_119),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_97),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_148),
.C(n_133),
.Y(n_160)
);

HAxp5_ASAP7_75t_SL g158 ( 
.A(n_140),
.B(n_141),
.CON(n_158),
.SN(n_158)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_142),
.A2(n_111),
.B1(n_131),
.B2(n_114),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_129),
.B(n_81),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_145),
.B(n_149),
.Y(n_156)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_107),
.A2(n_99),
.B1(n_82),
.B2(n_100),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_108),
.B(n_99),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_120),
.A2(n_75),
.B(n_7),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_122),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_142),
.Y(n_170)
);

XNOR2x1_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_148),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_137),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_157),
.A2(n_151),
.B1(n_141),
.B2(n_143),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_136),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_164),
.C(n_140),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g162 ( 
.A(n_144),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_136),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_121),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_166),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_156),
.B(n_123),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_175),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_170),
.B(n_171),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_173),
.A2(n_179),
.B1(n_180),
.B2(n_125),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_153),
.C(n_160),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_161),
.A2(n_164),
.B(n_167),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_155),
.Y(n_176)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_176),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_143),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_178),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_163),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_158),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_186),
.C(n_172),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_152),
.C(n_159),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_188),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_157),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_189),
.A2(n_168),
.B1(n_127),
.B2(n_117),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_170),
.C(n_172),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_179),
.Y(n_196)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_183),
.Y(n_192)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_192),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_187),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_177),
.C(n_168),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_196),
.C(n_197),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_180),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_198),
.A2(n_189),
.B1(n_191),
.B2(n_117),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_201),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_187),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_202),
.A2(n_198),
.B1(n_195),
.B2(n_158),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_203),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_200),
.C(n_201),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_206),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_193),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_207),
.A2(n_105),
.B(n_132),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_209),
.B(n_210),
.C(n_205),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_211),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_208),
.A2(n_6),
.B(n_8),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_212),
.Y(n_214)
);

BUFx24_ASAP7_75t_SL g215 ( 
.A(n_214),
.Y(n_215)
);


endmodule