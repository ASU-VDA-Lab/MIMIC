module fake_jpeg_30338_n_216 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_216);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_6),
.B(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_11),
.B(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_53),
.Y(n_63)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

CKINVDCx9p33_ASAP7_75t_R g45 ( 
.A(n_22),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_45),
.Y(n_66)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g47 ( 
.A(n_23),
.Y(n_47)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_33),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_0),
.Y(n_82)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_56),
.Y(n_68)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_55),
.B(n_32),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_0),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_35),
.B1(n_32),
.B2(n_34),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_59),
.A2(n_83),
.B1(n_3),
.B2(n_4),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_43),
.A2(n_34),
.B1(n_25),
.B2(n_30),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_61),
.A2(n_65),
.B1(n_77),
.B2(n_78),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_44),
.B(n_46),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_62),
.A2(n_40),
.B(n_37),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_38),
.A2(n_17),
.B1(n_29),
.B2(n_28),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_82),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_39),
.A2(n_17),
.B1(n_29),
.B2(n_28),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_41),
.A2(n_27),
.B1(n_18),
.B2(n_20),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_48),
.B(n_26),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_79),
.B(n_57),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_54),
.A2(n_27),
.B1(n_18),
.B2(n_20),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_80),
.A2(n_85),
.B1(n_2),
.B2(n_3),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_47),
.A2(n_30),
.B1(n_1),
.B2(n_2),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_84),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_50),
.B1(n_53),
.B2(n_51),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_50),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_97),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_24),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_92),
.Y(n_116)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_91),
.A2(n_110),
.B1(n_86),
.B2(n_81),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_57),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_95),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_69),
.B(n_57),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_94),
.B(n_58),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_14),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_52),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_114),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_1),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_66),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_104),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_70),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_107),
.Y(n_124)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_103),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_67),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_62),
.B(n_49),
.C(n_45),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_58),
.C(n_7),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_10),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_113),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_111),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_4),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_13),
.Y(n_123)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_75),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_90),
.A2(n_101),
.B1(n_97),
.B2(n_108),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_118),
.A2(n_128),
.B1(n_130),
.B2(n_133),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_123),
.B(n_112),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_86),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_100),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_74),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_135),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_90),
.A2(n_81),
.B1(n_60),
.B2(n_76),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_107),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_91),
.A2(n_76),
.B1(n_70),
.B2(n_74),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_104),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_110),
.C(n_114),
.Y(n_149)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_141),
.Y(n_170)
);

AOI322xp5_ASAP7_75t_SL g142 ( 
.A1(n_121),
.A2(n_99),
.A3(n_123),
.B1(n_116),
.B2(n_98),
.C1(n_118),
.C2(n_126),
.Y(n_142)
);

BUFx24_ASAP7_75t_SL g168 ( 
.A(n_142),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_145),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_146),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_94),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_98),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_89),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_148),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_103),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_155),
.Y(n_161)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_156),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_133),
.A2(n_128),
.B(n_132),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_152),
.A2(n_153),
.B(n_132),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_132),
.A2(n_96),
.B(n_102),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_119),
.A2(n_125),
.B1(n_130),
.B2(n_137),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_154),
.A2(n_134),
.B1(n_106),
.B2(n_117),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_96),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

OAI32xp33_ASAP7_75t_L g158 ( 
.A1(n_146),
.A2(n_137),
.A3(n_124),
.B1(n_136),
.B2(n_105),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_154),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_134),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_160),
.B(n_164),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_151),
.A2(n_106),
.B1(n_113),
.B2(n_127),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_169),
.A2(n_172),
.B(n_148),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_138),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_171),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_151),
.A2(n_127),
.B1(n_113),
.B2(n_9),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_173),
.A2(n_176),
.B1(n_175),
.B2(n_181),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_147),
.C(n_144),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_179),
.C(n_181),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_159),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_177),
.B(n_182),
.Y(n_185)
);

XNOR2x1_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_149),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_180),
.A2(n_169),
.B1(n_158),
.B2(n_166),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_155),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_156),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_157),
.A2(n_152),
.B(n_153),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_183),
.A2(n_164),
.B(n_172),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_143),
.C(n_140),
.Y(n_184)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_184),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_174),
.Y(n_195)
);

AO21x1_ASAP7_75t_L g198 ( 
.A1(n_187),
.A2(n_167),
.B(n_139),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_180),
.A2(n_170),
.B1(n_165),
.B2(n_162),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_189),
.A2(n_193),
.B1(n_184),
.B2(n_170),
.Y(n_199)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_182),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_192),
.Y(n_200)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_187),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_199),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_197),
.C(n_190),
.Y(n_201)
);

NOR2x1_ASAP7_75t_SL g196 ( 
.A(n_193),
.B(n_168),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_196),
.A2(n_198),
.B(n_185),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_179),
.C(n_175),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_205),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_204),
.Y(n_206)
);

O2A1O1Ixp5_ASAP7_75t_L g204 ( 
.A1(n_198),
.A2(n_189),
.B(n_186),
.C(n_188),
.Y(n_204)
);

MAJx2_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_200),
.C(n_195),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_202),
.A2(n_141),
.B(n_150),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_208),
.B(n_209),
.Y(n_210)
);

NAND4xp25_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_5),
.C(n_8),
.D(n_9),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_8),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_212),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_207),
.A2(n_8),
.B1(n_9),
.B2(n_202),
.Y(n_212)
);

FAx1_ASAP7_75t_SL g213 ( 
.A(n_212),
.B(n_207),
.CI(n_210),
.CON(n_213),
.SN(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_213),
.B(n_214),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_213),
.Y(n_216)
);


endmodule