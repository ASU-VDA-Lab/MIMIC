module fake_jpeg_2034_n_150 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_150);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_19),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_39),
.B(n_0),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_59),
.A2(n_51),
.B(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_61),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_56),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_61),
.A2(n_38),
.B1(n_44),
.B2(n_46),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_72),
.B1(n_49),
.B2(n_57),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_38),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_60),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_47),
.B1(n_41),
.B2(n_46),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_47),
.B1(n_42),
.B2(n_49),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_52),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_75),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_54),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_77),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_58),
.B(n_60),
.C(n_59),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_63),
.A2(n_62),
.B1(n_67),
.B2(n_71),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_84),
.B1(n_81),
.B2(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_87),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_86),
.Y(n_99)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

O2A1O1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_56),
.B(n_43),
.C(n_62),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_1),
.B(n_2),
.Y(n_102)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_43),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_64),
.B1(n_63),
.B2(n_50),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_89),
.A2(n_100),
.B1(n_4),
.B2(n_5),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_75),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_92),
.B(n_3),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_64),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_94),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_0),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_37),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_6),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_98),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_86),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_87),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_97),
.C(n_102),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_102),
.Y(n_105)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_104),
.Y(n_126)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_109),
.Y(n_127)
);

OAI21x1_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_12),
.B(n_13),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_4),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_108),
.B(n_117),
.Y(n_129)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_116),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_15),
.B1(n_32),
.B2(n_33),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_95),
.A2(n_21),
.B1(n_35),
.B2(n_34),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_114),
.A2(n_36),
.B(n_112),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_115),
.A2(n_89),
.B1(n_98),
.B2(n_14),
.Y(n_121)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_99),
.B(n_7),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_9),
.B(n_10),
.Y(n_118)
);

OA21x2_ASAP7_75t_L g124 ( 
.A1(n_118),
.A2(n_12),
.B(n_13),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_24),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_10),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_14),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_121),
.A2(n_105),
.B1(n_118),
.B2(n_106),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_113),
.B(n_27),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_130),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_125),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_124),
.A2(n_132),
.B(n_114),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_17),
.C(n_28),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_131),
.A2(n_115),
.B1(n_110),
.B2(n_104),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_133),
.A2(n_136),
.B(n_138),
.Y(n_140)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_127),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_135),
.A2(n_128),
.B(n_121),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_124),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_142),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_139),
.A2(n_138),
.B1(n_126),
.B2(n_135),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_144),
.B(n_129),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_143),
.Y(n_146)
);

NAND2x1_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_143),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_140),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_SL g149 ( 
.A1(n_148),
.A2(n_124),
.B(n_122),
.C(n_137),
.Y(n_149)
);

BUFx24_ASAP7_75t_SL g150 ( 
.A(n_149),
.Y(n_150)
);


endmodule