module fake_jpeg_442_n_189 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_189);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_189;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx11_ASAP7_75t_SL g62 ( 
.A(n_34),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_20),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_70),
.Y(n_74)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_54),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_65),
.Y(n_78)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_75),
.B(n_53),
.Y(n_91)
);

AO22x1_ASAP7_75t_SL g76 ( 
.A1(n_71),
.A2(n_60),
.B1(n_56),
.B2(n_63),
.Y(n_76)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_57),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_77),
.B(n_82),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_64),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_67),
.A2(n_56),
.B1(n_51),
.B2(n_59),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_79),
.A2(n_81),
.B1(n_83),
.B2(n_53),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_66),
.A2(n_51),
.B1(n_59),
.B2(n_52),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_50),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_69),
.A2(n_58),
.B1(n_63),
.B2(n_61),
.Y(n_83)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_80),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_87),
.B(n_89),
.Y(n_107)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_50),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_95),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_96),
.Y(n_108)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_44),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_61),
.B1(n_53),
.B2(n_55),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_74),
.B1(n_77),
.B2(n_75),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_94),
.A2(n_101),
.B1(n_49),
.B2(n_1),
.Y(n_110)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_74),
.Y(n_99)
);

INVx5_ASAP7_75t_SL g120 ( 
.A(n_99),
.Y(n_120)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_100),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_76),
.A2(n_53),
.B1(n_49),
.B2(n_2),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_103),
.A2(n_110),
.B1(n_26),
.B2(n_25),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_97),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_114),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_46),
.C(n_45),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_11),
.C(n_12),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_SL g112 ( 
.A1(n_85),
.A2(n_30),
.B(n_43),
.C(n_41),
.Y(n_112)
);

A2O1A1O1Ixp25_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_4),
.B(n_5),
.C(n_6),
.D(n_7),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_0),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_1),
.B(n_2),
.Y(n_115)
);

O2A1O1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_115),
.A2(n_111),
.B(n_112),
.C(n_121),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_3),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_118),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_96),
.B(n_3),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_117),
.B(n_33),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_88),
.Y(n_118)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_121),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_101),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_105),
.C(n_18),
.Y(n_156)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_126),
.B(n_134),
.Y(n_150)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_129),
.A2(n_108),
.B(n_103),
.Y(n_143)
);

BUFx24_ASAP7_75t_SL g130 ( 
.A(n_104),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_130),
.B(n_132),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_102),
.A2(n_100),
.B1(n_94),
.B2(n_6),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_135),
.B1(n_138),
.B2(n_106),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_4),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_110),
.A2(n_39),
.B1(n_36),
.B2(n_35),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_133),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_5),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_120),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_137),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_10),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_28),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_140),
.C(n_11),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_152),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_145),
.B(n_146),
.Y(n_168)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_21),
.C(n_19),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_156),
.C(n_140),
.Y(n_161)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_105),
.B1(n_13),
.B2(n_14),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_153),
.A2(n_12),
.B1(n_13),
.B2(n_16),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_124),
.Y(n_155)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_126),
.B(n_17),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_156),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_151),
.C(n_160),
.Y(n_174)
);

OAI321xp33_ASAP7_75t_L g163 ( 
.A1(n_150),
.A2(n_129),
.A3(n_133),
.B1(n_15),
.B2(n_16),
.C(n_17),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_163),
.A2(n_144),
.B1(n_149),
.B2(n_154),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_166),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_158),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_172),
.C(n_173),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_171),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_159),
.B(n_144),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_142),
.Y(n_173)
);

FAx1_ASAP7_75t_SL g176 ( 
.A(n_174),
.B(n_162),
.CI(n_164),
.CON(n_176),
.SN(n_176)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_172),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_175),
.A2(n_167),
.B1(n_164),
.B2(n_162),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_178),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_177),
.C(n_170),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_177),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_176),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_184),
.B(n_179),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_179),
.B(n_175),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_176),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_187),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_180),
.C(n_178),
.Y(n_189)
);


endmodule