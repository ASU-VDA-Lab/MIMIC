module fake_jpeg_14634_n_101 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_101);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_101;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_24),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_47),
.Y(n_53)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_51),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_50),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_46),
.B(n_38),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_59),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_48),
.B(n_45),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_60),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_44),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_33),
.Y(n_61)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_55),
.B(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_68),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_0),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_74),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_56),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_1),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_59),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_5),
.B(n_7),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_3),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_13),
.C(n_15),
.Y(n_82)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_76),
.A2(n_77),
.B(n_72),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_8),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_16),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_84),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_66),
.Y(n_85)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

BUFx4f_ASAP7_75t_SL g86 ( 
.A(n_79),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_87),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_63),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_75),
.Y(n_92)
);

OA21x2_ASAP7_75t_SL g94 ( 
.A1(n_92),
.A2(n_93),
.B(n_89),
.Y(n_94)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_80),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

AOI21x1_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_88),
.B(n_22),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_21),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_23),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_25),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_26),
.Y(n_101)
);


endmodule