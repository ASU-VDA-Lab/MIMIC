module fake_jpeg_21531_n_262 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_262);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_262;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx4_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_3),
.B(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_1),
.B(n_11),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_27),
.B(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_35),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx5_ASAP7_75t_SL g67 ( 
.A(n_37),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_33),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_43),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_17),
.B1(n_28),
.B2(n_27),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_46),
.A2(n_56),
.B1(n_62),
.B2(n_70),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_22),
.B(n_17),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_64),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_49),
.B(n_51),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_57),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_17),
.B1(n_28),
.B2(n_25),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_54),
.A2(n_32),
.B1(n_42),
.B2(n_34),
.Y(n_89)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_68),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_43),
.A2(n_28),
.B1(n_25),
.B2(n_19),
.Y(n_56)
);

NOR2x1_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_20),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_66),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_44),
.A2(n_25),
.B1(n_19),
.B2(n_23),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_19),
.B1(n_23),
.B2(n_29),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_63),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_30),
.C(n_26),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_39),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_71),
.B(n_73),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_66),
.B(n_40),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_76),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_42),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_24),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_84),
.Y(n_109)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_49),
.B(n_39),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_87),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_24),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_86),
.Y(n_130)
);

OAI32xp33_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_30),
.A3(n_32),
.B1(n_39),
.B2(n_42),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_88),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_89),
.A2(n_104),
.B1(n_16),
.B2(n_13),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_56),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_91),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_62),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_33),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_94),
.C(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_103),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_61),
.A2(n_32),
.B(n_33),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_60),
.A2(n_34),
.B1(n_24),
.B2(n_3),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_95),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_34),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_98),
.Y(n_129)
);

AOI32xp33_ASAP7_75t_L g98 ( 
.A1(n_60),
.A2(n_9),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_0),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_105),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_10),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_52),
.B(n_0),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_106),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_60),
.B1(n_52),
.B2(n_67),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_110),
.A2(n_113),
.B1(n_115),
.B2(n_127),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_52),
.B1(n_67),
.B2(n_50),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_86),
.A2(n_67),
.B1(n_50),
.B2(n_7),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_76),
.A2(n_5),
.B(n_6),
.Y(n_117)
);

MAJx2_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_94),
.C(n_83),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_85),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_123),
.A2(n_126),
.B1(n_98),
.B2(n_99),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_72),
.B(n_16),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_132),
.C(n_134),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_82),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_74),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_131),
.B(n_80),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_82),
.B(n_12),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_73),
.B(n_75),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_101),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_79),
.B(n_15),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_140),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_137),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_133),
.B(n_101),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_138),
.B(n_141),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_83),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_121),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_120),
.B(n_80),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_142),
.B(n_154),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_143),
.A2(n_129),
.B1(n_124),
.B2(n_134),
.Y(n_164)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_145),
.A2(n_161),
.B1(n_132),
.B2(n_130),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_122),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_152),
.Y(n_171)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_151),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_83),
.C(n_92),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_125),
.C(n_134),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_78),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_155),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_124),
.A2(n_85),
.B1(n_92),
.B2(n_87),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_157),
.A2(n_108),
.B1(n_116),
.B2(n_128),
.Y(n_166)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_114),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_160),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_159),
.Y(n_163)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_164),
.A2(n_112),
.B1(n_104),
.B2(n_81),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_167),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_157),
.A2(n_123),
.B1(n_131),
.B2(n_130),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_184),
.C(n_139),
.Y(n_186)
);

AOI21x1_ASAP7_75t_L g172 ( 
.A1(n_140),
.A2(n_105),
.B(n_127),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_172),
.A2(n_178),
.B(n_158),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_175),
.A2(n_180),
.B(n_149),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_135),
.A2(n_132),
.B(n_111),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_147),
.A2(n_107),
.B1(n_111),
.B2(n_88),
.Y(n_180)
);

AOI221xp5_ASAP7_75t_L g183 ( 
.A1(n_143),
.A2(n_136),
.B1(n_135),
.B2(n_145),
.C(n_148),
.Y(n_183)
);

A2O1A1O1Ixp25_ASAP7_75t_L g198 ( 
.A1(n_183),
.A2(n_107),
.B(n_150),
.C(n_97),
.D(n_71),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_93),
.C(n_97),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_194),
.C(n_200),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_187),
.A2(n_190),
.B(n_193),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_181),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_188),
.B(n_202),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_171),
.A2(n_144),
.B(n_155),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_160),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_196),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_170),
.B(n_139),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_197),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_156),
.Y(n_194)
);

XNOR2x1_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_156),
.Y(n_195)
);

OAI322xp33_ASAP7_75t_L g211 ( 
.A1(n_195),
.A2(n_198),
.A3(n_172),
.B1(n_175),
.B2(n_185),
.C1(n_167),
.C2(n_176),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_180),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_159),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_103),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_201),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_102),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_174),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_102),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_203),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_81),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_204),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_164),
.C(n_178),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_214),
.C(n_189),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_196),
.A2(n_185),
.B1(n_182),
.B2(n_173),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_210),
.A2(n_182),
.B1(n_201),
.B2(n_179),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_211),
.A2(n_198),
.B1(n_168),
.B2(n_165),
.Y(n_231)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_204),
.Y(n_212)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_179),
.C(n_176),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_216),
.Y(n_229)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_218),
.Y(n_227)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_202),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_165),
.Y(n_232)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_221),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_195),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_223),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_193),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_188),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_224),
.B(n_230),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_187),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_226),
.C(n_214),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_189),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_231),
.B(n_217),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_219),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_218),
.A2(n_163),
.B1(n_104),
.B2(n_168),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_233),
.A2(n_210),
.B1(n_163),
.B2(n_212),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_222),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_237),
.A2(n_240),
.B1(n_213),
.B2(n_221),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_241),
.Y(n_245)
);

OAI31xp33_ASAP7_75t_L g241 ( 
.A1(n_227),
.A2(n_215),
.A3(n_216),
.B(n_220),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_206),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_242),
.B(n_232),
.Y(n_246)
);

OAI221xp5_ASAP7_75t_L g243 ( 
.A1(n_234),
.A2(n_220),
.B1(n_217),
.B2(n_215),
.C(n_229),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_243),
.A2(n_248),
.B(n_241),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_236),
.B(n_226),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_244),
.B(n_246),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_235),
.C(n_225),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_249),
.B(n_250),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_245),
.A2(n_240),
.B1(n_239),
.B2(n_228),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_253),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_247),
.A2(n_207),
.B(n_239),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_251),
.B(n_223),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_251),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_257),
.A2(n_258),
.B(n_207),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_194),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_257),
.B(n_256),
.C(n_235),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_259),
.B(n_260),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_261),
.B(n_13),
.Y(n_262)
);


endmodule