module fake_jpeg_21932_n_219 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_219);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_219;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_41),
.Y(n_52)
);

BUFx4f_ASAP7_75t_SL g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_0),
.Y(n_63)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_38),
.B1(n_40),
.B2(n_31),
.Y(n_44)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_31),
.B1(n_25),
.B2(n_20),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_43),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_44),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_22),
.B1(n_23),
.B2(n_31),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_23),
.B1(n_25),
.B2(n_22),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_15),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_1),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_34),
.B(n_15),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_21),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_20),
.B1(n_19),
.B2(n_15),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_56),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_21),
.B1(n_30),
.B2(n_27),
.Y(n_54)
);

AO22x1_ASAP7_75t_SL g79 ( 
.A1(n_54),
.A2(n_62),
.B1(n_46),
.B2(n_17),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_29),
.B1(n_18),
.B2(n_30),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_55),
.A2(n_28),
.B(n_2),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_20),
.C(n_29),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVxp33_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_16),
.Y(n_60)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_27),
.B1(n_18),
.B2(n_16),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_1),
.Y(n_75)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_65),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_49),
.B(n_21),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_52),
.B(n_51),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_74),
.C(n_71),
.Y(n_101)
);

AO22x2_ASAP7_75t_SL g68 ( 
.A1(n_54),
.A2(n_28),
.B1(n_17),
.B2(n_21),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_68),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_54),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_75),
.Y(n_94)
);

NAND2x1_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_52),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_53),
.A2(n_21),
.B(n_28),
.C(n_17),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_78),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_55),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_79),
.A2(n_83),
.B1(n_63),
.B2(n_54),
.Y(n_84)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_60),
.B(n_21),
.Y(n_82)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_84),
.A2(n_99),
.B1(n_104),
.B2(n_67),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_86),
.B(n_1),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_90),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_66),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_93),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_78),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_96),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_62),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_45),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_98),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_105),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_45),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_64),
.A2(n_61),
.B1(n_59),
.B2(n_57),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_68),
.Y(n_118)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_79),
.Y(n_108)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_103),
.A2(n_79),
.B1(n_68),
.B2(n_73),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_115),
.B1(n_124),
.B2(n_105),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_108),
.A2(n_125),
.B(n_92),
.Y(n_135)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_110),
.Y(n_131)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_105),
.B1(n_50),
.B2(n_80),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_87),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_114),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_90),
.A2(n_68),
.B1(n_71),
.B2(n_58),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_123),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_120),
.Y(n_129)
);

OAI32xp33_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_89),
.A3(n_102),
.B1(n_98),
.B2(n_95),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_69),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_126),
.Y(n_134)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_102),
.A2(n_28),
.B1(n_69),
.B2(n_50),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_85),
.B(n_2),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_119),
.A2(n_101),
.B(n_86),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_127),
.A2(n_132),
.B(n_135),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_113),
.A2(n_84),
.B1(n_101),
.B2(n_104),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_138),
.B1(n_110),
.B2(n_6),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_111),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_142),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_123),
.A2(n_92),
.B(n_94),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_122),
.B(n_94),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_124),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_139),
.B1(n_109),
.B2(n_106),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_108),
.A2(n_121),
.B(n_119),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_116),
.A2(n_2),
.B(n_3),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_125),
.Y(n_147)
);

NOR4xp25_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_112),
.C(n_120),
.D(n_115),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_141),
.B(n_4),
.Y(n_163)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_126),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_144),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_107),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_145),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_3),
.Y(n_146)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_161),
.Y(n_165)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_150),
.A2(n_154),
.B(n_162),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_118),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_163),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_137),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_153),
.Y(n_175)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_158),
.A2(n_136),
.B1(n_134),
.B2(n_144),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_4),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_4),
.Y(n_162)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_129),
.C(n_127),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_168),
.C(n_176),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_128),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_177),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_139),
.C(n_141),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_169),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_133),
.C(n_142),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_135),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_158),
.B1(n_131),
.B2(n_152),
.Y(n_179)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_165),
.B(n_132),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_181),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_149),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_172),
.A2(n_131),
.B1(n_154),
.B2(n_150),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_182),
.A2(n_130),
.B1(n_177),
.B2(n_138),
.Y(n_193)
);

AOI31xp67_ASAP7_75t_L g184 ( 
.A1(n_169),
.A2(n_140),
.A3(n_147),
.B(n_162),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_170),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_173),
.A2(n_159),
.B(n_146),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_186),
.A2(n_188),
.B(n_176),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_164),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_166),
.C(n_168),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_189),
.B(n_191),
.Y(n_201)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_170),
.C(n_174),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_186),
.Y(n_192)
);

NAND4xp25_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_195),
.C(n_187),
.D(n_182),
.Y(n_198)
);

NAND2x1_ASAP7_75t_SL g204 ( 
.A(n_193),
.B(n_189),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_167),
.Y(n_195)
);

NOR2xp67_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_6),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_198),
.A2(n_203),
.B1(n_204),
.B2(n_193),
.Y(n_205)
);

NAND4xp25_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_178),
.C(n_185),
.D(n_9),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_199),
.B(n_9),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_194),
.A2(n_6),
.B(n_7),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_7),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_208),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_191),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_206),
.B(n_207),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_195),
.C(n_11),
.Y(n_209)
);

NAND2x1p5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_10),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_209),
.A2(n_200),
.B1(n_204),
.B2(n_12),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_211),
.B(n_213),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_210),
.A2(n_212),
.B(n_207),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_215),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_10),
.C(n_11),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_216),
.B(n_12),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_217),
.Y(n_219)
);


endmodule