module real_jpeg_32956_n_17 (n_8, n_0, n_2, n_132, n_125, n_10, n_9, n_129, n_12, n_124, n_130, n_134, n_6, n_128, n_133, n_11, n_14, n_131, n_7, n_3, n_127, n_5, n_4, n_1, n_126, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_132;
input n_125;
input n_10;
input n_9;
input n_129;
input n_12;
input n_124;
input n_130;
input n_134;
input n_6;
input n_128;
input n_133;
input n_11;
input n_14;
input n_131;
input n_7;
input n_3;
input n_127;
input n_5;
input n_4;
input n_1;
input n_126;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_0),
.B(n_27),
.Y(n_115)
);

FAx1_ASAP7_75t_SL g17 ( 
.A(n_1),
.B(n_18),
.CI(n_23),
.CON(n_17),
.SN(n_17)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_2),
.B(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_3),
.B(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_3),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_4),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_5),
.B(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

AOI221xp5_ASAP7_75t_L g43 ( 
.A1(n_8),
.A2(n_12),
.B1(n_44),
.B2(n_49),
.C(n_52),
.Y(n_43)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_9),
.Y(n_86)
);

AOI322xp5_ASAP7_75t_L g109 ( 
.A1(n_9),
.A2(n_78),
.A3(n_80),
.B1(n_88),
.B2(n_110),
.C1(n_112),
.C2(n_134),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_10),
.Y(n_85)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_11),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_11),
.B(n_90),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_12),
.B(n_44),
.C(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_13),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_13),
.B(n_94),
.Y(n_107)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_14),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_14),
.B(n_101),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_15),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_15),
.B(n_118),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

OAI21x1_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_116),
.B(n_121),
.Y(n_23)
);

AOI21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_32),
.B(n_115),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVxp67_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

AOI31xp67_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_71),
.A3(n_99),
.B(n_105),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_66),
.C(n_67),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_56),
.B(n_65),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_43),
.B1(n_54),
.B2(n_55),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_45),
.B(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_126),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_64),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_64),
.Y(n_65)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_70),
.B(n_119),
.Y(n_118)
);

NOR3xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_87),
.C(n_93),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_72),
.A2(n_106),
.B(n_109),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_78),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NOR3xp33_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_93),
.C(n_111),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_86),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_130),
.Y(n_80)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OA21x2_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_107),
.B(n_108),
.Y(n_106)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2x1_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_104),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_124),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_125),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_127),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_128),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_129),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_131),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_132),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_133),
.Y(n_102)
);


endmodule