module fake_jpeg_1938_n_218 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_218);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_218;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_34),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_9),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_1),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_27),
.Y(n_77)
);

BUFx2_ASAP7_75t_R g78 ( 
.A(n_61),
.Y(n_78)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g96 ( 
.A(n_79),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_0),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_77),
.Y(n_94)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_58),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_83),
.B(n_78),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_82),
.A2(n_64),
.B1(n_58),
.B2(n_59),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_86),
.A2(n_95),
.B1(n_98),
.B2(n_72),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_89),
.B(n_92),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_83),
.A2(n_75),
.B1(n_68),
.B2(n_72),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_56),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_79),
.A2(n_85),
.B1(n_68),
.B2(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_57),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_84),
.A2(n_64),
.B1(n_76),
.B2(n_67),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_65),
.B1(n_76),
.B2(n_67),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_104),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_91),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_102),
.B(n_91),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_70),
.C(n_62),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_11),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_91),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_73),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_107),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_74),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_3),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_63),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_114),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_99),
.Y(n_110)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_71),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_54),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_118),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_61),
.B(n_53),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_10),
.Y(n_137)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_65),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_116),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_122),
.B1(n_124),
.B2(n_126),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_53),
.B1(n_84),
.B2(n_68),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_56),
.B1(n_60),
.B2(n_69),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_105),
.A2(n_56),
.B1(n_1),
.B2(n_2),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_128),
.B(n_13),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_108),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_132),
.B1(n_133),
.B2(n_136),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_106),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_118),
.A2(n_5),
.B1(n_7),
.B2(n_10),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_113),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_12),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_140),
.B(n_14),
.Y(n_152)
);

NAND3xp33_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_125),
.C(n_134),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_144),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_111),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_145),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_137),
.A2(n_110),
.B(n_117),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_132),
.B(n_112),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_21),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_12),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_154),
.Y(n_184)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_148),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_127),
.A2(n_13),
.B(n_14),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_161),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_150),
.B(n_152),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_15),
.B(n_17),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_153),
.A2(n_29),
.B(n_30),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_15),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_38),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_162),
.C(n_164),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_131),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_158),
.B(n_160),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_119),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_159),
.A2(n_162),
.B1(n_155),
.B2(n_151),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_136),
.B(n_18),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_19),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_40),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_20),
.Y(n_163)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_163),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_42),
.Y(n_164)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_148),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_168),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_141),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_156),
.A2(n_43),
.B(n_22),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_170),
.A2(n_173),
.B(n_159),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_183),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_156),
.A2(n_21),
.B(n_26),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_155),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_181),
.B(n_182),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_165),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_151),
.A2(n_32),
.B1(n_35),
.B2(n_37),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_164),
.C(n_157),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_167),
.C(n_174),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_167),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_192),
.Y(n_197)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_176),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_195),
.Y(n_196)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_179),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_192),
.A2(n_171),
.B1(n_183),
.B2(n_169),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_198),
.A2(n_199),
.B1(n_201),
.B2(n_187),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_189),
.A2(n_175),
.B1(n_178),
.B2(n_184),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_203),
.C(n_44),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_191),
.A2(n_177),
.B1(n_170),
.B2(n_181),
.Y(n_201)
);

OAI21x1_ASAP7_75t_SL g209 ( 
.A1(n_204),
.A2(n_206),
.B(n_203),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_197),
.A2(n_188),
.B(n_173),
.Y(n_205)
);

AO21x1_ASAP7_75t_L g211 ( 
.A1(n_205),
.A2(n_207),
.B(n_200),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_L g206 ( 
.A1(n_197),
.A2(n_189),
.B1(n_202),
.B2(n_190),
.Y(n_206)
);

AO21x1_ASAP7_75t_L g207 ( 
.A1(n_196),
.A2(n_172),
.B(n_186),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_208),
.A2(n_45),
.B(n_46),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_209),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_210),
.B(n_211),
.Y(n_213)
);

FAx1_ASAP7_75t_SL g214 ( 
.A(n_212),
.B(n_206),
.CI(n_207),
.CON(n_214),
.SN(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_213),
.C(n_49),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_47),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_50),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_51),
.Y(n_218)
);


endmodule