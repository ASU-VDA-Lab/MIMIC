module fake_jpeg_19659_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVxp33_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_39),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx4f_ASAP7_75t_SL g90 ( 
.A(n_46),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_63),
.Y(n_101)
);

BUFx16f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_69),
.Y(n_103)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_38),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_67),
.B(n_88),
.Y(n_123)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_43),
.B1(n_39),
.B2(n_35),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_73),
.A2(n_26),
.B1(n_17),
.B2(n_20),
.Y(n_107)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_74),
.A2(n_68),
.B1(n_66),
.B2(n_71),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_45),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_75),
.B(n_80),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_41),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_79),
.C(n_31),
.Y(n_102)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_82),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_39),
.C(n_37),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_40),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_61),
.A2(n_43),
.B1(n_36),
.B2(n_35),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_81),
.A2(n_17),
.B1(n_20),
.B2(n_26),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_40),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_43),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_92),
.Y(n_96)
);

CKINVDCx12_ASAP7_75t_R g84 ( 
.A(n_46),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_85),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_52),
.B(n_24),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_24),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_87),
.Y(n_116)
);

CKINVDCx12_ASAP7_75t_R g87 ( 
.A(n_47),
.Y(n_87)
);

NAND2xp33_ASAP7_75t_SL g88 ( 
.A(n_52),
.B(n_42),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_25),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_91),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_36),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_19),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_94),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_37),
.B1(n_42),
.B2(n_25),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_100),
.A2(n_109),
.B1(n_115),
.B2(n_122),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_120),
.Y(n_131)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_117),
.Y(n_125)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_74),
.A2(n_16),
.B1(n_30),
.B2(n_21),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_79),
.A2(n_19),
.B1(n_30),
.B2(n_21),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_67),
.B(n_31),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_31),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_121),
.Y(n_139)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_18),
.C(n_22),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_31),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_88),
.A2(n_32),
.B1(n_28),
.B2(n_29),
.Y(n_122)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_68),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_95),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_126),
.B(n_141),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_123),
.A2(n_117),
.B(n_102),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_128),
.A2(n_136),
.B(n_120),
.Y(n_160)
);

INVx4_ASAP7_75t_SL g129 ( 
.A(n_99),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_135),
.Y(n_162)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_R g136 ( 
.A(n_123),
.B(n_97),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_97),
.A2(n_34),
.B1(n_69),
.B2(n_81),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_101),
.B1(n_100),
.B2(n_107),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_96),
.A2(n_77),
.B1(n_76),
.B2(n_70),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_138),
.A2(n_124),
.B1(n_108),
.B2(n_106),
.Y(n_169)
);

AND2x6_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_90),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_105),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_142),
.B(n_143),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_104),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_90),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_146),
.Y(n_172)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_90),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

XNOR2x1_ASAP7_75t_SL g152 ( 
.A(n_115),
.B(n_118),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_152),
.A2(n_139),
.B(n_125),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_98),
.B(n_111),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_23),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_130),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_155),
.B(n_170),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_129),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_141),
.A2(n_121),
.B(n_98),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_158),
.A2(n_164),
.B(n_165),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_160),
.A2(n_166),
.B(n_168),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_101),
.B(n_122),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_133),
.A2(n_109),
.B(n_119),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_104),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_169),
.A2(n_173),
.B1(n_181),
.B2(n_140),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_147),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_112),
.B1(n_76),
.B2(n_66),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_128),
.A2(n_18),
.B1(n_22),
.B2(n_32),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_127),
.A2(n_136),
.B(n_125),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_176),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_144),
.A2(n_32),
.B1(n_28),
.B2(n_22),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_147),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_177),
.B(n_179),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_64),
.C(n_22),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_186),
.C(n_132),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_135),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_180),
.B(n_167),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_138),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_127),
.A2(n_23),
.B(n_1),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_183),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_28),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_126),
.Y(n_185)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_185),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_131),
.B(n_64),
.C(n_72),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_187),
.A2(n_218),
.B1(n_181),
.B2(n_165),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_184),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_188),
.B(n_198),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_186),
.Y(n_190)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_143),
.Y(n_192)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_163),
.B(n_10),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_194),
.B(n_199),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_195),
.A2(n_210),
.B1(n_170),
.B2(n_177),
.Y(n_226)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_196),
.Y(n_240)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_154),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_140),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_154),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_203),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_209),
.Y(n_225)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

XNOR2x2_ASAP7_75t_SL g204 ( 
.A(n_160),
.B(n_150),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_206),
.Y(n_231)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_157),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_171),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_208),
.Y(n_241)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_157),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_161),
.B(n_23),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_161),
.A2(n_132),
.B1(n_150),
.B2(n_72),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_178),
.Y(n_219)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_213),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_167),
.B(n_7),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_216),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_163),
.B(n_7),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_7),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_217),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_0),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_191),
.C(n_196),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_221),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_212),
.B(n_175),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_222),
.B(n_223),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_197),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_226),
.A2(n_232),
.B1(n_213),
.B2(n_201),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_188),
.A2(n_197),
.B1(n_201),
.B2(n_173),
.Y(n_229)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_195),
.A2(n_159),
.B1(n_166),
.B2(n_155),
.Y(n_232)
);

NOR4xp25_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_168),
.C(n_158),
.D(n_166),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_233),
.B(n_218),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_164),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_243),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_204),
.A2(n_182),
.B(n_179),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_237),
.A2(n_205),
.B(n_189),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_208),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_239),
.Y(n_247)
);

AOI22x1_ASAP7_75t_L g242 ( 
.A1(n_204),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_189),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_191),
.B(n_8),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_241),
.Y(n_244)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_248),
.C(n_260),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_193),
.C(n_203),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_241),
.Y(n_249)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

INVx13_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_207),
.Y(n_253)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_253),
.Y(n_278)
);

AOI211xp5_ASAP7_75t_SL g277 ( 
.A1(n_254),
.A2(n_242),
.B(n_237),
.C(n_243),
.Y(n_277)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_224),
.Y(n_256)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_256),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_194),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_257),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_230),
.A2(n_205),
.B1(n_210),
.B2(n_211),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_258),
.A2(n_263),
.B(n_264),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_222),
.B(n_193),
.C(n_200),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_220),
.A2(n_198),
.B1(n_211),
.B2(n_209),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_231),
.Y(n_267)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_223),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_273),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_272),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_232),
.C(n_234),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_264),
.C(n_262),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_259),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_231),
.Y(n_273)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_225),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_261),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_245),
.B(n_240),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_281),
.B(n_228),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_285),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_270),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_235),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_287),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_282),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_291),
.Y(n_301)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_265),
.C(n_267),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_250),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_294),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_276),
.A2(n_246),
.B1(n_252),
.B2(n_247),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_258),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_296),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_269),
.A2(n_247),
.B1(n_226),
.B2(n_239),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_266),
.A2(n_254),
.B(n_242),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_297),
.A2(n_277),
.B(n_273),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_292),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_299),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_302),
.B(n_8),
.Y(n_314)
);

INVx11_ASAP7_75t_L g303 ( 
.A(n_287),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_303),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g305 ( 
.A(n_288),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_307),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_285),
.A2(n_271),
.B1(n_280),
.B2(n_275),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_283),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_289),
.B(n_279),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_6),
.C(n_13),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_307),
.A2(n_283),
.B(n_290),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_310),
.A2(n_301),
.B(n_317),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_300),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_298),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_305),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_289),
.C(n_272),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_313),
.B(n_314),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_306),
.C(n_304),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_321),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_303),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_323),
.A2(n_324),
.B(n_316),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_316),
.A2(n_313),
.B(n_318),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_325),
.A2(n_327),
.B(n_319),
.Y(n_328)
);

AOI322xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_326),
.A3(n_9),
.B1(n_5),
.B2(n_11),
.C1(n_13),
.C2(n_14),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_329),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_330),
.Y(n_331)
);

A2O1A1O1Ixp25_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_9),
.B(n_3),
.C(n_4),
.D(n_2),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_3),
.Y(n_333)
);

OAI311xp33_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_4),
.A3(n_9),
.B1(n_305),
.C1(n_316),
.Y(n_334)
);


endmodule