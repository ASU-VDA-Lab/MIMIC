module fake_jpeg_5779_n_140 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_140);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx3_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_30),
.Y(n_39)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_33),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

CKINVDCx6p67_ASAP7_75t_R g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_0),
.Y(n_33)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_25),
.Y(n_34)
);

INVx5_ASAP7_75t_SL g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_22),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_28),
.A2(n_18),
.B1(n_13),
.B2(n_19),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_19),
.B1(n_13),
.B2(n_21),
.Y(n_60)
);

NAND3xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_26),
.C(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_45),
.B(n_17),
.Y(n_66)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_44),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_51),
.Y(n_73)
);

OAI32xp33_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_34),
.A3(n_32),
.B1(n_28),
.B2(n_29),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_56),
.Y(n_72)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_54),
.B(n_63),
.Y(n_69)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_21),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_40),
.B(n_33),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_58),
.Y(n_78)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_61),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_60),
.A2(n_41),
.B(n_34),
.Y(n_68)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_65),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_26),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_14),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_66),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_35),
.Y(n_67)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_82),
.B1(n_59),
.B2(n_51),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_56),
.A2(n_47),
.B(n_38),
.C(n_30),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_70),
.B(n_71),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_47),
.B(n_38),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_15),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_47),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_83),
.B1(n_61),
.B2(n_53),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_30),
.B1(n_46),
.B2(n_36),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_27),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_54),
.A2(n_36),
.B(n_27),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_84),
.Y(n_98)
);

FAx1_ASAP7_75t_SL g106 ( 
.A(n_85),
.B(n_69),
.CI(n_75),
.CON(n_106),
.SN(n_106)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_92),
.B1(n_83),
.B2(n_98),
.Y(n_99)
);

NOR2x1p5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_62),
.Y(n_87)
);

AO21x1_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_70),
.B(n_84),
.Y(n_105)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_89),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_80),
.Y(n_89)
);

OA21x2_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_65),
.B(n_22),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_93),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_73),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_91),
.B(n_95),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_72),
.A2(n_48),
.B1(n_15),
.B2(n_7),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_94),
.A2(n_97),
.B(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_75),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_96),
.B(n_77),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_106),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_76),
.B1(n_78),
.B2(n_83),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_78),
.B1(n_69),
.B2(n_68),
.Y(n_101)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_107),
.B(n_109),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_95),
.A2(n_81),
.B(n_48),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_103),
.B(n_88),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_117),
.B(n_0),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_85),
.C(n_92),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_115),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_90),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_108),
.A2(n_90),
.B1(n_89),
.B2(n_93),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_116),
.A2(n_106),
.B1(n_3),
.B2(n_4),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_0),
.C(n_1),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_112),
.A2(n_102),
.B(n_105),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_122),
.Y(n_128)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_114),
.A2(n_106),
.B1(n_3),
.B2(n_5),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_120),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_121),
.B(n_117),
.Y(n_124)
);

INVxp33_ASAP7_75t_SL g122 ( 
.A(n_116),
.Y(n_122)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_113),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_123),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_129),
.B(n_125),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_128),
.A2(n_122),
.B1(n_113),
.B2(n_115),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_130),
.A2(n_131),
.B(n_10),
.C(n_11),
.Y(n_135)
);

OAI31xp33_ASAP7_75t_L g131 ( 
.A1(n_128),
.A2(n_111),
.A3(n_6),
.B(n_9),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_134),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_132),
.A2(n_127),
.B1(n_126),
.B2(n_11),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_135),
.A2(n_10),
.B(n_12),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_5),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_136),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_130),
.Y(n_140)
);


endmodule