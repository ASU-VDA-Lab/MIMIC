module fake_jpeg_17275_n_149 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_149);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_149;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_36),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_38),
.B(n_39),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_14),
.B(n_1),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_24),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_30),
.B1(n_26),
.B2(n_20),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_44),
.A2(n_48),
.B1(n_52),
.B2(n_61),
.Y(n_77)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_26),
.B1(n_20),
.B2(n_14),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_49),
.B(n_6),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_33),
.A2(n_15),
.B1(n_22),
.B2(n_29),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_15),
.B1(n_22),
.B2(n_29),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_54),
.A2(n_58),
.B1(n_62),
.B2(n_43),
.Y(n_71)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_41),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_31),
.B1(n_32),
.B2(n_24),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_31),
.A2(n_25),
.B1(n_23),
.B2(n_21),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_32),
.A2(n_23),
.B1(n_21),
.B2(n_18),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_47),
.B(n_49),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_69),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_70),
.Y(n_87)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_42),
.B1(n_18),
.B2(n_16),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_47),
.B(n_38),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_74),
.Y(n_88)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_67),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_40),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_63),
.Y(n_85)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_80),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_79),
.B1(n_7),
.B2(n_8),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_45),
.B(n_7),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_82),
.Y(n_91)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_59),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_53),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_63),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_56),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_56),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_92),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_74),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_95),
.B(n_65),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_55),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_96),
.B(n_8),
.Y(n_104)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

NOR2xp67_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_71),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_107),
.B(n_84),
.Y(n_121)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_104),
.B1(n_96),
.B2(n_88),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_93),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_112),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_82),
.C(n_63),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_108),
.C(n_111),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_75),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_110),
.B(n_113),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_75),
.C(n_40),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_90),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_87),
.B(n_60),
.Y(n_113)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_100),
.A2(n_94),
.B1(n_95),
.B2(n_97),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_102),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_117),
.B(n_99),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_112),
.A2(n_94),
.B(n_95),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_120),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_111),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_123),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_99),
.B1(n_72),
.B2(n_83),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_125),
.B(n_122),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_108),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_127),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_120),
.C(n_105),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_109),
.C(n_102),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_118),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_124),
.A2(n_115),
.B(n_123),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_132),
.A2(n_134),
.B(n_130),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_135),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_124),
.A2(n_115),
.B(n_117),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_103),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_126),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_140),
.C(n_128),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_141),
.A2(n_106),
.B1(n_128),
.B2(n_101),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_139),
.B(n_91),
.Y(n_142)
);

NAND3xp33_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_143),
.C(n_13),
.Y(n_146)
);

AOI322xp5_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_116),
.A3(n_106),
.B1(n_89),
.B2(n_59),
.C1(n_13),
.C2(n_11),
.Y(n_145)
);

INVxp33_ASAP7_75t_L g147 ( 
.A(n_145),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_147),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_146),
.Y(n_149)
);


endmodule