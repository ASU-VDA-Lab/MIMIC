module fake_netlist_1_1780_n_35 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_35);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_35;
wire n_20;
wire n_34;
wire n_28;
wire n_8;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_6), .Y(n_8) );
BUFx3_ASAP7_75t_L g9 ( .A(n_1), .Y(n_9) );
AND2x6_ASAP7_75t_L g10 ( .A(n_7), .B(n_3), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_5), .Y(n_11) );
NAND2xp33_ASAP7_75t_SL g12 ( .A(n_4), .B(n_3), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_4), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_11), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_9), .Y(n_15) );
BUFx3_ASAP7_75t_L g16 ( .A(n_10), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_13), .B(n_2), .Y(n_17) );
NOR2xp33_ASAP7_75t_R g18 ( .A(n_8), .B(n_0), .Y(n_18) );
AOI21x1_ASAP7_75t_L g19 ( .A1(n_14), .A2(n_10), .B(n_12), .Y(n_19) );
NAND3xp33_ASAP7_75t_L g20 ( .A(n_17), .B(n_12), .C(n_10), .Y(n_20) );
INVx5_ASAP7_75t_L g21 ( .A(n_14), .Y(n_21) );
CKINVDCx14_ASAP7_75t_R g22 ( .A(n_18), .Y(n_22) );
OAI22xp33_ASAP7_75t_L g23 ( .A1(n_20), .A2(n_15), .B1(n_16), .B2(n_10), .Y(n_23) );
INVxp33_ASAP7_75t_SL g24 ( .A(n_22), .Y(n_24) );
INVxp67_ASAP7_75t_L g25 ( .A(n_19), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_25), .B(n_21), .Y(n_26) );
AND2x2_ASAP7_75t_L g27 ( .A(n_25), .B(n_15), .Y(n_27) );
CKINVDCx5p33_ASAP7_75t_R g28 ( .A(n_27), .Y(n_28) );
NOR2xp33_ASAP7_75t_L g29 ( .A(n_26), .B(n_24), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
NAND2xp5_ASAP7_75t_L g31 ( .A(n_29), .B(n_23), .Y(n_31) );
AOI22xp33_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_21), .B1(n_16), .B2(n_2), .Y(n_32) );
NAND2x1p5_ASAP7_75t_L g33 ( .A(n_31), .B(n_21), .Y(n_33) );
AND2x2_ASAP7_75t_SL g34 ( .A(n_32), .B(n_0), .Y(n_34) );
AOI22xp33_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_1), .B1(n_33), .B2(n_31), .Y(n_35) );
endmodule