module real_aes_14461_n_9 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_1, n_9);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_1;
output n_9;
wire n_17;
wire n_28;
wire n_22;
wire n_13;
wire n_24;
wire n_41;
wire n_34;
wire n_12;
wire n_19;
wire n_40;
wire n_25;
wire n_32;
wire n_30;
wire n_14;
wire n_11;
wire n_16;
wire n_37;
wire n_35;
wire n_39;
wire n_15;
wire n_27;
wire n_23;
wire n_38;
wire n_29;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_10;
wire n_33;
wire n_36;
BUFx10_ASAP7_75t_L g29 ( .A(n_0), .Y(n_29) );
INVx1_ASAP7_75t_L g31 ( .A(n_1), .Y(n_31) );
INVx2_ASAP7_75t_L g36 ( .A(n_2), .Y(n_36) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_3), .Y(n_17) );
AOI21xp33_ASAP7_75t_L g9 ( .A1(n_4), .A2(n_10), .B(n_22), .Y(n_9) );
NAND3xp33_ASAP7_75t_L g12 ( .A(n_5), .B(n_13), .C(n_16), .Y(n_12) );
BUFx3_ASAP7_75t_L g34 ( .A(n_6), .Y(n_34) );
INVx3_ASAP7_75t_L g15 ( .A(n_7), .Y(n_15) );
INVx1_ASAP7_75t_L g21 ( .A(n_8), .Y(n_21) );
INVxp33_ASAP7_75t_L g10 ( .A(n_11), .Y(n_10) );
NOR2xp33_ASAP7_75t_SL g11 ( .A(n_12), .B(n_18), .Y(n_11) );
BUFx3_ASAP7_75t_L g13 ( .A(n_14), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_15), .Y(n_14) );
INVx1_ASAP7_75t_L g16 ( .A(n_17), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_17), .B(n_25), .Y(n_24) );
INVx1_ASAP7_75t_L g18 ( .A(n_19), .Y(n_18) );
BUFx2_ASAP7_75t_L g19 ( .A(n_20), .Y(n_19) );
INVx1_ASAP7_75t_L g25 ( .A(n_20), .Y(n_25) );
HB1xp67_ASAP7_75t_L g20 ( .A(n_21), .Y(n_20) );
AND2x2_ASAP7_75t_L g22 ( .A(n_23), .B(n_26), .Y(n_22) );
INVxp67_ASAP7_75t_L g23 ( .A(n_24), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_27), .B(n_37), .Y(n_26) );
NAND3xp33_ASAP7_75t_L g27 ( .A(n_28), .B(n_30), .C(n_32), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_29), .Y(n_28) );
AND2x4_ASAP7_75t_L g38 ( .A(n_30), .B(n_39), .Y(n_38) );
INVx1_ASAP7_75t_L g30 ( .A(n_31), .Y(n_30) );
BUFx6f_ASAP7_75t_L g32 ( .A(n_33), .Y(n_32) );
OR2x2_ASAP7_75t_L g33 ( .A(n_34), .B(n_35), .Y(n_33) );
AND2x2_ASAP7_75t_L g41 ( .A(n_34), .B(n_35), .Y(n_41) );
INVx1_ASAP7_75t_L g35 ( .A(n_36), .Y(n_35) );
INVx2_ASAP7_75t_SL g37 ( .A(n_38), .Y(n_37) );
INVx1_ASAP7_75t_L g39 ( .A(n_40), .Y(n_39) );
INVx1_ASAP7_75t_L g40 ( .A(n_41), .Y(n_40) );
endmodule