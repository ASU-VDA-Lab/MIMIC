module fake_jpeg_14446_n_183 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_183);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_183;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_10),
.B(n_6),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_11),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_36),
.B(n_50),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_46),
.Y(n_57)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_23),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_47),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

OR2x4_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_11),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_52),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_51),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_22),
.B(n_0),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_15),
.B(n_7),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_54),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_69),
.Y(n_91)
);

NOR2x1_ASAP7_75t_R g58 ( 
.A(n_40),
.B(n_21),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_58),
.B(n_59),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_39),
.A2(n_29),
.B1(n_17),
.B2(n_18),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_62),
.A2(n_74),
.B1(n_75),
.B2(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_14),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_63),
.B(n_64),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_34),
.B(n_14),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_53),
.A2(n_29),
.B1(n_17),
.B2(n_18),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_71),
.B1(n_81),
.B2(n_76),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_83),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_15),
.B1(n_31),
.B2(n_19),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_44),
.A2(n_19),
.B1(n_2),
.B2(n_3),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_34),
.B(n_8),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_77),
.B(n_79),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_33),
.B(n_1),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_35),
.B(n_4),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_47),
.A2(n_4),
.B1(n_5),
.B2(n_41),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_84),
.A2(n_81),
.B(n_80),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_43),
.B(n_5),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_85),
.B(n_80),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_50),
.A2(n_5),
.B1(n_22),
.B2(n_16),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_88),
.A2(n_102),
.B1(n_61),
.B2(n_72),
.Y(n_123)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_91),
.B(n_94),
.Y(n_120)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_71),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_SL g95 ( 
.A1(n_58),
.A2(n_71),
.B(n_55),
.C(n_67),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_59),
.B(n_56),
.C(n_82),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_76),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_97),
.B(n_78),
.Y(n_125)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_84),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_82),
.Y(n_112)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_108),
.Y(n_110)
);

INVx3_ASAP7_75t_SL g107 ( 
.A(n_73),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_109),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_112),
.B(n_122),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_73),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_102),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_56),
.B(n_106),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_78),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_123),
.A2(n_98),
.B1(n_109),
.B2(n_104),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_127),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_72),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_96),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_87),
.Y(n_137)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_130),
.B(n_131),
.Y(n_153)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_116),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_134),
.Y(n_154)
);

AO22x1_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_95),
.B1(n_109),
.B2(n_92),
.Y(n_135)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_137),
.B(n_139),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_103),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_143),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_93),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

AOI32xp33_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_107),
.A3(n_105),
.B1(n_90),
.B2(n_56),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_141),
.B(n_124),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_110),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_138),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_132),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_149),
.A2(n_153),
.B(n_131),
.Y(n_160)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_144),
.C(n_135),
.Y(n_165)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_156),
.B(n_157),
.Y(n_166)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_143),
.C(n_136),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_162),
.C(n_163),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_SL g159 ( 
.A1(n_150),
.A2(n_142),
.B(n_135),
.C(n_130),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_160),
.B(n_152),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_161),
.A2(n_148),
.B1(n_151),
.B2(n_154),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_124),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_124),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_155),
.B(n_111),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_165),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_167),
.A2(n_161),
.B1(n_151),
.B2(n_145),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_169),
.A2(n_152),
.B(n_159),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_171),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_159),
.C(n_134),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_172),
.B(n_173),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_117),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_174),
.A2(n_166),
.B(n_140),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_177),
.A2(n_173),
.B(n_172),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_178),
.B(n_179),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_175),
.A2(n_133),
.B(n_129),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_176),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_114),
.B1(n_121),
.B2(n_126),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_182),
.A2(n_119),
.B(n_114),
.Y(n_183)
);


endmodule