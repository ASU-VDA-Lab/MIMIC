module real_aes_18339_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1225;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_1404;
wire n_402;
wire n_602;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_265;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1403;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1431;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_1085;
wire n_276;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_1049;
wire n_559;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_1352;
wire n_729;
wire n_1280;
wire n_1323;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_SL g883 ( .A1(n_0), .A2(n_67), .B1(n_485), .B2(n_487), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_0), .A2(n_229), .B1(n_587), .B2(n_633), .Y(n_894) );
OAI211xp5_ASAP7_75t_L g1361 ( .A1(n_1), .A2(n_1356), .B(n_1362), .C(n_1363), .Y(n_1361) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1), .Y(n_1383) );
INVx1_ASAP7_75t_L g889 ( .A(n_2), .Y(n_889) );
OAI211xp5_ASAP7_75t_L g442 ( .A1(n_3), .A2(n_443), .B(n_445), .C(n_456), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_3), .B(n_477), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g1405 ( .A1(n_4), .A2(n_114), .B1(n_1406), .B2(n_1408), .Y(n_1405) );
AOI22xp33_ASAP7_75t_SL g1424 ( .A1(n_4), .A2(n_116), .B1(n_586), .B2(n_633), .Y(n_1424) );
AOI22xp5_ASAP7_75t_SL g1138 ( .A1(n_5), .A2(n_232), .B1(n_1131), .B2(n_1139), .Y(n_1138) );
INVx1_ASAP7_75t_L g297 ( .A(n_6), .Y(n_297) );
AO22x1_ASAP7_75t_L g371 ( .A1(n_6), .A2(n_131), .B1(n_372), .B2(n_374), .Y(n_371) );
AND2x2_ASAP7_75t_L g266 ( .A(n_7), .B(n_267), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_7), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g383 ( .A(n_7), .B(n_206), .Y(n_383) );
INVx1_ASAP7_75t_L g402 ( .A(n_7), .Y(n_402) );
INVx1_ASAP7_75t_L g318 ( .A(n_8), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_8), .A2(n_95), .B1(n_367), .B2(n_369), .Y(n_366) );
INVx1_ASAP7_75t_L g759 ( .A(n_9), .Y(n_759) );
AOI221xp5_ASAP7_75t_L g881 ( .A1(n_10), .A2(n_135), .B1(n_669), .B2(n_878), .C(n_882), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_10), .A2(n_58), .B1(n_587), .B2(n_898), .Y(n_897) );
AOI22xp33_ASAP7_75t_SL g1403 ( .A1(n_11), .A2(n_145), .B1(n_339), .B2(n_1404), .Y(n_1403) );
AOI221xp5_ASAP7_75t_L g1421 ( .A1(n_11), .A2(n_17), .B1(n_577), .B2(n_583), .C(n_1422), .Y(n_1421) );
AOI22xp33_ASAP7_75t_SL g539 ( .A1(n_12), .A2(n_118), .B1(n_482), .B2(n_540), .Y(n_539) );
INVxp67_ASAP7_75t_SL g607 ( .A(n_12), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_13), .A2(n_140), .B1(n_920), .B2(n_922), .Y(n_919) );
AOI22xp33_ASAP7_75t_SL g956 ( .A1(n_13), .A2(n_234), .B1(n_482), .B2(n_957), .Y(n_956) );
CKINVDCx5p33_ASAP7_75t_R g874 ( .A(n_14), .Y(n_874) );
CKINVDCx5p33_ASAP7_75t_R g1076 ( .A(n_15), .Y(n_1076) );
INVx2_ASAP7_75t_L g1126 ( .A(n_16), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_16), .B(n_1127), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1134 ( .A(n_16), .B(n_98), .Y(n_1134) );
AOI22xp33_ASAP7_75t_SL g1412 ( .A1(n_17), .A2(n_32), .B1(n_554), .B2(n_877), .Y(n_1412) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_18), .A2(n_220), .B1(n_540), .B2(n_552), .Y(n_551) );
AOI221xp5_ASAP7_75t_L g576 ( .A1(n_18), .A2(n_118), .B1(n_577), .B2(n_579), .C(n_582), .Y(n_576) );
INVx1_ASAP7_75t_L g1401 ( .A(n_19), .Y(n_1401) );
OAI22xp33_ASAP7_75t_L g1413 ( .A1(n_20), .A2(n_193), .B1(n_556), .B2(n_560), .Y(n_1413) );
INVx1_ASAP7_75t_L g1427 ( .A(n_20), .Y(n_1427) );
XNOR2xp5_ASAP7_75t_L g623 ( .A(n_21), .B(n_624), .Y(n_623) );
AOI22xp5_ASAP7_75t_SL g1153 ( .A1(n_21), .A2(n_122), .B1(n_1131), .B2(n_1139), .Y(n_1153) );
INVx1_ASAP7_75t_L g1081 ( .A(n_22), .Y(n_1081) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_23), .A2(n_211), .B1(n_417), .B2(n_569), .Y(n_568) );
XOR2x2_ASAP7_75t_L g747 ( .A(n_24), .B(n_748), .Y(n_747) );
AOI22xp5_ASAP7_75t_SL g1143 ( .A1(n_25), .A2(n_226), .B1(n_1128), .B2(n_1133), .Y(n_1143) );
INVx1_ASAP7_75t_L g914 ( .A(n_26), .Y(n_914) );
OAI22xp5_ASAP7_75t_L g939 ( .A1(n_26), .A2(n_222), .B1(n_417), .B2(n_569), .Y(n_939) );
INVx1_ASAP7_75t_L g1026 ( .A(n_27), .Y(n_1026) );
OAI22xp33_ASAP7_75t_L g1044 ( .A1(n_27), .A2(n_154), .B1(n_556), .B2(n_960), .Y(n_1044) );
OAI221xp5_ASAP7_75t_L g1034 ( .A1(n_28), .A2(n_52), .B1(n_597), .B2(n_1003), .C(n_1035), .Y(n_1034) );
INVx1_ASAP7_75t_L g1052 ( .A(n_28), .Y(n_1052) );
OAI211xp5_ASAP7_75t_L g457 ( .A1(n_29), .A2(n_458), .B(n_462), .C(n_464), .Y(n_457) );
INVx1_ASAP7_75t_L g520 ( .A(n_29), .Y(n_520) );
CKINVDCx5p33_ASAP7_75t_R g966 ( .A(n_30), .Y(n_966) );
OAI22xp33_ASAP7_75t_L g1359 ( .A1(n_31), .A2(n_163), .B1(n_822), .B2(n_1360), .Y(n_1359) );
OAI22xp33_ASAP7_75t_L g1373 ( .A1(n_31), .A2(n_163), .B1(n_834), .B2(n_1374), .Y(n_1373) );
A2O1A1Ixp33_ASAP7_75t_L g1430 ( .A1(n_32), .A2(n_1342), .B(n_1431), .C(n_1438), .Y(n_1430) );
AOI22xp5_ASAP7_75t_L g1122 ( .A1(n_33), .A2(n_157), .B1(n_1123), .B2(n_1128), .Y(n_1122) );
INVx1_ASAP7_75t_L g1337 ( .A(n_34), .Y(n_1337) );
INVx1_ASAP7_75t_L g776 ( .A(n_35), .Y(n_776) );
OAI22xp5_ASAP7_75t_L g1417 ( .A1(n_36), .A2(n_57), .B1(n_477), .B2(n_569), .Y(n_1417) );
OAI211xp5_ASAP7_75t_L g1419 ( .A1(n_36), .A2(n_995), .B(n_1420), .C(n_1425), .Y(n_1419) );
AOI22xp33_ASAP7_75t_L g1220 ( .A1(n_37), .A2(n_90), .B1(n_1131), .B2(n_1149), .Y(n_1220) );
INVx1_ASAP7_75t_L g740 ( .A(n_38), .Y(n_740) );
XOR2x2_ASAP7_75t_L g528 ( .A(n_39), .B(n_529), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g1130 ( .A1(n_39), .A2(n_160), .B1(n_1131), .B2(n_1133), .Y(n_1130) );
AOI21xp33_ASAP7_75t_L g644 ( .A1(n_40), .A2(n_645), .B(n_646), .Y(n_644) );
INVx1_ASAP7_75t_L g656 ( .A(n_40), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g1161 ( .A1(n_41), .A2(n_76), .B1(n_1123), .B2(n_1131), .Y(n_1161) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_42), .A2(n_63), .B1(n_409), .B2(n_447), .Y(n_446) );
AOI22xp33_ASAP7_75t_SL g481 ( .A1(n_42), .A2(n_243), .B1(n_482), .B2(n_483), .Y(n_481) );
INVx1_ASAP7_75t_L g991 ( .A(n_43), .Y(n_991) );
INVx1_ASAP7_75t_L g289 ( .A(n_44), .Y(n_289) );
INVx1_ASAP7_75t_L g302 ( .A(n_44), .Y(n_302) );
INVx1_ASAP7_75t_L g1327 ( .A(n_45), .Y(n_1327) );
INVxp67_ASAP7_75t_SL g1017 ( .A(n_46), .Y(n_1017) );
AND4x1_ASAP7_75t_L g1054 ( .A(n_46), .B(n_1019), .C(n_1022), .D(n_1042), .Y(n_1054) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_47), .A2(n_181), .B1(n_409), .B2(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g657 ( .A(n_47), .Y(n_657) );
OAI22xp33_ASAP7_75t_L g555 ( .A1(n_48), .A2(n_158), .B1(n_556), .B2(n_560), .Y(n_555) );
INVx1_ASAP7_75t_L g590 ( .A(n_48), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g1165 ( .A1(n_49), .A2(n_241), .B1(n_1123), .B2(n_1128), .Y(n_1165) );
INVxp67_ASAP7_75t_SL g929 ( .A(n_50), .Y(n_929) );
AOI22xp33_ASAP7_75t_SL g953 ( .A1(n_50), .A2(n_117), .B1(n_545), .B2(n_954), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g1409 ( .A1(n_51), .A2(n_116), .B1(n_1408), .B2(n_1410), .Y(n_1409) );
AOI221xp5_ASAP7_75t_L g1432 ( .A1(n_51), .A2(n_114), .B1(n_1433), .B2(n_1435), .C(n_1436), .Y(n_1432) );
INVx1_ASAP7_75t_L g1053 ( .A(n_52), .Y(n_1053) );
INVx1_ASAP7_75t_L g1108 ( .A(n_53), .Y(n_1108) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_54), .A2(n_212), .B1(n_583), .B2(n_629), .C(n_630), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_54), .A2(n_246), .B1(n_482), .B2(n_501), .Y(n_662) );
INVx2_ASAP7_75t_L g285 ( .A(n_55), .Y(n_285) );
INVx1_ASAP7_75t_L g426 ( .A(n_56), .Y(n_426) );
AOI221xp5_ASAP7_75t_L g876 ( .A1(n_58), .A2(n_66), .B1(n_877), .B2(n_878), .C(n_879), .Y(n_876) );
NOR2xp33_ASAP7_75t_L g934 ( .A(n_59), .B(n_638), .Y(n_934) );
INVx1_ASAP7_75t_L g945 ( .A(n_59), .Y(n_945) );
AOI22xp5_ASAP7_75t_L g1144 ( .A1(n_60), .A2(n_65), .B1(n_1123), .B2(n_1131), .Y(n_1144) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_61), .A2(n_74), .B1(n_981), .B2(n_983), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_61), .A2(n_208), .B1(n_423), .B2(n_920), .Y(n_998) );
INVx1_ASAP7_75t_L g870 ( .A(n_62), .Y(n_870) );
AOI22xp33_ASAP7_75t_SL g490 ( .A1(n_63), .A2(n_94), .B1(n_342), .B2(n_482), .Y(n_490) );
INVx1_ASAP7_75t_L g869 ( .A(n_64), .Y(n_869) );
AOI221xp5_ASAP7_75t_L g893 ( .A1(n_66), .A2(n_135), .B1(n_455), .B2(n_578), .C(n_580), .Y(n_893) );
AOI221xp5_ASAP7_75t_L g899 ( .A1(n_67), .A2(n_69), .B1(n_580), .B2(n_618), .C(n_629), .Y(n_899) );
AOI22xp33_ASAP7_75t_SL g1067 ( .A1(n_68), .A2(n_167), .B1(n_540), .B2(n_1068), .Y(n_1067) );
AOI22xp33_ASAP7_75t_SL g1097 ( .A1(n_68), .A2(n_215), .B1(n_633), .B2(n_1033), .Y(n_1097) );
AOI22xp33_ASAP7_75t_SL g880 ( .A1(n_69), .A2(n_229), .B1(n_485), .B2(n_487), .Y(n_880) );
AOI22xp5_ASAP7_75t_L g1160 ( .A1(n_70), .A2(n_173), .B1(n_1128), .B2(n_1139), .Y(n_1160) );
OAI22xp5_ASAP7_75t_L g1021 ( .A1(n_71), .A2(n_189), .B1(n_417), .B2(n_569), .Y(n_1021) );
OAI211xp5_ASAP7_75t_L g1023 ( .A1(n_71), .A2(n_995), .B(n_1024), .C(n_1027), .Y(n_1023) );
OAI222xp33_ASAP7_75t_L g337 ( .A1(n_72), .A2(n_186), .B1(n_338), .B2(n_346), .C1(n_348), .C2(n_352), .Y(n_337) );
INVx1_ASAP7_75t_L g384 ( .A(n_72), .Y(n_384) );
INVx1_ASAP7_75t_L g1366 ( .A(n_73), .Y(n_1366) );
OAI211xp5_ASAP7_75t_L g1375 ( .A1(n_73), .A2(n_1376), .B(n_1377), .C(n_1381), .Y(n_1375) );
AOI21xp33_ASAP7_75t_L g1006 ( .A1(n_74), .A2(n_449), .B(n_454), .Y(n_1006) );
OAI211xp5_ASAP7_75t_L g806 ( .A1(n_75), .A2(n_789), .B(n_807), .C(n_809), .Y(n_806) );
INVx1_ASAP7_75t_L g856 ( .A(n_75), .Y(n_856) );
INVx1_ASAP7_75t_L g536 ( .A(n_77), .Y(n_536) );
OAI221xp5_ASAP7_75t_L g596 ( .A1(n_77), .A2(n_86), .B1(n_597), .B2(n_601), .C(n_604), .Y(n_596) );
OAI22xp33_ASAP7_75t_L g992 ( .A1(n_78), .A2(n_82), .B1(n_560), .B2(n_959), .Y(n_992) );
INVx1_ASAP7_75t_L g1000 ( .A(n_78), .Y(n_1000) );
INVx1_ASAP7_75t_L g1340 ( .A(n_79), .Y(n_1340) );
INVx1_ASAP7_75t_L g1339 ( .A(n_80), .Y(n_1339) );
AOI22xp33_ASAP7_75t_SL g987 ( .A1(n_81), .A2(n_237), .B1(n_877), .B2(n_976), .Y(n_987) );
AOI22xp33_ASAP7_75t_SL g1007 ( .A1(n_81), .A2(n_156), .B1(n_1008), .B2(n_1009), .Y(n_1007) );
INVx1_ASAP7_75t_L g1001 ( .A(n_82), .Y(n_1001) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_83), .Y(n_309) );
XOR2xp5_ASAP7_75t_L g1393 ( .A(n_84), .B(n_1394), .Y(n_1393) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_85), .A2(n_239), .B1(n_372), .B2(n_1033), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g1049 ( .A1(n_85), .A2(n_107), .B1(n_545), .B2(n_1048), .Y(n_1049) );
INVx1_ASAP7_75t_L g533 ( .A(n_86), .Y(n_533) );
INVx1_ASAP7_75t_L g699 ( .A(n_87), .Y(n_699) );
AOI221xp5_ASAP7_75t_L g719 ( .A1(n_87), .A2(n_200), .B1(n_669), .B2(n_720), .C(n_721), .Y(n_719) );
AOI22xp33_ASAP7_75t_SL g1070 ( .A1(n_88), .A2(n_248), .B1(n_717), .B2(n_954), .Y(n_1070) );
AOI21xp33_ASAP7_75t_L g1094 ( .A1(n_88), .A2(n_618), .B(n_1095), .Y(n_1094) );
HB1xp67_ASAP7_75t_L g1110 ( .A(n_89), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1124 ( .A(n_89), .B(n_1108), .Y(n_1124) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_91), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g873 ( .A(n_92), .Y(n_873) );
AOI22xp5_ASAP7_75t_L g1147 ( .A1(n_93), .A2(n_147), .B1(n_1123), .B2(n_1128), .Y(n_1147) );
AOI221xp5_ASAP7_75t_SL g453 ( .A1(n_94), .A2(n_243), .B1(n_369), .B2(n_454), .C(n_455), .Y(n_453) );
INVx1_ASAP7_75t_L g312 ( .A(n_95), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g641 ( .A(n_96), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g1082 ( .A1(n_97), .A2(n_235), .B1(n_560), .B2(n_959), .Y(n_1082) );
INVx1_ASAP7_75t_L g1089 ( .A(n_97), .Y(n_1089) );
INVx1_ASAP7_75t_L g1127 ( .A(n_98), .Y(n_1127) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_98), .B(n_1126), .Y(n_1132) );
AOI22xp5_ASAP7_75t_L g1140 ( .A1(n_99), .A2(n_172), .B1(n_1123), .B2(n_1128), .Y(n_1140) );
OAI22xp33_ASAP7_75t_L g735 ( .A1(n_100), .A2(n_209), .B1(n_281), .B2(n_736), .Y(n_735) );
INVxp67_ASAP7_75t_SL g739 ( .A(n_100), .Y(n_739) );
INVxp67_ASAP7_75t_SL g1038 ( .A(n_101), .Y(n_1038) );
AOI22xp33_ASAP7_75t_SL g1050 ( .A1(n_101), .A2(n_191), .B1(n_723), .B2(n_957), .Y(n_1050) );
CKINVDCx5p33_ASAP7_75t_R g469 ( .A(n_102), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g1020 ( .A(n_103), .Y(n_1020) );
INVx1_ASAP7_75t_L g815 ( .A(n_104), .Y(n_815) );
OAI211xp5_ASAP7_75t_L g849 ( .A1(n_104), .A2(n_756), .B(n_850), .C(n_853), .Y(n_849) );
INVxp67_ASAP7_75t_SL g926 ( .A(n_105), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_105), .A2(n_233), .B1(n_950), .B2(n_951), .Y(n_949) );
OAI211xp5_ASAP7_75t_SL g915 ( .A1(n_106), .A2(n_601), .B(n_916), .C(n_925), .Y(n_915) );
INVx1_ASAP7_75t_L g943 ( .A(n_106), .Y(n_943) );
AOI221xp5_ASAP7_75t_L g1039 ( .A1(n_107), .A2(n_202), .B1(n_367), .B2(n_618), .C(n_1040), .Y(n_1039) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_108), .B(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g315 ( .A(n_108), .Y(n_315) );
INVx1_ASAP7_75t_L g331 ( .A(n_108), .Y(n_331) );
OAI22xp33_ASAP7_75t_L g1367 ( .A1(n_109), .A2(n_217), .B1(n_1368), .B2(n_1369), .Y(n_1367) );
OAI22xp5_ASAP7_75t_L g1384 ( .A1(n_109), .A2(n_217), .B1(n_1385), .B2(n_1386), .Y(n_1384) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_110), .A2(n_126), .B1(n_458), .B2(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g499 ( .A(n_110), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_111), .A2(n_136), .B1(n_684), .B2(n_685), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_111), .A2(n_185), .B1(n_487), .B2(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g325 ( .A(n_112), .Y(n_325) );
NAND2xp33_ASAP7_75t_SL g410 ( .A(n_112), .B(n_369), .Y(n_410) );
INVx1_ASAP7_75t_L g705 ( .A(n_113), .Y(n_705) );
INVx1_ASAP7_75t_L g913 ( .A(n_115), .Y(n_913) );
OAI22xp33_ASAP7_75t_L g958 ( .A1(n_115), .A2(n_242), .B1(n_959), .B2(n_960), .Y(n_958) );
INVxp67_ASAP7_75t_SL g917 ( .A(n_117), .Y(n_917) );
INVx1_ASAP7_75t_L g752 ( .A(n_119), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_120), .A2(n_208), .B1(n_983), .B2(n_985), .Y(n_984) );
INVx1_ASAP7_75t_L g1005 ( .A(n_120), .Y(n_1005) );
INVx1_ASAP7_75t_L g775 ( .A(n_121), .Y(n_775) );
INVx1_ASAP7_75t_L g636 ( .A(n_123), .Y(n_636) );
INVxp67_ASAP7_75t_SL g1065 ( .A(n_124), .Y(n_1065) );
OAI211xp5_ASAP7_75t_L g1084 ( .A1(n_124), .A2(n_573), .B(n_1085), .C(n_1088), .Y(n_1084) );
AOI22xp33_ASAP7_75t_SL g1071 ( .A1(n_125), .A2(n_230), .B1(n_717), .B2(n_954), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1087 ( .A1(n_125), .A2(n_248), .B1(n_587), .B2(n_1008), .Y(n_1087) );
INVx1_ASAP7_75t_L g516 ( .A(n_126), .Y(n_516) );
INVx1_ASAP7_75t_L g1219 ( .A(n_127), .Y(n_1219) );
CKINVDCx16_ASAP7_75t_R g341 ( .A(n_128), .Y(n_341) );
INVx1_ASAP7_75t_L g1329 ( .A(n_129), .Y(n_1329) );
INVx1_ASAP7_75t_L g1333 ( .A(n_130), .Y(n_1333) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_131), .A2(n_327), .B(n_330), .Y(n_326) );
NAND5xp2_ASAP7_75t_L g440 ( .A(n_132), .B(n_441), .C(n_478), .D(n_502), .E(n_511), .Y(n_440) );
INVx1_ASAP7_75t_L g524 ( .A(n_132), .Y(n_524) );
INVx1_ASAP7_75t_L g415 ( .A(n_133), .Y(n_415) );
AOI22xp33_ASAP7_75t_SL g647 ( .A1(n_134), .A2(n_246), .B1(n_374), .B2(n_585), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_134), .A2(n_212), .B1(n_482), .B2(n_669), .Y(n_668) );
AOI22xp33_ASAP7_75t_SL g715 ( .A1(n_136), .A2(n_231), .B1(n_716), .B2(n_717), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_137), .A2(n_238), .B1(n_542), .B2(n_545), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_137), .A2(n_174), .B1(n_585), .B2(n_586), .Y(n_584) );
INVx1_ASAP7_75t_L g635 ( .A(n_138), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g1148 ( .A1(n_139), .A2(n_165), .B1(n_1131), .B2(n_1149), .Y(n_1148) );
AOI22xp33_ASAP7_75t_SL g947 ( .A1(n_140), .A2(n_159), .B1(n_482), .B2(n_948), .Y(n_947) );
BUFx3_ASAP7_75t_L g291 ( .A(n_141), .Y(n_291) );
INVx1_ASAP7_75t_L g1062 ( .A(n_142), .Y(n_1062) );
OAI221xp5_ASAP7_75t_L g1091 ( .A1(n_142), .A2(n_143), .B1(n_638), .B2(n_639), .C(n_1092), .Y(n_1091) );
INVx1_ASAP7_75t_L g1063 ( .A(n_143), .Y(n_1063) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_144), .A2(n_215), .B1(n_540), .B2(n_1073), .Y(n_1072) );
AOI221xp5_ASAP7_75t_L g1086 ( .A1(n_144), .A2(n_167), .B1(n_578), .B2(n_583), .C(n_645), .Y(n_1086) );
NAND2xp5_ASAP7_75t_L g1437 ( .A(n_145), .B(n_1326), .Y(n_1437) );
INVxp67_ASAP7_75t_L g964 ( .A(n_146), .Y(n_964) );
AOI22xp33_ASAP7_75t_SL g975 ( .A1(n_148), .A2(n_156), .B1(n_976), .B2(n_977), .Y(n_975) );
AOI221xp5_ASAP7_75t_L g997 ( .A1(n_148), .A2(n_237), .B1(n_367), .B2(n_583), .C(n_933), .Y(n_997) );
AOI22xp5_ASAP7_75t_L g1166 ( .A1(n_149), .A2(n_197), .B1(n_1131), .B2(n_1139), .Y(n_1166) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_150), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_151), .A2(n_184), .B1(n_372), .B2(n_409), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_151), .A2(n_179), .B1(n_487), .B2(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g891 ( .A(n_152), .Y(n_891) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_153), .A2(n_185), .B1(n_685), .B2(n_695), .C(n_697), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g718 ( .A1(n_153), .A2(n_192), .B1(n_330), .B2(n_482), .C(n_540), .Y(n_718) );
INVx1_ASAP7_75t_L g1025 ( .A(n_154), .Y(n_1025) );
OAI21xp5_ASAP7_75t_SL g901 ( .A1(n_155), .A2(n_675), .B(n_902), .Y(n_901) );
INVx1_ASAP7_75t_L g593 ( .A(n_158), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g930 ( .A1(n_159), .A2(n_234), .B1(n_583), .B2(n_931), .C(n_933), .Y(n_930) );
INVx1_ASAP7_75t_L g969 ( .A(n_161), .Y(n_969) );
OAI221xp5_ASAP7_75t_SL g1002 ( .A1(n_161), .A2(n_236), .B1(n_597), .B2(n_1003), .C(n_1004), .Y(n_1002) );
INVx1_ASAP7_75t_L g273 ( .A(n_162), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_162), .B(n_281), .Y(n_280) );
XOR2x2_ASAP7_75t_L g906 ( .A(n_164), .B(n_907), .Y(n_906) );
INVx1_ASAP7_75t_L g767 ( .A(n_166), .Y(n_767) );
INVx1_ASAP7_75t_L g1324 ( .A(n_168), .Y(n_1324) );
OAI221xp5_ASAP7_75t_L g637 ( .A1(n_169), .A2(n_214), .B1(n_638), .B2(n_639), .C(n_640), .Y(n_637) );
OAI22xp33_ASAP7_75t_L g670 ( .A1(n_169), .A2(n_214), .B1(n_535), .B2(n_671), .Y(n_670) );
OAI22xp33_ASAP7_75t_L g819 ( .A1(n_170), .A2(n_188), .B1(n_820), .B2(n_823), .Y(n_819) );
OAI22xp33_ASAP7_75t_L g831 ( .A1(n_170), .A2(n_188), .B1(n_832), .B2(n_837), .Y(n_831) );
INVx1_ASAP7_75t_L g754 ( .A(n_171), .Y(n_754) );
XOR2x2_ASAP7_75t_L g1317 ( .A(n_173), .B(n_1318), .Y(n_1317) );
AOI22xp33_ASAP7_75t_L g1388 ( .A1(n_173), .A2(n_1389), .B1(n_1392), .B2(n_1441), .Y(n_1388) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_174), .A2(n_244), .B1(n_542), .B2(n_545), .Y(n_541) );
INVx1_ASAP7_75t_L g510 ( .A(n_175), .Y(n_510) );
INVx1_ASAP7_75t_L g1365 ( .A(n_176), .Y(n_1365) );
INVxp67_ASAP7_75t_SL g1036 ( .A(n_177), .Y(n_1036) );
AOI22xp33_ASAP7_75t_SL g1046 ( .A1(n_177), .A2(n_201), .B1(n_554), .B2(n_948), .Y(n_1046) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_178), .Y(n_270) );
AOI221xp5_ASAP7_75t_L g448 ( .A1(n_179), .A2(n_223), .B1(n_367), .B2(n_369), .C(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g810 ( .A(n_180), .Y(n_810) );
INVx1_ASAP7_75t_L g667 ( .A(n_181), .Y(n_667) );
INVx1_ASAP7_75t_L g938 ( .A(n_182), .Y(n_938) );
CKINVDCx5p33_ASAP7_75t_R g1416 ( .A(n_183), .Y(n_1416) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_184), .A2(n_223), .B1(n_485), .B2(n_487), .Y(n_484) );
NOR2xp33_ASAP7_75t_R g392 ( .A(n_186), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g762 ( .A(n_187), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g1057 ( .A(n_190), .B(n_1058), .Y(n_1057) );
AOI22xp5_ASAP7_75t_L g1077 ( .A1(n_190), .A2(n_1078), .B1(n_1079), .B2(n_1098), .Y(n_1077) );
INVx1_ASAP7_75t_L g1100 ( .A(n_190), .Y(n_1100) );
AOI221xp5_ASAP7_75t_L g1028 ( .A1(n_191), .A2(n_201), .B1(n_931), .B2(n_1029), .C(n_1031), .Y(n_1028) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_192), .A2(n_200), .B1(n_399), .B2(n_689), .C(n_691), .Y(n_688) );
INVx1_ASAP7_75t_L g1426 ( .A(n_193), .Y(n_1426) );
INVx1_ASAP7_75t_L g768 ( .A(n_194), .Y(n_768) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_195), .A2(n_207), .B1(n_799), .B2(n_803), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_195), .A2(n_207), .B1(n_841), .B2(n_843), .Y(n_840) );
INVx1_ASAP7_75t_L g1336 ( .A(n_196), .Y(n_1336) );
INVx1_ASAP7_75t_L g255 ( .A(n_197), .Y(n_255) );
INVx1_ASAP7_75t_L g1399 ( .A(n_198), .Y(n_1399) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_199), .A2(n_245), .B1(n_417), .B2(n_675), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_202), .A2(n_239), .B1(n_545), .B2(n_1048), .Y(n_1047) );
INVxp67_ASAP7_75t_SL g708 ( .A(n_203), .Y(n_708) );
OAI221xp5_ASAP7_75t_L g734 ( .A1(n_203), .A2(n_205), .B1(n_333), .B2(n_348), .C(n_352), .Y(n_734) );
INVx1_ASAP7_75t_L g673 ( .A(n_204), .Y(n_673) );
OAI221xp5_ASAP7_75t_L g693 ( .A1(n_205), .A2(n_213), .B1(n_379), .B2(n_386), .C(n_411), .Y(n_693) );
INVx1_ASAP7_75t_L g267 ( .A(n_206), .Y(n_267) );
BUFx3_ASAP7_75t_L g365 ( .A(n_206), .Y(n_365) );
INVxp67_ASAP7_75t_SL g704 ( .A(n_209), .Y(n_704) );
CKINVDCx5p33_ASAP7_75t_R g466 ( .A(n_210), .Y(n_466) );
OAI211xp5_ASAP7_75t_L g572 ( .A1(n_211), .A2(n_573), .B(n_575), .C(n_589), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_213), .A2(n_216), .B1(n_725), .B2(n_728), .Y(n_724) );
INVxp67_ASAP7_75t_SL g710 ( .A(n_216), .Y(n_710) );
INVx1_ASAP7_75t_L g264 ( .A(n_218), .Y(n_264) );
INVx2_ASAP7_75t_L g357 ( .A(n_218), .Y(n_357) );
INVx1_ASAP7_75t_L g397 ( .A(n_218), .Y(n_397) );
XNOR2x1_ASAP7_75t_L g865 ( .A(n_219), .B(n_866), .Y(n_865) );
INVxp67_ASAP7_75t_SL g613 ( .A(n_220), .Y(n_613) );
CKINVDCx5p33_ASAP7_75t_R g567 ( .A(n_221), .Y(n_567) );
INVx1_ASAP7_75t_L g303 ( .A(n_224), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_224), .A2(n_247), .B1(n_372), .B2(n_409), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g1152 ( .A1(n_225), .A2(n_240), .B1(n_1123), .B2(n_1128), .Y(n_1152) );
INVxp67_ASAP7_75t_SL g972 ( .A(n_227), .Y(n_972) );
OAI211xp5_ASAP7_75t_SL g994 ( .A1(n_227), .A2(n_995), .B(n_996), .C(n_999), .Y(n_994) );
INVx1_ASAP7_75t_L g1217 ( .A(n_228), .Y(n_1217) );
INVx1_ASAP7_75t_L g1093 ( .A(n_230), .Y(n_1093) );
INVx1_ASAP7_75t_L g698 ( .A(n_231), .Y(n_698) );
AOI21xp5_ASAP7_75t_L g923 ( .A1(n_233), .A2(n_449), .B(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g1090 ( .A(n_235), .Y(n_1090) );
INVx1_ASAP7_75t_L g970 ( .A(n_236), .Y(n_970) );
AOI221xp5_ASAP7_75t_L g614 ( .A1(n_238), .A2(n_244), .B1(n_615), .B2(n_616), .C(n_618), .Y(n_614) );
INVx1_ASAP7_75t_L g911 ( .A(n_242), .Y(n_911) );
OAI211xp5_ASAP7_75t_L g626 ( .A1(n_245), .A2(n_573), .B(n_627), .C(n_634), .Y(n_626) );
INVx1_ASAP7_75t_L g320 ( .A(n_247), .Y(n_320) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_744), .B(n_1103), .C(n_1114), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g1103 ( .A1(n_250), .A2(n_744), .B(n_1104), .Y(n_1103) );
AO22x1_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_620), .B1(n_742), .B2(n_743), .Y(n_250) );
INVx1_ASAP7_75t_L g743 ( .A(n_251), .Y(n_743) );
XNOR2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_435), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
XNOR2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
NOR2x1_ASAP7_75t_L g256 ( .A(n_257), .B(n_358), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_279), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_260), .B1(n_273), .B2(n_274), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g338 ( .A1(n_259), .A2(n_339), .B1(n_341), .B2(n_342), .Y(n_338) );
INVx3_ASAP7_75t_L g712 ( .A(n_260), .Y(n_712) );
AND2x4_ASAP7_75t_L g260 ( .A(n_261), .B(n_265), .Y(n_260) );
AND2x4_ASAP7_75t_L g274 ( .A(n_261), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g379 ( .A(n_262), .B(n_380), .Y(n_379) );
INVxp67_ASAP7_75t_L g419 ( .A(n_262), .Y(n_419) );
OR2x2_ASAP7_75t_L g570 ( .A(n_262), .B(n_380), .Y(n_570) );
INVx1_ASAP7_75t_L g863 ( .A(n_262), .Y(n_863) );
BUFx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g403 ( .A(n_263), .Y(n_403) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g592 ( .A(n_265), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_265), .A2(n_595), .B1(n_635), .B2(n_636), .Y(n_634) );
BUFx6f_ASAP7_75t_L g890 ( .A(n_265), .Y(n_890) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_268), .Y(n_265) );
AND2x2_ASAP7_75t_L g275 ( .A(n_266), .B(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_266), .B(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g444 ( .A(n_266), .B(n_423), .Y(n_444) );
BUFx2_ASAP7_75t_L g472 ( .A(n_266), .Y(n_472) );
AND2x4_ASAP7_75t_L g574 ( .A(n_266), .B(n_374), .Y(n_574) );
AND2x4_ASAP7_75t_L g595 ( .A(n_266), .B(n_276), .Y(n_595) );
AND2x4_ASAP7_75t_SL g600 ( .A(n_266), .B(n_369), .Y(n_600) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_267), .Y(n_839) );
INVx3_ASAP7_75t_L g373 ( .A(n_268), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_268), .B(n_383), .Y(n_430) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_268), .Y(n_447) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
OR2x2_ASAP7_75t_L g407 ( .A(n_269), .B(n_272), .Y(n_407) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_269), .Y(n_468) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g277 ( .A(n_270), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g370 ( .A(n_270), .B(n_272), .Y(n_370) );
INVx2_ASAP7_75t_L g376 ( .A(n_270), .Y(n_376) );
INVx1_ASAP7_75t_L g382 ( .A(n_270), .Y(n_382) );
NAND2x1_ASAP7_75t_L g395 ( .A(n_270), .B(n_272), .Y(n_395) );
OR2x2_ASAP7_75t_L g461 ( .A(n_270), .B(n_272), .Y(n_461) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g278 ( .A(n_272), .Y(n_278) );
AND2x2_ASAP7_75t_L g375 ( .A(n_272), .B(n_376), .Y(n_375) );
BUFx2_ASAP7_75t_L g391 ( .A(n_272), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_272), .B(n_376), .Y(n_612) );
INVx2_ASAP7_75t_L g509 ( .A(n_274), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_274), .B(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g581 ( .A(n_276), .Y(n_581) );
INVx1_ASAP7_75t_L g631 ( .A(n_276), .Y(n_631) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g368 ( .A(n_277), .Y(n_368) );
BUFx3_ASAP7_75t_L g645 ( .A(n_277), .Y(n_645) );
AND2x4_ASAP7_75t_L g838 ( .A(n_277), .B(n_839), .Y(n_838) );
OAI31xp33_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_292), .A3(n_337), .B(n_356), .Y(n_279) );
OR2x6_ASAP7_75t_SL g281 ( .A(n_282), .B(n_286), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_283), .Y(n_347) );
AND2x4_ASAP7_75t_L g433 ( .A(n_283), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g508 ( .A(n_284), .B(n_403), .Y(n_508) );
INVx1_ASAP7_75t_L g727 ( .A(n_284), .Y(n_727) );
BUFx3_ASAP7_75t_L g314 ( .A(n_285), .Y(n_314) );
INVx3_ASAP7_75t_L g332 ( .A(n_285), .Y(n_332) );
NAND2xp33_ASAP7_75t_SL g653 ( .A(n_285), .B(n_315), .Y(n_653) );
INVx3_ASAP7_75t_L g506 ( .A(n_286), .Y(n_506) );
INVx1_ASAP7_75t_L g716 ( .A(n_286), .Y(n_716) );
BUFx2_ASAP7_75t_L g982 ( .A(n_286), .Y(n_982) );
BUFx2_ASAP7_75t_L g1407 ( .A(n_286), .Y(n_1407) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_287), .Y(n_311) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_287), .Y(n_486) );
BUFx8_ASAP7_75t_L g544 ( .A(n_287), .Y(n_544) );
AND2x4_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
INVxp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g296 ( .A(n_289), .Y(n_296) );
AND2x4_ASAP7_75t_L g328 ( .A(n_290), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g295 ( .A(n_291), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_291), .B(n_302), .Y(n_301) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_291), .Y(n_308) );
AND2x4_ASAP7_75t_L g344 ( .A(n_291), .B(n_345), .Y(n_344) );
OAI221xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_304), .B1(n_316), .B2(n_321), .C(n_333), .Y(n_292) );
OAI22xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_297), .B1(n_298), .B2(n_303), .Y(n_293) );
HB1xp67_ASAP7_75t_L g781 ( .A(n_294), .Y(n_781) );
INVx1_ASAP7_75t_L g795 ( .A(n_294), .Y(n_795) );
BUFx4f_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g558 ( .A(n_295), .Y(n_558) );
OR2x4_ASAP7_75t_L g801 ( .A(n_295), .B(n_802), .Y(n_801) );
OR2x4_ASAP7_75t_L g822 ( .A(n_295), .B(n_332), .Y(n_822) );
BUFx3_ASAP7_75t_L g1349 ( .A(n_295), .Y(n_1349) );
INVx1_ASAP7_75t_L g329 ( .A(n_296), .Y(n_329) );
INVx3_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx3_ASAP7_75t_L g319 ( .A(n_299), .Y(n_319) );
CKINVDCx8_ASAP7_75t_R g666 ( .A(n_299), .Y(n_666) );
INVx3_ASAP7_75t_L g796 ( .A(n_299), .Y(n_796) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g519 ( .A(n_300), .Y(n_519) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
BUFx2_ASAP7_75t_L g661 ( .A(n_301), .Y(n_661) );
INVx1_ASAP7_75t_L g307 ( .A(n_302), .Y(n_307) );
INVx2_ASAP7_75t_L g345 ( .A(n_302), .Y(n_345) );
OAI221xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_309), .B1(n_310), .B2(n_312), .C(n_313), .Y(n_304) );
OR2x6_ASAP7_75t_L g333 ( .A(n_305), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g1351 ( .A(n_305), .Y(n_1351) );
BUFx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_306), .Y(n_324) );
BUFx3_ASAP7_75t_L g790 ( .A(n_306), .Y(n_790) );
NAND2x1p5_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
BUFx2_ASAP7_75t_L g818 ( .A(n_307), .Y(n_818) );
INVx2_ASAP7_75t_L g351 ( .A(n_308), .Y(n_351) );
AND2x4_ASAP7_75t_L g434 ( .A(n_308), .B(n_355), .Y(n_434) );
BUFx2_ASAP7_75t_L g814 ( .A(n_308), .Y(n_814) );
OAI211xp5_ASAP7_75t_L g404 ( .A1(n_309), .A2(n_405), .B(n_408), .C(n_410), .Y(n_404) );
INVx2_ASAP7_75t_L g720 ( .A(n_310), .Y(n_720) );
INVx3_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_SL g317 ( .A(n_311), .Y(n_317) );
HB1xp67_ASAP7_75t_L g950 ( .A(n_311), .Y(n_950) );
INVx2_ASAP7_75t_SL g955 ( .A(n_311), .Y(n_955) );
INVx5_ASAP7_75t_L g1411 ( .A(n_311), .Y(n_1411) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
AND3x4_ASAP7_75t_L g480 ( .A(n_314), .B(n_315), .C(n_356), .Y(n_480) );
INVx3_ASAP7_75t_L g813 ( .A(n_314), .Y(n_813) );
INVx1_ASAP7_75t_L g336 ( .A(n_315), .Y(n_336) );
HB1xp67_ASAP7_75t_L g827 ( .A(n_315), .Y(n_827) );
OAI22xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_318), .B1(n_319), .B2(n_320), .Y(n_316) );
OAI22xp5_ASAP7_75t_L g785 ( .A1(n_319), .A2(n_752), .B1(n_767), .B2(n_786), .Y(n_785) );
OAI21xp5_ASAP7_75t_SL g321 ( .A1(n_322), .A2(n_325), .B(n_326), .Y(n_321) );
INVx3_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx3_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g513 ( .A(n_324), .B(n_508), .Y(n_513) );
BUFx6f_ASAP7_75t_L g784 ( .A(n_324), .Y(n_784) );
INVx4_ASAP7_75t_L g1357 ( .A(n_324), .Y(n_1357) );
BUFx2_ASAP7_75t_L g723 ( .A(n_327), .Y(n_723) );
BUFx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx8_ASAP7_75t_L g340 ( .A(n_328), .Y(n_340) );
NAND2x1p5_ASAP7_75t_L g418 ( .A(n_328), .B(n_335), .Y(n_418) );
BUFx3_ASAP7_75t_L g554 ( .A(n_328), .Y(n_554) );
AND2x2_ASAP7_75t_L g726 ( .A(n_328), .B(n_727), .Y(n_726) );
OR2x6_ASAP7_75t_L g492 ( .A(n_330), .B(n_363), .Y(n_492) );
OR2x2_ASAP7_75t_L g879 ( .A(n_330), .B(n_363), .Y(n_879) );
NAND2x1p5_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
NAND3x1_ASAP7_75t_L g549 ( .A(n_331), .B(n_332), .C(n_550), .Y(n_549) );
AND2x4_ASAP7_75t_L g335 ( .A(n_332), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g802 ( .A(n_332), .Y(n_802) );
OR2x6_ASAP7_75t_L g805 ( .A(n_332), .B(n_661), .Y(n_805) );
AND2x4_ASAP7_75t_L g808 ( .A(n_332), .B(n_344), .Y(n_808) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x6_ASAP7_75t_L g349 ( .A(n_335), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g353 ( .A(n_335), .B(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_L g495 ( .A(n_335), .B(n_429), .Y(n_495) );
AND2x4_ASAP7_75t_L g514 ( .A(n_339), .B(n_515), .Y(n_514) );
AND2x4_ASAP7_75t_L g677 ( .A(n_339), .B(n_515), .Y(n_677) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx8_ASAP7_75t_L g482 ( .A(n_340), .Y(n_482) );
INVx2_ASAP7_75t_L g878 ( .A(n_340), .Y(n_878) );
INVx3_ASAP7_75t_L g1073 ( .A(n_340), .Y(n_1073) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_341), .A2(n_378), .B1(n_384), .B2(n_385), .Y(n_377) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g669 ( .A(n_343), .Y(n_669) );
INVx1_ASAP7_75t_L g957 ( .A(n_343), .Y(n_957) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx2_ASAP7_75t_L g483 ( .A(n_344), .Y(n_483) );
BUFx2_ASAP7_75t_L g501 ( .A(n_344), .Y(n_501) );
BUFx3_ASAP7_75t_L g540 ( .A(n_344), .Y(n_540) );
AND2x2_ASAP7_75t_L g729 ( .A(n_344), .B(n_727), .Y(n_729) );
BUFx2_ASAP7_75t_L g877 ( .A(n_344), .Y(n_877) );
BUFx2_ASAP7_75t_L g948 ( .A(n_344), .Y(n_948) );
INVx1_ASAP7_75t_L g355 ( .A(n_345), .Y(n_355) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx4_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x4_ASAP7_75t_SL g494 ( .A(n_350), .B(n_495), .Y(n_494) );
NAND2x1_ASAP7_75t_L g535 ( .A(n_350), .B(n_495), .Y(n_535) );
AND2x2_ASAP7_75t_L g944 ( .A(n_350), .B(n_495), .Y(n_944) );
AND2x2_ASAP7_75t_L g1400 ( .A(n_350), .B(n_495), .Y(n_1400) );
INVx3_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g498 ( .A(n_354), .Y(n_498) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g475 ( .A(n_356), .Y(n_475) );
INVx2_ASAP7_75t_SL g619 ( .A(n_356), .Y(n_619) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx2_ASAP7_75t_L g363 ( .A(n_357), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_357), .B(n_383), .Y(n_388) );
NAND3xp33_ASAP7_75t_L g358 ( .A(n_359), .B(n_414), .C(n_425), .Y(n_358) );
NOR3xp33_ASAP7_75t_SL g359 ( .A(n_360), .B(n_392), .C(n_398), .Y(n_359) );
OAI21xp5_ASAP7_75t_SL g360 ( .A1(n_361), .A2(n_371), .B(n_377), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_362), .B(n_366), .Y(n_361) );
OAI221xp5_ASAP7_75t_L g697 ( .A1(n_362), .A2(n_690), .B1(n_692), .B2(n_698), .C(n_699), .Y(n_697) );
INVx2_ASAP7_75t_L g757 ( .A(n_362), .Y(n_757) );
INVx2_ASAP7_75t_L g1322 ( .A(n_362), .Y(n_1322) );
AND2x4_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx1_ASAP7_75t_L g432 ( .A(n_363), .Y(n_432) );
AND2x4_ASAP7_75t_L g401 ( .A(n_365), .B(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g451 ( .A(n_365), .Y(n_451) );
BUFx2_ASAP7_75t_L g848 ( .A(n_365), .Y(n_848) );
AND2x4_ASAP7_75t_L g859 ( .A(n_365), .B(n_381), .Y(n_859) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g454 ( .A(n_368), .Y(n_454) );
BUFx6f_ASAP7_75t_L g578 ( .A(n_369), .Y(n_578) );
AND2x6_ASAP7_75t_L g588 ( .A(n_369), .B(n_383), .Y(n_588) );
BUFx3_ASAP7_75t_L g615 ( .A(n_369), .Y(n_615) );
BUFx3_ASAP7_75t_L g629 ( .A(n_369), .Y(n_629) );
AND2x2_ASAP7_75t_L g851 ( .A(n_369), .B(n_852), .Y(n_851) );
BUFx3_ASAP7_75t_L g933 ( .A(n_369), .Y(n_933) );
INVx1_ASAP7_75t_L g1030 ( .A(n_369), .Y(n_1030) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g1380 ( .A(n_370), .Y(n_1380) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_SL g585 ( .A(n_373), .Y(n_585) );
INVx2_ASAP7_75t_L g633 ( .A(n_373), .Y(n_633) );
INVx1_ASAP7_75t_L g898 ( .A(n_373), .Y(n_898) );
BUFx2_ASAP7_75t_L g922 ( .A(n_374), .Y(n_922) );
INVx1_ASAP7_75t_L g1010 ( .A(n_374), .Y(n_1010) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx3_ASAP7_75t_L g409 ( .A(n_375), .Y(n_409) );
INVx2_ASAP7_75t_L g424 ( .A(n_375), .Y(n_424) );
BUFx3_ASAP7_75t_L g587 ( .A(n_375), .Y(n_587) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g471 ( .A(n_383), .Y(n_471) );
AND2x2_ASAP7_75t_L g900 ( .A(n_383), .B(n_465), .Y(n_900) );
INVx2_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
NAND2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_389), .Y(n_386) );
INVx1_ASAP7_75t_L g413 ( .A(n_387), .Y(n_413) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
BUFx2_ASAP7_75t_L g465 ( .A(n_391), .Y(n_465) );
INVx1_ASAP7_75t_L g603 ( .A(n_391), .Y(n_603) );
AND2x4_ASAP7_75t_L g855 ( .A(n_391), .B(n_848), .Y(n_855) );
AND2x2_ASAP7_75t_L g1382 ( .A(n_391), .B(n_848), .Y(n_1382) );
OR2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_396), .Y(n_393) );
INVx2_ASAP7_75t_SL g643 ( .A(n_394), .Y(n_643) );
OR2x2_ASAP7_75t_L g707 ( .A(n_394), .B(n_396), .Y(n_707) );
BUFx3_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_395), .Y(n_412) );
INVx1_ASAP7_75t_L g422 ( .A(n_396), .Y(n_422) );
INVx1_ASAP7_75t_L g429 ( .A(n_397), .Y(n_429) );
INVx1_ASAP7_75t_L g550 ( .A(n_397), .Y(n_550) );
OAI21xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_404), .B(n_411), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_SL g400 ( .A(n_401), .B(n_403), .Y(n_400) );
INVx4_ASAP7_75t_L g455 ( .A(n_401), .Y(n_455) );
INVx4_ASAP7_75t_L g583 ( .A(n_401), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_401), .B(n_772), .Y(n_771) );
INVx1_ASAP7_75t_SL g1031 ( .A(n_401), .Y(n_1031) );
AND2x4_ASAP7_75t_L g1344 ( .A(n_401), .B(n_772), .Y(n_1344) );
AND2x4_ASAP7_75t_L g450 ( .A(n_402), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g862 ( .A(n_402), .Y(n_862) );
OR2x2_ASAP7_75t_L g652 ( .A(n_403), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g773 ( .A(n_403), .Y(n_773) );
HB1xp67_ASAP7_75t_L g829 ( .A(n_403), .Y(n_829) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g1335 ( .A(n_406), .Y(n_1335) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
BUFx3_ASAP7_75t_L g690 ( .A(n_407), .Y(n_690) );
BUFx2_ASAP7_75t_L g753 ( .A(n_407), .Y(n_753) );
BUFx2_ASAP7_75t_L g1332 ( .A(n_407), .Y(n_1332) );
OR2x6_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
INVx4_ASAP7_75t_L g463 ( .A(n_412), .Y(n_463) );
BUFx4f_ASAP7_75t_L g474 ( .A(n_412), .Y(n_474) );
BUFx4f_ASAP7_75t_L g692 ( .A(n_412), .Y(n_692) );
BUFx6f_ASAP7_75t_L g756 ( .A(n_412), .Y(n_756) );
BUFx4f_ASAP7_75t_L g918 ( .A(n_412), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_420), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
OR2x6_ASAP7_75t_L g477 ( .A(n_418), .B(n_419), .Y(n_477) );
INVx2_ASAP7_75t_L g733 ( .A(n_418), .Y(n_733) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AOI222xp33_ASAP7_75t_L g700 ( .A1(n_421), .A2(n_701), .B1(n_704), .B2(n_705), .C1(n_706), .C2(n_708), .Y(n_700) );
AND2x4_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
INVx3_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g1033 ( .A(n_424), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_431), .Y(n_427) );
AND2x4_ASAP7_75t_L g566 ( .A(n_428), .B(n_518), .Y(n_566) );
OR2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_L g702 ( .A(n_429), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_430), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
BUFx2_ASAP7_75t_L g886 ( .A(n_432), .Y(n_886) );
INVx1_ASAP7_75t_L g1041 ( .A(n_432), .Y(n_1041) );
INVx3_ASAP7_75t_L g736 ( .A(n_433), .Y(n_736) );
BUFx12f_ASAP7_75t_L g487 ( .A(n_434), .Y(n_487) );
BUFx3_ASAP7_75t_L g545 ( .A(n_434), .Y(n_545) );
BUFx2_ASAP7_75t_L g717 ( .A(n_434), .Y(n_717) );
INVx5_ASAP7_75t_L g952 ( .A(n_434), .Y(n_952) );
BUFx3_ASAP7_75t_L g1408 ( .A(n_434), .Y(n_1408) );
XNOR2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_528), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NAND3xp33_ASAP7_75t_L g439 ( .A(n_440), .B(n_521), .C(n_525), .Y(n_439) );
INVx1_ASAP7_75t_L g522 ( .A(n_441), .Y(n_522) );
AOI21x1_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_475), .B(n_476), .Y(n_441) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AOI221xp5_ASAP7_75t_L g892 ( .A1(n_444), .A2(n_588), .B1(n_869), .B2(n_893), .C(n_894), .Y(n_892) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_448), .B1(n_452), .B2(n_453), .Y(n_445) );
INVx3_ASAP7_75t_L g921 ( .A(n_447), .Y(n_921) );
BUFx6f_ASAP7_75t_L g1008 ( .A(n_447), .Y(n_1008) );
INVx3_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g618 ( .A(n_450), .Y(n_618) );
INVx1_ASAP7_75t_L g646 ( .A(n_450), .Y(n_646) );
INVx2_ASAP7_75t_L g1436 ( .A(n_450), .Y(n_1436) );
INVxp67_ASAP7_75t_L g836 ( .A(n_451), .Y(n_836) );
INVx1_ASAP7_75t_L g852 ( .A(n_451), .Y(n_852) );
INVx2_ASAP7_75t_L g617 ( .A(n_454), .Y(n_617) );
INVx1_ASAP7_75t_L g932 ( .A(n_454), .Y(n_932) );
HB1xp67_ASAP7_75t_L g1435 ( .A(n_454), .Y(n_1435) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_470), .B1(n_472), .B2(n_473), .Y(n_456) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
BUFx6f_ASAP7_75t_L g606 ( .A(n_459), .Y(n_606) );
BUFx4f_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx3_ASAP7_75t_L g687 ( .A(n_460), .Y(n_687) );
INVx2_ASAP7_75t_L g835 ( .A(n_460), .Y(n_835) );
INVx3_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OAI211xp5_ASAP7_75t_L g1092 ( .A1(n_462), .A2(n_1093), .B(n_1094), .C(n_1097), .Y(n_1092) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g1376 ( .A(n_463), .Y(n_1376) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_466), .B1(n_467), .B2(n_469), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g493 ( .A1(n_466), .A2(n_494), .B1(n_496), .B2(n_499), .C(n_500), .Y(n_493) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AOI222xp33_ASAP7_75t_L g511 ( .A1(n_469), .A2(n_512), .B1(n_514), .B2(n_516), .C1(n_517), .C2(n_520), .Y(n_511) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NOR2x1_ASAP7_75t_L g602 ( .A(n_471), .B(n_603), .Y(n_602) );
BUFx2_ASAP7_75t_L g648 ( .A(n_475), .Y(n_648) );
BUFx2_ASAP7_75t_L g737 ( .A(n_475), .Y(n_737) );
INVx3_ASAP7_75t_L g868 ( .A(n_477), .Y(n_868) );
INVx5_ASAP7_75t_L g973 ( .A(n_477), .Y(n_973) );
INVx1_ASAP7_75t_L g523 ( .A(n_478), .Y(n_523) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_493), .Y(n_478) );
AOI33xp33_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .A3(n_484), .B1(n_488), .B2(n_490), .B3(n_491), .Y(n_479) );
AOI33xp33_ASAP7_75t_L g538 ( .A1(n_480), .A2(n_539), .A3(n_541), .B1(n_546), .B2(n_547), .B3(n_551), .Y(n_538) );
INVx1_ASAP7_75t_L g882 ( .A(n_480), .Y(n_882) );
AOI33xp33_ASAP7_75t_L g946 ( .A1(n_480), .A2(n_547), .A3(n_947), .B1(n_949), .B2(n_953), .B3(n_956), .Y(n_946) );
BUFx3_ASAP7_75t_L g979 ( .A(n_480), .Y(n_979) );
AOI33xp33_ASAP7_75t_L g1045 ( .A1(n_480), .A2(n_792), .A3(n_1046), .B1(n_1047), .B2(n_1049), .B3(n_1050), .Y(n_1045) );
AOI33xp33_ASAP7_75t_L g1066 ( .A1(n_480), .A2(n_1067), .A3(n_1070), .B1(n_1071), .B2(n_1072), .B3(n_1074), .Y(n_1066) );
BUFx2_ASAP7_75t_L g976 ( .A(n_482), .Y(n_976) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_486), .Y(n_489) );
INVx2_ASAP7_75t_L g786 ( .A(n_486), .Y(n_786) );
AND2x4_ASAP7_75t_L g824 ( .A(n_486), .B(n_802), .Y(n_824) );
INVx1_ASAP7_75t_L g788 ( .A(n_489), .Y(n_788) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g872 ( .A1(n_494), .A2(n_496), .B1(n_873), .B2(n_874), .Y(n_872) );
AND2x4_ASAP7_75t_SL g496 ( .A(n_495), .B(n_497), .Y(n_496) );
AND2x4_ASAP7_75t_L g500 ( .A(n_495), .B(n_501), .Y(n_500) );
AND2x4_ASAP7_75t_L g537 ( .A(n_495), .B(n_497), .Y(n_537) );
INVx1_ASAP7_75t_L g671 ( .A(n_496), .Y(n_671) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx3_ASAP7_75t_L g563 ( .A(n_500), .Y(n_563) );
NOR3xp33_ASAP7_75t_L g649 ( .A(n_500), .B(n_650), .C(n_670), .Y(n_649) );
INVx3_ASAP7_75t_L g962 ( .A(n_500), .Y(n_962) );
HB1xp67_ASAP7_75t_L g1414 ( .A(n_500), .Y(n_1414) );
BUFx2_ASAP7_75t_L g1404 ( .A(n_501), .Y(n_1404) );
INVx1_ASAP7_75t_L g527 ( .A(n_502), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_510), .Y(n_502) );
NAND2x1_ASAP7_75t_L g503 ( .A(n_504), .B(n_509), .Y(n_503) );
INVx2_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_505), .A2(n_514), .B1(n_889), .B2(n_891), .Y(n_902) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
INVx2_ASAP7_75t_L g1353 ( .A(n_506), .Y(n_1353) );
INVxp67_ASAP7_75t_L g559 ( .A(n_507), .Y(n_559) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g515 ( .A(n_508), .Y(n_515) );
OR2x2_ASAP7_75t_L g518 ( .A(n_508), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g526 ( .A(n_511), .Y(n_526) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x4_ASAP7_75t_L g569 ( .A(n_513), .B(n_570), .Y(n_569) );
AND2x4_ASAP7_75t_L g675 ( .A(n_513), .B(n_570), .Y(n_675) );
AND2x4_ASAP7_75t_L g561 ( .A(n_515), .B(n_544), .Y(n_561) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B(n_524), .Y(n_521) );
OAI21xp33_ASAP7_75t_L g525 ( .A1(n_524), .A2(n_526), .B(n_527), .Y(n_525) );
NAND3xp33_ASAP7_75t_L g529 ( .A(n_530), .B(n_564), .C(n_571), .Y(n_529) );
NOR3xp33_ASAP7_75t_L g530 ( .A(n_531), .B(n_555), .C(n_562), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_538), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_534), .B1(n_536), .B2(n_537), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g1061 ( .A1(n_534), .A2(n_537), .B1(n_1062), .B2(n_1063), .Y(n_1061) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_537), .A2(n_943), .B1(n_944), .B2(n_945), .Y(n_942) );
AOI22xp5_ASAP7_75t_L g968 ( .A1(n_537), .A2(n_944), .B1(n_969), .B2(n_970), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_537), .A2(n_944), .B1(n_1052), .B2(n_1053), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g1398 ( .A1(n_537), .A2(n_1399), .B1(n_1400), .B2(n_1401), .Y(n_1398) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx3_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_SL g655 ( .A(n_544), .Y(n_655) );
INVx3_ASAP7_75t_L g986 ( .A(n_544), .Y(n_986) );
AOI33xp33_ASAP7_75t_L g1402 ( .A1(n_547), .A2(n_979), .A3(n_1403), .B1(n_1405), .B2(n_1409), .B3(n_1412), .Y(n_1402) );
BUFx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
BUFx2_ASAP7_75t_L g792 ( .A(n_548), .Y(n_792) );
BUFx2_ASAP7_75t_L g1074 ( .A(n_548), .Y(n_1074) );
INVx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx3_ASAP7_75t_L g664 ( .A(n_549), .Y(n_664) );
OAI33xp33_ASAP7_75t_L g1345 ( .A1(n_549), .A2(n_651), .A3(n_1346), .B1(n_1352), .B2(n_1354), .B3(n_1355), .Y(n_1345) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_SL g1069 ( .A(n_554), .Y(n_1069) );
OR2x6_ASAP7_75t_L g556 ( .A(n_557), .B(n_559), .Y(n_556) );
OR2x2_ASAP7_75t_L g959 ( .A(n_557), .B(n_559), .Y(n_959) );
INVx2_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_561), .A2(n_635), .B1(n_636), .B2(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g960 ( .A(n_561), .Y(n_960) );
INVx2_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
NAND3xp33_ASAP7_75t_SL g871 ( .A(n_563), .B(n_872), .C(n_875), .Y(n_871) );
AND4x1_ASAP7_75t_L g1042 ( .A(n_563), .B(n_1043), .C(n_1045), .D(n_1051), .Y(n_1042) );
AOI21xp33_ASAP7_75t_SL g564 ( .A1(n_565), .A2(n_567), .B(n_568), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g672 ( .A1(n_565), .A2(n_673), .B(n_674), .Y(n_672) );
AOI221xp5_ASAP7_75t_L g867 ( .A1(n_565), .A2(n_868), .B1(n_869), .B2(n_870), .C(n_871), .Y(n_867) );
AOI21xp33_ASAP7_75t_SL g937 ( .A1(n_565), .A2(n_938), .B(n_939), .Y(n_937) );
AOI211x1_ASAP7_75t_L g965 ( .A1(n_565), .A2(n_966), .B(n_967), .C(n_988), .Y(n_965) );
AOI21xp33_ASAP7_75t_L g1019 ( .A1(n_565), .A2(n_1020), .B(n_1021), .Y(n_1019) );
NAND2xp33_ASAP7_75t_L g1075 ( .A(n_565), .B(n_1076), .Y(n_1075) );
AOI21xp5_ASAP7_75t_L g1415 ( .A1(n_565), .A2(n_1416), .B(n_1417), .Y(n_1415) );
INVx8_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g990 ( .A(n_569), .Y(n_990) );
OAI21xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_596), .B(n_619), .Y(n_571) );
INVx2_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_574), .A2(n_890), .B1(n_913), .B2(n_914), .Y(n_912) );
INVx3_ASAP7_75t_L g995 ( .A(n_574), .Y(n_995) );
AOI21xp5_ASAP7_75t_SL g575 ( .A1(n_576), .A2(n_584), .B(n_588), .Y(n_575) );
BUFx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g1423 ( .A(n_580), .Y(n_1423) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
HB1xp67_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
BUFx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_588), .A2(n_628), .B(n_632), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g910 ( .A1(n_588), .A2(n_594), .B(n_911), .Y(n_910) );
AOI21xp5_ASAP7_75t_L g996 ( .A1(n_588), .A2(n_997), .B(n_998), .Y(n_996) );
AOI21xp5_ASAP7_75t_L g1027 ( .A1(n_588), .A2(n_1028), .B(n_1032), .Y(n_1027) );
AOI21xp5_ASAP7_75t_L g1085 ( .A1(n_588), .A2(n_1086), .B(n_1087), .Y(n_1085) );
AOI21xp5_ASAP7_75t_L g1420 ( .A1(n_588), .A2(n_1421), .B(n_1424), .Y(n_1420) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B1(n_593), .B2(n_594), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g1425 ( .A1(n_591), .A2(n_1426), .B1(n_1427), .B2(n_1428), .Y(n_1425) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_594), .A2(n_890), .B1(n_1000), .B2(n_1001), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_594), .A2(n_890), .B1(n_1025), .B2(n_1026), .Y(n_1024) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g888 ( .A1(n_595), .A2(n_889), .B1(n_890), .B2(n_891), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_595), .A2(n_890), .B1(n_1089), .B2(n_1090), .Y(n_1088) );
INVx1_ASAP7_75t_L g1429 ( .A(n_595), .Y(n_1429) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g638 ( .A(n_598), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g1438 ( .A1(n_598), .A2(n_602), .B1(n_1399), .B2(n_1401), .Y(n_1438) );
INVx4_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
BUFx3_ASAP7_75t_L g896 ( .A(n_600), .Y(n_896) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g639 ( .A(n_602), .Y(n_639) );
OAI221xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_607), .B1(n_608), .B2(n_613), .C(n_614), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g684 ( .A(n_608), .Y(n_684) );
BUFx2_ASAP7_75t_L g1037 ( .A(n_608), .Y(n_1037) );
BUFx6f_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx4_ASAP7_75t_L g765 ( .A(n_610), .Y(n_765) );
INVx2_ASAP7_75t_SL g928 ( .A(n_610), .Y(n_928) );
BUFx6f_ASAP7_75t_L g1342 ( .A(n_610), .Y(n_1342) );
INVx8_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
BUFx2_ASAP7_75t_L g696 ( .A(n_611), .Y(n_696) );
OR2x2_ASAP7_75t_L g847 ( .A(n_611), .B(n_848), .Y(n_847) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g924 ( .A(n_617), .Y(n_924) );
INVx1_ASAP7_75t_L g742 ( .A(n_620), .Y(n_742) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_622), .B1(n_678), .B2(n_741), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND4x1_ASAP7_75t_L g624 ( .A(n_625), .B(n_649), .C(n_672), .D(n_676), .Y(n_624) );
OAI21xp5_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_637), .B(n_648), .Y(n_625) );
INVx2_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
BUFx2_ASAP7_75t_L g1003 ( .A(n_639), .Y(n_1003) );
OAI211xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B(n_644), .C(n_647), .Y(n_640) );
OAI221xp5_ASAP7_75t_L g665 ( .A1(n_641), .A2(n_655), .B1(n_666), .B2(n_667), .C(n_668), .Y(n_665) );
OAI211xp5_ASAP7_75t_L g1004 ( .A1(n_642), .A2(n_1005), .B(n_1006), .C(n_1007), .Y(n_1004) );
OAI22xp5_ASAP7_75t_L g1334 ( .A1(n_642), .A2(n_1335), .B1(n_1336), .B2(n_1337), .Y(n_1334) );
INVx5_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g1096 ( .A(n_645), .Y(n_1096) );
OAI22xp5_ASAP7_75t_SL g650 ( .A1(n_651), .A2(n_654), .B1(n_663), .B2(n_665), .Y(n_650) );
BUFx8_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
BUFx4f_ASAP7_75t_L g779 ( .A(n_652), .Y(n_779) );
BUFx2_ASAP7_75t_L g721 ( .A(n_653), .Y(n_721) );
OAI221xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_656), .B1(n_657), .B2(n_658), .C(n_662), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g1354 ( .A1(n_658), .A2(n_788), .B1(n_1333), .B2(n_1340), .Y(n_1354) );
INVx3_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
BUFx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
CKINVDCx5p33_ASAP7_75t_R g663 ( .A(n_664), .Y(n_663) );
AOI33xp33_ASAP7_75t_L g974 ( .A1(n_664), .A2(n_975), .A3(n_979), .B1(n_980), .B2(n_984), .B3(n_987), .Y(n_974) );
OAI22xp5_ASAP7_75t_L g1352 ( .A1(n_666), .A2(n_1329), .B1(n_1339), .B2(n_1353), .Y(n_1352) );
INVx1_ASAP7_75t_L g741 ( .A(n_678), .Y(n_741) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
XNOR2x1_ASAP7_75t_L g679 ( .A(n_680), .B(n_740), .Y(n_679) );
OR2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_713), .Y(n_680) );
NAND3xp33_ASAP7_75t_SL g681 ( .A(n_682), .B(n_700), .C(n_709), .Y(n_681) );
AOI211xp5_ASAP7_75t_SL g682 ( .A1(n_683), .A2(n_688), .B(n_693), .C(n_694), .Y(n_682) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OAI221xp5_ASAP7_75t_L g925 ( .A1(n_686), .A2(n_926), .B1(n_927), .B2(n_929), .C(n_930), .Y(n_925) );
BUFx6f_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx2_ASAP7_75t_SL g761 ( .A(n_687), .Y(n_761) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVxp67_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AND2x4_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
AOI211xp5_ASAP7_75t_L g730 ( .A1(n_705), .A2(n_731), .B(n_734), .C(n_735), .Y(n_730) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
A2O1A1Ixp33_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_730), .B(n_737), .C(n_738), .Y(n_713) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_718), .B1(n_719), .B2(n_722), .C(n_724), .Y(n_714) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g936 ( .A(n_737), .Y(n_936) );
INVx1_ASAP7_75t_L g1440 ( .A(n_737), .Y(n_1440) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_1013), .B1(n_1014), .B2(n_1102), .Y(n_744) );
INVx1_ASAP7_75t_L g1102 ( .A(n_745), .Y(n_1102) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_904), .B1(n_905), .B2(n_1012), .Y(n_745) );
INVx1_ASAP7_75t_L g1012 ( .A(n_746), .Y(n_1012) );
AO22x1_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_864), .B1(n_865), .B2(n_903), .Y(n_746) );
INVx1_ASAP7_75t_L g903 ( .A(n_747), .Y(n_903) );
NAND3xp33_ASAP7_75t_L g748 ( .A(n_749), .B(n_797), .C(n_830), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_750), .B(n_777), .Y(n_749) );
OAI33xp33_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_757), .A3(n_758), .B1(n_766), .B2(n_769), .B3(n_774), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_753), .B1(n_754), .B2(n_755), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g774 ( .A1(n_753), .A2(n_763), .B1(n_775), .B2(n_776), .Y(n_774) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_754), .A2(n_768), .B1(n_788), .B2(n_789), .Y(n_787) );
HB1xp67_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
OAI22xp33_ASAP7_75t_L g766 ( .A1(n_756), .A2(n_760), .B1(n_767), .B2(n_768), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_760), .B1(n_762), .B2(n_763), .Y(n_758) );
OAI22xp33_ASAP7_75t_L g780 ( .A1(n_759), .A2(n_775), .B1(n_781), .B2(n_782), .Y(n_780) );
OAI221xp5_ASAP7_75t_L g1035 ( .A1(n_760), .A2(n_1036), .B1(n_1037), .B2(n_1038), .C(n_1039), .Y(n_1035) );
OAI22xp5_ASAP7_75t_L g1338 ( .A1(n_760), .A2(n_1339), .B1(n_1340), .B2(n_1341), .Y(n_1338) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_762), .A2(n_776), .B1(n_794), .B2(n_796), .Y(n_793) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
OAI33xp33_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_780), .A3(n_785), .B1(n_787), .B2(n_791), .B3(n_793), .Y(n_777) );
BUFx3_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx2_ASAP7_75t_SL g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g1048 ( .A(n_786), .Y(n_1048) );
BUFx6f_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
OAI31xp33_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_806), .A3(n_819), .B(n_825), .Y(n_797) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx2_ASAP7_75t_SL g800 ( .A(n_801), .Y(n_800) );
BUFx3_ASAP7_75t_L g1368 ( .A(n_801), .Y(n_1368) );
INVx2_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g1370 ( .A(n_805), .Y(n_1370) );
CKINVDCx8_ASAP7_75t_R g807 ( .A(n_808), .Y(n_807) );
CKINVDCx8_ASAP7_75t_R g1362 ( .A(n_808), .Y(n_1362) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_811), .B1(n_815), .B2(n_816), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_810), .A2(n_854), .B1(n_856), .B2(n_857), .Y(n_853) );
BUFx3_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
AND2x2_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .Y(n_812) );
AND2x4_ASAP7_75t_L g817 ( .A(n_813), .B(n_818), .Y(n_817) );
AND2x4_ASAP7_75t_L g1364 ( .A(n_813), .B(n_814), .Y(n_1364) );
BUFx6f_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g1363 ( .A1(n_817), .A2(n_1364), .B1(n_1365), .B2(n_1366), .Y(n_1363) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx2_ASAP7_75t_L g1360 ( .A(n_824), .Y(n_1360) );
AND2x2_ASAP7_75t_SL g825 ( .A(n_826), .B(n_828), .Y(n_825) );
AND2x2_ASAP7_75t_L g1371 ( .A(n_826), .B(n_828), .Y(n_1371) );
INVx1_ASAP7_75t_SL g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
OAI31xp33_ASAP7_75t_SL g830 ( .A1(n_831), .A2(n_840), .A3(n_849), .B(n_860), .Y(n_830) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g1112 ( .A(n_833), .B(n_1113), .Y(n_1112) );
AND2x4_ASAP7_75t_SL g1315 ( .A(n_833), .B(n_1316), .Y(n_1315) );
INVx3_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
OR2x6_ASAP7_75t_L g834 ( .A(n_835), .B(n_836), .Y(n_834) );
OR2x6_ASAP7_75t_L g842 ( .A(n_835), .B(n_839), .Y(n_842) );
INVxp67_ASAP7_75t_L g1326 ( .A(n_835), .Y(n_1326) );
INVx3_ASAP7_75t_SL g837 ( .A(n_838), .Y(n_837) );
INVx4_ASAP7_75t_L g1374 ( .A(n_838), .Y(n_1374) );
HB1xp67_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
BUFx6f_ASAP7_75t_L g1385 ( .A(n_842), .Y(n_1385) );
INVx2_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx2_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx2_ASAP7_75t_L g1387 ( .A(n_847), .Y(n_1387) );
INVx3_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
AND2x2_ASAP7_75t_L g1378 ( .A(n_852), .B(n_1379), .Y(n_1378) );
BUFx3_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g1381 ( .A1(n_857), .A2(n_1365), .B1(n_1382), .B2(n_1383), .Y(n_1381) );
INVx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
OAI31xp33_ASAP7_75t_L g1372 ( .A1(n_860), .A2(n_1373), .A3(n_1375), .B(n_1384), .Y(n_1372) );
BUFx3_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
AND2x4_ASAP7_75t_L g861 ( .A(n_862), .B(n_863), .Y(n_861) );
INVx1_ASAP7_75t_L g1113 ( .A(n_862), .Y(n_1113) );
NOR2xp33_ASAP7_75t_L g1316 ( .A(n_862), .B(n_1105), .Y(n_1316) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
AND2x2_ASAP7_75t_L g866 ( .A(n_867), .B(n_884), .Y(n_866) );
AOI222xp33_ASAP7_75t_L g895 ( .A1(n_873), .A2(n_874), .B1(n_896), .B2(n_897), .C1(n_899), .C2(n_900), .Y(n_895) );
AOI22xp5_ASAP7_75t_L g875 ( .A1(n_876), .A2(n_880), .B1(n_881), .B2(n_883), .Y(n_875) );
INVx1_ASAP7_75t_L g978 ( .A(n_877), .Y(n_978) );
AOI21xp5_ASAP7_75t_L g884 ( .A1(n_885), .A2(n_887), .B(n_901), .Y(n_884) );
OAI21xp5_ASAP7_75t_L g1083 ( .A1(n_885), .A2(n_1084), .B(n_1091), .Y(n_1083) );
INVx2_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx1_ASAP7_75t_L g1011 ( .A(n_886), .Y(n_1011) );
NAND3xp33_ASAP7_75t_L g887 ( .A(n_888), .B(n_892), .C(n_895), .Y(n_887) );
INVx2_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
XNOR2x2_ASAP7_75t_L g905 ( .A(n_906), .B(n_963), .Y(n_905) );
NAND3xp33_ASAP7_75t_L g907 ( .A(n_908), .B(n_937), .C(n_940), .Y(n_907) );
OAI31xp33_ASAP7_75t_L g908 ( .A1(n_909), .A2(n_915), .A3(n_934), .B(n_935), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_910), .B(n_912), .Y(n_909) );
OAI211xp5_ASAP7_75t_L g916 ( .A1(n_917), .A2(n_918), .B(n_919), .C(n_923), .Y(n_916) );
OAI22xp5_ASAP7_75t_L g1328 ( .A1(n_918), .A2(n_1329), .B1(n_1330), .B2(n_1333), .Y(n_1328) );
INVx2_ASAP7_75t_SL g920 ( .A(n_921), .Y(n_920) );
HB1xp67_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
OAI22xp33_ASAP7_75t_L g1323 ( .A1(n_928), .A2(n_1324), .B1(n_1325), .B2(n_1327), .Y(n_1323) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
NOR3xp33_ASAP7_75t_L g940 ( .A(n_941), .B(n_958), .C(n_961), .Y(n_940) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_942), .B(n_946), .Y(n_941) );
INVx2_ASAP7_75t_R g951 ( .A(n_952), .Y(n_951) );
INVx1_ASAP7_75t_L g983 ( .A(n_952), .Y(n_983) );
INVx2_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
INVx1_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
NAND4xp25_ASAP7_75t_SL g967 ( .A(n_962), .B(n_968), .C(n_971), .D(n_974), .Y(n_967) );
NAND4xp25_ASAP7_75t_SL g1060 ( .A(n_962), .B(n_1061), .C(n_1064), .D(n_1066), .Y(n_1060) );
XNOR2x2_ASAP7_75t_L g963 ( .A(n_964), .B(n_965), .Y(n_963) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_972), .B(n_973), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g1064 ( .A(n_973), .B(n_1065), .Y(n_1064) );
INVx1_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
INVx1_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
INVx1_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g988 ( .A(n_989), .B(n_993), .Y(n_988) );
AOI21xp5_ASAP7_75t_L g989 ( .A1(n_990), .A2(n_991), .B(n_992), .Y(n_989) );
AOI21xp5_ASAP7_75t_L g1080 ( .A1(n_990), .A2(n_1081), .B(n_1082), .Y(n_1080) );
OAI21xp33_ASAP7_75t_L g993 ( .A1(n_994), .A2(n_1002), .B(n_1011), .Y(n_993) );
INVx1_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
INVx2_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
OAI22x1_ASAP7_75t_L g1015 ( .A1(n_1016), .A2(n_1055), .B1(n_1056), .B2(n_1101), .Y(n_1015) );
INVx2_ASAP7_75t_L g1101 ( .A(n_1016), .Y(n_1101) );
AO21x2_ASAP7_75t_L g1016 ( .A1(n_1017), .A2(n_1018), .B(n_1054), .Y(n_1016) );
NAND3xp33_ASAP7_75t_SL g1018 ( .A(n_1019), .B(n_1022), .C(n_1042), .Y(n_1018) );
OAI21xp5_ASAP7_75t_L g1022 ( .A1(n_1023), .A2(n_1034), .B(n_1041), .Y(n_1022) );
INVx1_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
INVx1_ASAP7_75t_L g1040 ( .A(n_1030), .Y(n_1040) );
INVx1_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
INVx2_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
NAND2x1p5_ASAP7_75t_L g1056 ( .A(n_1057), .B(n_1077), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g1058 ( .A(n_1059), .B(n_1075), .Y(n_1058) );
INVxp67_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
NOR2xp33_ASAP7_75t_SL g1098 ( .A(n_1060), .B(n_1099), .Y(n_1098) );
INVx2_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g1099 ( .A(n_1075), .B(n_1100), .Y(n_1099) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
NAND2xp5_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1083), .Y(n_1079) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
OR2x2_ASAP7_75t_L g1104 ( .A(n_1105), .B(n_1111), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
NOR2xp33_ASAP7_75t_L g1106 ( .A(n_1107), .B(n_1109), .Y(n_1106) );
NOR2xp33_ASAP7_75t_L g1391 ( .A(n_1107), .B(n_1110), .Y(n_1391) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1107), .Y(n_1442) );
HB1xp67_ASAP7_75t_L g1107 ( .A(n_1108), .Y(n_1107) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
NOR2xp33_ASAP7_75t_L g1444 ( .A(n_1110), .B(n_1442), .Y(n_1444) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
OAI221xp5_ASAP7_75t_L g1114 ( .A1(n_1115), .A2(n_1309), .B1(n_1311), .B2(n_1317), .C(n_1388), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_1116), .B(n_1251), .Y(n_1115) );
OAI32xp33_ASAP7_75t_L g1116 ( .A1(n_1117), .A2(n_1180), .A3(n_1212), .B1(n_1226), .B2(n_1241), .Y(n_1116) );
OAI311xp33_ASAP7_75t_L g1117 ( .A1(n_1118), .A2(n_1145), .A3(n_1150), .B1(n_1154), .C1(n_1173), .Y(n_1117) );
NAND2xp5_ASAP7_75t_L g1118 ( .A(n_1119), .B(n_1135), .Y(n_1118) );
OR2x2_ASAP7_75t_L g1235 ( .A(n_1119), .B(n_1236), .Y(n_1235) );
CKINVDCx5p33_ASAP7_75t_R g1119 ( .A(n_1120), .Y(n_1119) );
NOR2xp33_ASAP7_75t_L g1186 ( .A(n_1120), .B(n_1187), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1120), .B(n_1172), .Y(n_1201) );
OR2x2_ASAP7_75t_L g1231 ( .A(n_1120), .B(n_1207), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1263 ( .A(n_1120), .B(n_1189), .Y(n_1263) );
NOR2xp33_ASAP7_75t_L g1292 ( .A(n_1120), .B(n_1203), .Y(n_1292) );
INVx4_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
NOR2xp33_ASAP7_75t_L g1157 ( .A(n_1121), .B(n_1158), .Y(n_1157) );
INVx4_ASAP7_75t_L g1177 ( .A(n_1121), .Y(n_1177) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1121), .Y(n_1206) );
NAND2xp5_ASAP7_75t_L g1223 ( .A(n_1121), .B(n_1191), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1121), .B(n_1183), .Y(n_1237) );
OR2x2_ASAP7_75t_L g1244 ( .A(n_1121), .B(n_1179), .Y(n_1244) );
OAI22xp5_ASAP7_75t_L g1245 ( .A1(n_1121), .A2(n_1177), .B1(n_1246), .B2(n_1247), .Y(n_1245) );
NOR2xp33_ASAP7_75t_L g1268 ( .A(n_1121), .B(n_1184), .Y(n_1268) );
NAND2xp5_ASAP7_75t_SL g1277 ( .A(n_1121), .B(n_1179), .Y(n_1277) );
AND2x4_ASAP7_75t_SL g1121 ( .A(n_1122), .B(n_1130), .Y(n_1121) );
AND2x4_ASAP7_75t_L g1123 ( .A(n_1124), .B(n_1125), .Y(n_1123) );
AND2x6_ASAP7_75t_L g1128 ( .A(n_1124), .B(n_1129), .Y(n_1128) );
AND2x6_ASAP7_75t_L g1131 ( .A(n_1124), .B(n_1132), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_1124), .B(n_1134), .Y(n_1133) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1124), .B(n_1134), .Y(n_1139) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1124), .B(n_1134), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1216 ( .A(n_1124), .B(n_1125), .Y(n_1216) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_1126), .B(n_1127), .Y(n_1125) );
INVx2_ASAP7_75t_L g1218 ( .A(n_1128), .Y(n_1218) );
OAI21xp5_ASAP7_75t_L g1441 ( .A1(n_1134), .A2(n_1442), .B(n_1443), .Y(n_1441) );
AOI222xp33_ASAP7_75t_L g1232 ( .A1(n_1135), .A2(n_1233), .B1(n_1234), .B2(n_1237), .C1(n_1238), .C2(n_1239), .Y(n_1232) );
O2A1O1Ixp33_ASAP7_75t_SL g1271 ( .A1(n_1135), .A2(n_1268), .B(n_1272), .C(n_1278), .Y(n_1271) );
O2A1O1Ixp33_ASAP7_75t_L g1293 ( .A1(n_1135), .A2(n_1294), .B(n_1295), .C(n_1296), .Y(n_1293) );
CKINVDCx5p33_ASAP7_75t_R g1135 ( .A(n_1136), .Y(n_1135) );
OR2x2_ASAP7_75t_L g1228 ( .A(n_1136), .B(n_1171), .Y(n_1228) );
OR2x2_ASAP7_75t_L g1136 ( .A(n_1137), .B(n_1141), .Y(n_1136) );
INVx2_ASAP7_75t_L g1185 ( .A(n_1137), .Y(n_1185) );
NAND2xp5_ASAP7_75t_L g1137 ( .A(n_1138), .B(n_1140), .Y(n_1137) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1141), .Y(n_1172) );
OR2x2_ASAP7_75t_L g1197 ( .A(n_1141), .B(n_1185), .Y(n_1197) );
NOR2xp33_ASAP7_75t_L g1298 ( .A(n_1141), .B(n_1299), .Y(n_1298) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
OR2x2_ASAP7_75t_L g1184 ( .A(n_1142), .B(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1142), .Y(n_1192) );
NAND2xp5_ASAP7_75t_L g1142 ( .A(n_1143), .B(n_1144), .Y(n_1142) );
NAND2xp5_ASAP7_75t_L g1200 ( .A(n_1145), .B(n_1201), .Y(n_1200) );
OAI211xp5_ASAP7_75t_L g1252 ( .A1(n_1145), .A2(n_1253), .B(n_1261), .C(n_1271), .Y(n_1252) );
OR2x2_ASAP7_75t_L g1289 ( .A(n_1145), .B(n_1184), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1145), .B(n_1259), .Y(n_1303) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1146), .Y(n_1145) );
INVx3_ASAP7_75t_L g1171 ( .A(n_1146), .Y(n_1171) );
OR2x2_ASAP7_75t_L g1240 ( .A(n_1146), .B(n_1185), .Y(n_1240) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1146), .B(n_1233), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1146), .B(n_1185), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_1147), .B(n_1148), .Y(n_1146) );
HB1xp67_ASAP7_75t_L g1310 ( .A(n_1149), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1150), .B(n_1159), .Y(n_1183) );
NOR2xp33_ASAP7_75t_L g1189 ( .A(n_1150), .B(n_1178), .Y(n_1189) );
OAI21xp33_ASAP7_75t_L g1205 ( .A1(n_1150), .A2(n_1206), .B(n_1207), .Y(n_1205) );
OR2x2_ASAP7_75t_L g1227 ( .A(n_1150), .B(n_1179), .Y(n_1227) );
INVx2_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
OR2x2_ASAP7_75t_L g1158 ( .A(n_1151), .B(n_1159), .Y(n_1158) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1151), .B(n_1159), .Y(n_1168) );
NAND2xp5_ASAP7_75t_L g1208 ( .A(n_1151), .B(n_1209), .Y(n_1208) );
NAND2x1p5_ASAP7_75t_L g1151 ( .A(n_1152), .B(n_1153), .Y(n_1151) );
OAI21xp5_ASAP7_75t_SL g1154 ( .A1(n_1155), .A2(n_1162), .B(n_1169), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
NAND3xp33_ASAP7_75t_SL g1290 ( .A(n_1156), .B(n_1286), .C(n_1291), .Y(n_1290) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1285 ( .A(n_1157), .B(n_1164), .Y(n_1285) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1158), .Y(n_1224) );
OR2x2_ASAP7_75t_L g1265 ( .A(n_1158), .B(n_1244), .Y(n_1265) );
OR2x2_ASAP7_75t_L g1273 ( .A(n_1158), .B(n_1178), .Y(n_1273) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1159), .Y(n_1204) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1159), .Y(n_1209) );
NAND2xp5_ASAP7_75t_L g1236 ( .A(n_1159), .B(n_1179), .Y(n_1236) );
OAI32xp33_ASAP7_75t_L g1301 ( .A1(n_1159), .A2(n_1188), .A3(n_1235), .B1(n_1240), .B2(n_1302), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_1160), .B(n_1161), .Y(n_1159) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
NOR2xp33_ASAP7_75t_L g1296 ( .A(n_1163), .B(n_1228), .Y(n_1296) );
OR2x2_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1167), .Y(n_1163) );
OR2x2_ASAP7_75t_L g1207 ( .A(n_1164), .B(n_1208), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1164), .B(n_1183), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1165), .B(n_1166), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1165), .B(n_1166), .Y(n_1179) );
NOR2x1_ASAP7_75t_L g1176 ( .A(n_1167), .B(n_1177), .Y(n_1176) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
NAND2xp5_ASAP7_75t_L g1242 ( .A(n_1168), .B(n_1243), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1168), .B(n_1276), .Y(n_1275) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
OR2x2_ASAP7_75t_L g1170 ( .A(n_1171), .B(n_1172), .Y(n_1170) );
CKINVDCx14_ASAP7_75t_R g1193 ( .A(n_1171), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1171), .B(n_1196), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1250 ( .A(n_1171), .B(n_1185), .Y(n_1250) );
OR2x2_ASAP7_75t_L g1279 ( .A(n_1171), .B(n_1197), .Y(n_1279) );
OR2x2_ASAP7_75t_L g1306 ( .A(n_1171), .B(n_1192), .Y(n_1306) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1172), .Y(n_1174) );
O2A1O1Ixp33_ASAP7_75t_L g1241 ( .A1(n_1172), .A2(n_1242), .B(n_1245), .C(n_1249), .Y(n_1241) );
NAND2xp5_ASAP7_75t_L g1173 ( .A(n_1174), .B(n_1175), .Y(n_1173) );
OAI21xp5_ASAP7_75t_L g1297 ( .A1(n_1175), .A2(n_1193), .B(n_1298), .Y(n_1297) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1178), .Y(n_1175) );
NOR2xp33_ASAP7_75t_L g1257 ( .A(n_1177), .B(n_1233), .Y(n_1257) );
CKINVDCx5p33_ASAP7_75t_R g1259 ( .A(n_1177), .Y(n_1259) );
O2A1O1Ixp33_ASAP7_75t_SL g1284 ( .A1(n_1177), .A2(n_1227), .B(n_1285), .C(n_1286), .Y(n_1284) );
NAND2xp5_ASAP7_75t_L g1308 ( .A(n_1177), .B(n_1215), .Y(n_1308) );
OAI221xp5_ASAP7_75t_L g1180 ( .A1(n_1178), .A2(n_1181), .B1(n_1193), .B2(n_1194), .C(n_1198), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1178), .B(n_1183), .Y(n_1182) );
OR2x2_ASAP7_75t_L g1248 ( .A(n_1178), .B(n_1208), .Y(n_1248) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
OR2x2_ASAP7_75t_L g1203 ( .A(n_1179), .B(n_1204), .Y(n_1203) );
AOI22xp5_ASAP7_75t_SL g1181 ( .A1(n_1182), .A2(n_1184), .B1(n_1186), .B2(n_1190), .Y(n_1181) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1182), .Y(n_1270) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1183), .Y(n_1256) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1184), .Y(n_1210) );
INVx2_ASAP7_75t_L g1225 ( .A(n_1185), .Y(n_1225) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1185), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1185), .B(n_1192), .Y(n_1260) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
HB1xp67_ASAP7_75t_L g1188 ( .A(n_1189), .Y(n_1188) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1191), .Y(n_1190) );
NAND2xp5_ASAP7_75t_SL g1229 ( .A(n_1191), .B(n_1230), .Y(n_1229) );
INVx2_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
NOR2xp33_ASAP7_75t_L g1264 ( .A(n_1192), .B(n_1265), .Y(n_1264) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
AOI22xp5_ASAP7_75t_L g1304 ( .A1(n_1195), .A2(n_1238), .B1(n_1246), .B2(n_1305), .Y(n_1304) );
O2A1O1Ixp33_ASAP7_75t_L g1300 ( .A1(n_1196), .A2(n_1246), .B(n_1263), .C(n_1301), .Y(n_1300) );
CKINVDCx5p33_ASAP7_75t_R g1196 ( .A(n_1197), .Y(n_1196) );
AOI221xp5_ASAP7_75t_L g1198 ( .A1(n_1199), .A2(n_1202), .B1(n_1205), .B2(n_1210), .C(n_1211), .Y(n_1198) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1201), .Y(n_1280) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
AOI22xp5_ASAP7_75t_L g1253 ( .A1(n_1204), .A2(n_1254), .B1(n_1257), .B2(n_1258), .Y(n_1253) );
NAND2xp5_ASAP7_75t_L g1255 ( .A(n_1208), .B(n_1256), .Y(n_1255) );
NAND2xp5_ASAP7_75t_L g1302 ( .A(n_1210), .B(n_1303), .Y(n_1302) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1212), .B(n_1221), .Y(n_1211) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1212), .Y(n_1281) );
INVx2_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
OAI221xp5_ASAP7_75t_L g1215 ( .A1(n_1216), .A2(n_1217), .B1(n_1218), .B2(n_1219), .C(n_1220), .Y(n_1215) );
NAND3xp33_ASAP7_75t_L g1221 ( .A(n_1222), .B(n_1224), .C(n_1225), .Y(n_1221) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1224), .B(n_1276), .Y(n_1295) );
OAI211xp5_ASAP7_75t_L g1226 ( .A1(n_1227), .A2(n_1228), .B(n_1229), .C(n_1232), .Y(n_1226) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1236), .Y(n_1238) );
CKINVDCx14_ASAP7_75t_R g1239 ( .A(n_1240), .Y(n_1239) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1244), .Y(n_1243) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1248), .Y(n_1247) );
AOI21xp5_ASAP7_75t_L g1278 ( .A1(n_1248), .A2(n_1279), .B(n_1280), .Y(n_1278) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1250), .Y(n_1249) );
AOI21xp5_ASAP7_75t_L g1251 ( .A1(n_1252), .A2(n_1281), .B(n_1282), .Y(n_1251) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1259), .B(n_1260), .Y(n_1258) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1260), .Y(n_1307) );
AOI211xp5_ASAP7_75t_L g1261 ( .A1(n_1262), .A2(n_1263), .B(n_1264), .C(n_1266), .Y(n_1261) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1262), .Y(n_1269) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1265), .Y(n_1294) );
AOI21xp33_ASAP7_75t_L g1266 ( .A1(n_1267), .A2(n_1269), .B(n_1270), .Y(n_1266) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
NAND2xp5_ASAP7_75t_L g1272 ( .A(n_1273), .B(n_1274), .Y(n_1272) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
NAND5xp2_ASAP7_75t_SL g1282 ( .A(n_1283), .B(n_1293), .C(n_1297), .D(n_1300), .E(n_1304), .Y(n_1282) );
OAI21xp5_ASAP7_75t_SL g1283 ( .A1(n_1284), .A2(n_1288), .B(n_1290), .Y(n_1283) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
INVxp67_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1295), .Y(n_1299) );
AOI21xp33_ASAP7_75t_L g1305 ( .A1(n_1306), .A2(n_1307), .B(n_1308), .Y(n_1305) );
INVx4_ASAP7_75t_L g1309 ( .A(n_1310), .Y(n_1309) );
CKINVDCx20_ASAP7_75t_R g1311 ( .A(n_1312), .Y(n_1311) );
CKINVDCx20_ASAP7_75t_R g1312 ( .A(n_1313), .Y(n_1312) );
INVx3_ASAP7_75t_L g1313 ( .A(n_1314), .Y(n_1313) );
BUFx3_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
NAND3xp33_ASAP7_75t_L g1318 ( .A(n_1319), .B(n_1358), .C(n_1372), .Y(n_1318) );
NOR2xp33_ASAP7_75t_L g1319 ( .A(n_1320), .B(n_1345), .Y(n_1319) );
OAI33xp33_ASAP7_75t_L g1320 ( .A1(n_1321), .A2(n_1323), .A3(n_1328), .B1(n_1334), .B2(n_1338), .B3(n_1343), .Y(n_1320) );
BUFx6f_ASAP7_75t_L g1321 ( .A(n_1322), .Y(n_1321) );
OAI22xp33_ASAP7_75t_L g1346 ( .A1(n_1324), .A2(n_1336), .B1(n_1347), .B2(n_1350), .Y(n_1346) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
OAI22xp33_ASAP7_75t_L g1355 ( .A1(n_1327), .A2(n_1337), .B1(n_1347), .B2(n_1356), .Y(n_1355) );
INVx2_ASAP7_75t_L g1330 ( .A(n_1331), .Y(n_1330) );
INVx4_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
INVx5_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
CKINVDCx5p33_ASAP7_75t_R g1343 ( .A(n_1344), .Y(n_1343) );
INVx2_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1349), .Y(n_1348) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1351), .Y(n_1350) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
OAI31xp33_ASAP7_75t_L g1358 ( .A1(n_1359), .A2(n_1361), .A3(n_1367), .B(n_1371), .Y(n_1358) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1370), .Y(n_1369) );
INVx2_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1380), .Y(n_1379) );
BUFx2_ASAP7_75t_L g1434 ( .A(n_1380), .Y(n_1434) );
INVx2_ASAP7_75t_L g1386 ( .A(n_1387), .Y(n_1386) );
BUFx3_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
BUFx3_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
INVxp33_ASAP7_75t_L g1392 ( .A(n_1393), .Y(n_1392) );
HB1xp67_ASAP7_75t_L g1394 ( .A(n_1395), .Y(n_1394) );
NAND3xp33_ASAP7_75t_L g1395 ( .A(n_1396), .B(n_1415), .C(n_1418), .Y(n_1395) );
NOR3xp33_ASAP7_75t_L g1396 ( .A(n_1397), .B(n_1413), .C(n_1414), .Y(n_1396) );
NAND2xp5_ASAP7_75t_L g1397 ( .A(n_1398), .B(n_1402), .Y(n_1397) );
INVx2_ASAP7_75t_L g1406 ( .A(n_1407), .Y(n_1406) );
INVx8_ASAP7_75t_L g1410 ( .A(n_1411), .Y(n_1410) );
OAI21xp5_ASAP7_75t_L g1418 ( .A1(n_1419), .A2(n_1430), .B(n_1439), .Y(n_1418) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1423), .Y(n_1422) );
INVx1_ASAP7_75t_L g1428 ( .A(n_1429), .Y(n_1428) );
NAND2xp5_ASAP7_75t_L g1431 ( .A(n_1432), .B(n_1437), .Y(n_1431) );
INVx2_ASAP7_75t_L g1433 ( .A(n_1434), .Y(n_1433) );
INVx2_ASAP7_75t_L g1439 ( .A(n_1440), .Y(n_1439) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1444), .Y(n_1443) );
endmodule