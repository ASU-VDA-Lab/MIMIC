module real_jpeg_4536_n_30 (n_17, n_8, n_0, n_21, n_168, n_2, n_29, n_10, n_175, n_9, n_12, n_24, n_170, n_176, n_6, n_28, n_171, n_169, n_177, n_23, n_11, n_14, n_172, n_25, n_7, n_22, n_18, n_3, n_174, n_5, n_4, n_173, n_1, n_26, n_27, n_20, n_19, n_16, n_15, n_13, n_30);

input n_17;
input n_8;
input n_0;
input n_21;
input n_168;
input n_2;
input n_29;
input n_10;
input n_175;
input n_9;
input n_12;
input n_24;
input n_170;
input n_176;
input n_6;
input n_28;
input n_171;
input n_169;
input n_177;
input n_23;
input n_11;
input n_14;
input n_172;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_174;
input n_5;
input n_4;
input n_173;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_16;
input n_15;
input n_13;

output n_30;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_131;
wire n_47;
wire n_163;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_150;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_0),
.B(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_1),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_2),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_2),
.B(n_131),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_3),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_4),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_4),
.B(n_122),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_5),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_5),
.B(n_64),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_6),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_7),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_8),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_9),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_11),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_12),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_12),
.B(n_109),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_14),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_14),
.B(n_71),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_16),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_16),
.B(n_54),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_17),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_17),
.B(n_96),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_18),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_18),
.B(n_58),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_19),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_20),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_21),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_22),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_23),
.B(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_24),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_25),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_26),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_26),
.B(n_75),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_27),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_27),
.B(n_152),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_28),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_28),
.B(n_48),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_29),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_29),
.B(n_148),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_29),
.B(n_41),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_29),
.B(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_161),
.Y(n_30)
);

AO21x1_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_39),
.B(n_160),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_38),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_33),
.B(n_38),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_42),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_36),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_38),
.B(n_166),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_43),
.B(n_159),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_146),
.B(n_156),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_124),
.B(n_140),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_66),
.B(n_112),
.C(n_121),
.Y(n_45)
);

NOR4xp25_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_53),
.C(n_57),
.D(n_63),
.Y(n_46)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_52),
.Y(n_150)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_53),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_105),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_57),
.A2(n_116),
.B(n_117),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_60),
.B(n_110),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_60),
.B(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_60),
.B(n_164),
.Y(n_163)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_89),
.Y(n_88)
);

OAI21x1_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_108),
.B(n_111),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_103),
.B(n_107),
.Y(n_67)
);

AO221x1_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_78),
.B1(n_100),
.B2(n_101),
.C(n_102),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_74),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

AO21x1_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_85),
.B(n_99),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_84),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_84),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_123),
.Y(n_122)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_95),
.B(n_98),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_90),
.B(n_94),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_93),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_93),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_106),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_106),
.Y(n_107)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

A2O1A1O1Ixp25_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B(n_118),
.C(n_119),
.D(n_120),
.Y(n_113)
);

NAND3xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_129),
.C(n_134),
.Y(n_124)
);

A2O1A1O1Ixp25_ASAP7_75t_L g140 ( 
.A1(n_125),
.A2(n_134),
.B(n_141),
.C(n_144),
.D(n_145),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_127),
.Y(n_145)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_130),
.A2(n_142),
.B(n_143),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_133),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_139),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_139),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_L g156 ( 
.A1(n_151),
.A2(n_157),
.B(n_158),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_163),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_168),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_169),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_170),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_171),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_172),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_173),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_174),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_175),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_176),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_177),
.Y(n_110)
);


endmodule