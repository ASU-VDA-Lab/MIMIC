module fake_netlist_5_1283_n_1731 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1731);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1731;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1633;
wire n_1236;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1363;
wire n_1668;
wire n_1301;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1439;
wire n_1312;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1478;
wire n_1339;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_139),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_128),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_1),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_50),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_159),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_68),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_136),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_167),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_37),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_32),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_120),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_123),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_69),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_107),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_26),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_14),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_25),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_91),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_67),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_165),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_84),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_23),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_5),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_48),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_112),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_96),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_121),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_1),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_83),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_103),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_88),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_23),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_114),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_5),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_95),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_20),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_109),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_147),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_61),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_48),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_25),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_97),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_146),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_29),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_122),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_110),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_115),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_161),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_26),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_102),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_33),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_24),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_134),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_89),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_86),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_49),
.Y(n_227)
);

BUFx2_ASAP7_75t_SL g228 ( 
.A(n_137),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_141),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_111),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_59),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_53),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_85),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_58),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_14),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_155),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_78),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_71),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_15),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_164),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_92),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_148),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_135),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_133),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_99),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_150),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_3),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_129),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_31),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_149),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_163),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_34),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_8),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_118),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_81),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_76),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_74),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_62),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_168),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_21),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_33),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_131),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_58),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_27),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_32),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_94),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_156),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_113),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_15),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_152),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_166),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_7),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_11),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_47),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_125),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_57),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_19),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_38),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_66),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_73),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_70),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_82),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_45),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_35),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_126),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_50),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_39),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_130),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_10),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_53),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_9),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_116),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_12),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_55),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_41),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_162),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_38),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_36),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_19),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_63),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_65),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_54),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_57),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_4),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_80),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_45),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_157),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_56),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_105),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_29),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_20),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_27),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_7),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_44),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_51),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_154),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_55),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_21),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_37),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_0),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_142),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_54),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_49),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_79),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_51),
.Y(n_325)
);

BUFx10_ASAP7_75t_L g326 ( 
.A(n_30),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_17),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_4),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_34),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_108),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_13),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_46),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_17),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_39),
.Y(n_334)
);

INVx2_ASAP7_75t_SL g335 ( 
.A(n_30),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_143),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_41),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_101),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_187),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_187),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_170),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_171),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_242),
.B(n_0),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_242),
.B(n_224),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_187),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_218),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_177),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_224),
.B(n_300),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_300),
.B(n_2),
.Y(n_349)
);

CKINVDCx14_ASAP7_75t_R g350 ( 
.A(n_297),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_187),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_187),
.Y(n_352)
);

INVxp33_ASAP7_75t_L g353 ( 
.A(n_180),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_266),
.Y(n_354)
);

BUFx6f_ASAP7_75t_SL g355 ( 
.A(n_181),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_178),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_247),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_297),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_182),
.Y(n_359)
);

INVxp33_ASAP7_75t_SL g360 ( 
.A(n_186),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_288),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_247),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_247),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_183),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_247),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_254),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_247),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_254),
.Y(n_368)
);

NOR2xp67_ASAP7_75t_L g369 ( 
.A(n_276),
.B(n_2),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_252),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_252),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_184),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_252),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_252),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_332),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_252),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_255),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_298),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_332),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_298),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_255),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_188),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_190),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_191),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_326),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_195),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_298),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_326),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_298),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_169),
.B(n_3),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_196),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_197),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_298),
.Y(n_393)
);

INVxp33_ASAP7_75t_SL g394 ( 
.A(n_179),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_172),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_326),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_199),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_201),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_206),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_208),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_210),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_172),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_215),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_215),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_216),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_235),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_217),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_235),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_219),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_221),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_239),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_192),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_181),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_193),
.Y(n_414)
);

INVxp33_ASAP7_75t_SL g415 ( 
.A(n_194),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_198),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_239),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_233),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_236),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_304),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_304),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_237),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_238),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_240),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_339),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_341),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_346),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_375),
.Y(n_428)
);

OA21x2_ASAP7_75t_L g429 ( 
.A1(n_339),
.A2(n_173),
.B(n_169),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_340),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_340),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_385),
.B(n_326),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_354),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_342),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_345),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_345),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_347),
.Y(n_437)
);

OAI21x1_ASAP7_75t_L g438 ( 
.A1(n_351),
.A2(n_279),
.B(n_257),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_351),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_361),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_352),
.Y(n_441)
);

NOR2xp67_ASAP7_75t_L g442 ( 
.A(n_352),
.B(n_243),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_357),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_379),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_348),
.B(n_241),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_357),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_362),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_356),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_362),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_366),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_363),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_413),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_363),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_359),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_365),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_365),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_364),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_367),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_367),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_412),
.Y(n_460)
);

OA21x2_ASAP7_75t_L g461 ( 
.A1(n_370),
.A2(n_176),
.B(n_173),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_370),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_383),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_386),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_371),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_414),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_371),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_373),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_373),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_374),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_374),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_376),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_397),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_372),
.Y(n_474)
);

INVx5_ASAP7_75t_L g475 ( 
.A(n_413),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_382),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_376),
.Y(n_477)
);

OA21x2_ASAP7_75t_L g478 ( 
.A1(n_378),
.A2(n_189),
.B(n_176),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_378),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_380),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_384),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_391),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_392),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_380),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_398),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_405),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_399),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_387),
.B(n_181),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_344),
.B(n_245),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_387),
.B(n_251),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_400),
.Y(n_491)
);

NAND2xp33_ASAP7_75t_R g492 ( 
.A(n_360),
.B(n_205),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_389),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_389),
.Y(n_494)
);

OA21x2_ASAP7_75t_L g495 ( 
.A1(n_393),
.A2(n_200),
.B(n_189),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_401),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_349),
.B(n_246),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_393),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_395),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_395),
.Y(n_500)
);

CKINVDCx6p67_ASAP7_75t_R g501 ( 
.A(n_418),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_430),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_445),
.B(n_407),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_488),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_430),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_428),
.B(n_416),
.Y(n_506)
);

AND2x6_ASAP7_75t_L g507 ( 
.A(n_490),
.B(n_251),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_497),
.B(n_257),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_L g509 ( 
.A1(n_497),
.A2(n_343),
.B1(n_390),
.B2(n_350),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_488),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_489),
.B(n_394),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_488),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_501),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_452),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_489),
.A2(n_358),
.B1(n_369),
.B2(n_234),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_488),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_445),
.B(n_409),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_430),
.Y(n_518)
);

BUFx10_ASAP7_75t_L g519 ( 
.A(n_426),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_441),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_452),
.B(n_279),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_460),
.B(n_415),
.Y(n_522)
);

NAND2xp33_ASAP7_75t_L g523 ( 
.A(n_490),
.B(n_316),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_460),
.B(n_410),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_441),
.Y(n_525)
);

INVx4_ASAP7_75t_L g526 ( 
.A(n_475),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_466),
.B(n_419),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_452),
.B(n_338),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_427),
.B(n_368),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g530 ( 
.A(n_450),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_475),
.B(n_422),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_435),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_466),
.B(n_423),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_441),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_475),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_501),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_431),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_431),
.Y(n_538)
);

NAND2x1p5_ASAP7_75t_L g539 ( 
.A(n_475),
.B(n_251),
.Y(n_539)
);

INVx5_ASAP7_75t_L g540 ( 
.A(n_425),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_449),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_490),
.B(n_402),
.Y(n_542)
);

INVx1_ASAP7_75t_SL g543 ( 
.A(n_463),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_475),
.Y(n_544)
);

INVx5_ASAP7_75t_L g545 ( 
.A(n_425),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_434),
.B(n_424),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_449),
.Y(n_547)
);

AO22x2_ASAP7_75t_L g548 ( 
.A1(n_432),
.A2(n_234),
.B1(n_335),
.B2(n_202),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_492),
.A2(n_381),
.B1(n_377),
.B2(n_388),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_492),
.A2(n_396),
.B1(n_355),
.B2(n_213),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_475),
.B(n_175),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_475),
.B(n_338),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_436),
.Y(n_553)
);

INVx6_ASAP7_75t_L g554 ( 
.A(n_435),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_442),
.B(n_443),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_443),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_428),
.B(n_353),
.Y(n_557)
);

AND2x6_ASAP7_75t_L g558 ( 
.A(n_446),
.B(n_200),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_446),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_442),
.B(n_256),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_435),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_501),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_429),
.A2(n_335),
.B1(n_315),
.B2(n_319),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_437),
.A2(n_448),
.B1(n_457),
.B2(n_454),
.Y(n_564)
);

INVxp67_ASAP7_75t_SL g565 ( 
.A(n_435),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_449),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_435),
.Y(n_567)
);

OR2x6_ASAP7_75t_L g568 ( 
.A(n_444),
.B(n_228),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_474),
.B(n_316),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_435),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_429),
.A2(n_315),
.B1(n_319),
.B2(n_325),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_439),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_476),
.B(n_355),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_481),
.B(n_355),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_482),
.B(n_316),
.Y(n_575)
);

AND2x6_ASAP7_75t_L g576 ( 
.A(n_451),
.B(n_203),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_483),
.B(n_316),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_485),
.B(n_324),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_451),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_456),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_487),
.B(n_207),
.Y(n_581)
);

INVx5_ASAP7_75t_L g582 ( 
.A(n_425),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_491),
.B(n_316),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_455),
.Y(n_584)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_439),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_439),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_496),
.B(n_212),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_439),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_439),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_455),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_444),
.B(n_253),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_450),
.B(n_322),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_500),
.B(n_402),
.Y(n_593)
);

NOR3xp33_ASAP7_75t_L g594 ( 
.A(n_500),
.B(n_269),
.C(n_265),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_499),
.B(n_203),
.Y(n_595)
);

AND2x2_ASAP7_75t_SL g596 ( 
.A(n_429),
.B(n_204),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_456),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_458),
.B(n_272),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_433),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_455),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_447),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_429),
.A2(n_258),
.B1(n_275),
.B2(n_270),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_499),
.B(n_403),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_458),
.B(n_467),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_499),
.B(n_204),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_470),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_447),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_459),
.Y(n_608)
);

BUFx10_ASAP7_75t_L g609 ( 
.A(n_498),
.Y(n_609)
);

BUFx10_ASAP7_75t_L g610 ( 
.A(n_498),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_459),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_429),
.A2(n_325),
.B1(n_223),
.B2(n_323),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_447),
.Y(n_613)
);

INVx4_ASAP7_75t_L g614 ( 
.A(n_447),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_470),
.B(n_209),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_440),
.Y(n_616)
);

A2O1A1Ixp33_ASAP7_75t_L g617 ( 
.A1(n_438),
.A2(n_223),
.B(n_314),
.C(n_277),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_464),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_477),
.B(n_209),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_447),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_477),
.A2(n_286),
.B1(n_278),
.B2(n_283),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_447),
.Y(n_622)
);

NOR2x1p5_ASAP7_75t_L g623 ( 
.A(n_479),
.B(n_323),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_461),
.A2(n_223),
.B1(n_174),
.B2(n_334),
.Y(n_624)
);

BUFx4f_ASAP7_75t_L g625 ( 
.A(n_461),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_479),
.B(n_214),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_459),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_484),
.B(n_248),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_484),
.B(n_214),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_494),
.B(n_250),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_494),
.B(n_225),
.Y(n_631)
);

BUFx4f_ASAP7_75t_L g632 ( 
.A(n_461),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_465),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_493),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_493),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_465),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_465),
.Y(n_637)
);

INVx1_ASAP7_75t_SL g638 ( 
.A(n_473),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_468),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_453),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_493),
.B(n_267),
.Y(n_641)
);

INVx4_ASAP7_75t_L g642 ( 
.A(n_453),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_453),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_453),
.B(n_268),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_461),
.A2(n_261),
.B1(n_185),
.B2(n_334),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_461),
.A2(n_261),
.B1(n_185),
.B2(n_202),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_462),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_462),
.B(n_280),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_616),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_596),
.A2(n_495),
.B1(n_478),
.B2(n_264),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_511),
.B(n_478),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_504),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_578),
.B(n_281),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_502),
.Y(n_654)
);

OAI221xp5_ASAP7_75t_L g655 ( 
.A1(n_509),
.A2(n_314),
.B1(n_227),
.B2(n_277),
.C(n_222),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_514),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_503),
.B(n_478),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_502),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_514),
.Y(n_659)
);

NAND3xp33_ASAP7_75t_L g660 ( 
.A(n_515),
.B(n_294),
.C(n_274),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_517),
.B(n_478),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_623),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_596),
.A2(n_495),
.B1(n_478),
.B2(n_174),
.Y(n_663)
);

INVxp67_ASAP7_75t_L g664 ( 
.A(n_557),
.Y(n_664)
);

OAI22xp5_ASAP7_75t_L g665 ( 
.A1(n_510),
.A2(n_259),
.B1(n_336),
.B2(n_262),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_512),
.B(n_495),
.Y(n_666)
);

INVxp67_ASAP7_75t_L g667 ( 
.A(n_591),
.Y(n_667)
);

NAND3xp33_ASAP7_75t_L g668 ( 
.A(n_524),
.B(n_533),
.C(n_527),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_516),
.B(n_495),
.Y(n_669)
);

AO221x1_ASAP7_75t_L g670 ( 
.A1(n_548),
.A2(n_295),
.B1(n_227),
.B2(n_232),
.C(n_249),
.Y(n_670)
);

BUFx12f_ASAP7_75t_L g671 ( 
.A(n_519),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_508),
.B(n_495),
.Y(n_672)
);

A2O1A1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_625),
.A2(n_438),
.B(n_230),
.C(n_321),
.Y(n_673)
);

OR2x6_ASAP7_75t_L g674 ( 
.A(n_599),
.B(n_228),
.Y(n_674)
);

INVx8_ASAP7_75t_L g675 ( 
.A(n_568),
.Y(n_675)
);

AND2x6_ASAP7_75t_SL g676 ( 
.A(n_522),
.B(n_220),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_581),
.B(n_587),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_542),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_505),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_550),
.B(n_282),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_609),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_569),
.B(n_284),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_560),
.B(n_285),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_507),
.A2(n_296),
.B1(n_292),
.B2(n_330),
.Y(n_684)
);

AND2x6_ASAP7_75t_SL g685 ( 
.A(n_546),
.B(n_220),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_537),
.B(n_462),
.Y(n_686)
);

INVx4_ASAP7_75t_L g687 ( 
.A(n_567),
.Y(n_687)
);

INVx6_ASAP7_75t_L g688 ( 
.A(n_609),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_505),
.Y(n_689)
);

NOR3x1_ASAP7_75t_L g690 ( 
.A(n_530),
.B(n_249),
.C(n_222),
.Y(n_690)
);

BUFx6f_ASAP7_75t_SL g691 ( 
.A(n_519),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_569),
.B(n_287),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_542),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_571),
.A2(n_264),
.B1(n_273),
.B2(n_232),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_609),
.B(n_301),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_616),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_575),
.B(n_290),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_538),
.B(n_462),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_575),
.B(n_291),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_645),
.A2(n_320),
.B1(n_318),
.B2(n_311),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_610),
.B(n_305),
.Y(n_701)
);

INVxp67_ASAP7_75t_L g702 ( 
.A(n_592),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_518),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_593),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_553),
.B(n_425),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_610),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_556),
.Y(n_707)
);

AOI221xp5_ASAP7_75t_L g708 ( 
.A1(n_548),
.A2(n_211),
.B1(n_260),
.B2(n_337),
.C(n_263),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_559),
.B(n_425),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_579),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_577),
.B(n_293),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_SL g712 ( 
.A(n_519),
.B(n_486),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_580),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_597),
.Y(n_714)
);

NOR2xp67_ASAP7_75t_L g715 ( 
.A(n_564),
.B(n_307),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_577),
.B(n_299),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_606),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_604),
.B(n_555),
.Y(n_718)
);

AND2x6_ASAP7_75t_SL g719 ( 
.A(n_568),
.B(n_273),
.Y(n_719)
);

BUFx6f_ASAP7_75t_SL g720 ( 
.A(n_568),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_646),
.A2(n_320),
.B1(n_289),
.B2(n_295),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_628),
.B(n_630),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_518),
.Y(n_723)
);

A2O1A1Ixp33_ASAP7_75t_L g724 ( 
.A1(n_625),
.A2(n_438),
.B(n_226),
.C(n_259),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_603),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_520),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_507),
.B(n_425),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_506),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_583),
.B(n_302),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_507),
.B(n_469),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_520),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_525),
.Y(n_732)
);

BUFx2_ASAP7_75t_L g733 ( 
.A(n_568),
.Y(n_733)
);

A2O1A1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_625),
.A2(n_321),
.B(n_229),
.C(n_230),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_534),
.Y(n_735)
);

O2A1O1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_617),
.A2(n_318),
.B(n_311),
.C(n_289),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_573),
.B(n_403),
.Y(n_737)
);

OAI21xp33_ASAP7_75t_L g738 ( 
.A1(n_548),
.A2(n_328),
.B(n_303),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_583),
.B(n_306),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_610),
.B(n_226),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_SL g741 ( 
.A(n_513),
.B(n_331),
.Y(n_741)
);

BUFx3_ASAP7_75t_L g742 ( 
.A(n_558),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_634),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_574),
.B(n_229),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_541),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_507),
.B(n_469),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_594),
.B(n_231),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_521),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_598),
.B(n_231),
.Y(n_749)
);

NAND2xp33_ASAP7_75t_L g750 ( 
.A(n_558),
.B(n_244),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_641),
.B(n_308),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_602),
.B(n_549),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_624),
.A2(n_336),
.B1(n_262),
.B2(n_271),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_547),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_547),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_635),
.B(n_469),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_566),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_632),
.B(n_244),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_566),
.Y(n_759)
);

OR2x2_ASAP7_75t_L g760 ( 
.A(n_543),
.B(n_310),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_521),
.B(n_312),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_528),
.B(n_313),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_528),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_563),
.B(n_469),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_565),
.B(n_469),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_567),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_632),
.B(n_469),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_621),
.B(n_317),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_584),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_632),
.B(n_271),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_644),
.B(n_309),
.Y(n_771)
);

A2O1A1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_617),
.A2(n_612),
.B(n_523),
.C(n_595),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_584),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_648),
.B(n_309),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_590),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_590),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_600),
.Y(n_777)
);

BUFx8_ASAP7_75t_L g778 ( 
.A(n_513),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_615),
.B(n_327),
.Y(n_779)
);

NAND2xp33_ASAP7_75t_L g780 ( 
.A(n_558),
.B(n_329),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_558),
.A2(n_576),
.B1(n_523),
.B2(n_551),
.Y(n_781)
);

INVx8_ASAP7_75t_L g782 ( 
.A(n_558),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_558),
.A2(n_333),
.B1(n_480),
.B2(n_471),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_532),
.B(n_480),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_600),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_615),
.B(n_6),
.Y(n_786)
);

NOR3xp33_ASAP7_75t_L g787 ( 
.A(n_638),
.B(n_420),
.C(n_406),
.Y(n_787)
);

O2A1O1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_619),
.A2(n_420),
.B(n_406),
.C(n_408),
.Y(n_788)
);

O2A1O1Ixp5_ASAP7_75t_L g789 ( 
.A1(n_619),
.A2(n_480),
.B(n_472),
.C(n_471),
.Y(n_789)
);

NAND2x1p5_ASAP7_75t_L g790 ( 
.A(n_595),
.B(n_472),
.Y(n_790)
);

NOR2x1p5_ASAP7_75t_L g791 ( 
.A(n_536),
.B(n_417),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_608),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_611),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_618),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_SL g795 ( 
.A(n_536),
.B(n_417),
.Y(n_795)
);

INVxp33_ASAP7_75t_L g796 ( 
.A(n_529),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_611),
.Y(n_797)
);

AND2x6_ASAP7_75t_SL g798 ( 
.A(n_618),
.B(n_404),
.Y(n_798)
);

NOR3xp33_ASAP7_75t_L g799 ( 
.A(n_562),
.B(n_421),
.C(n_411),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_626),
.B(n_6),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_627),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_627),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_562),
.B(n_539),
.Y(n_803)
);

NAND2x1_ASAP7_75t_L g804 ( 
.A(n_554),
.B(n_472),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_626),
.B(n_8),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_633),
.Y(n_806)
);

AND2x6_ASAP7_75t_SL g807 ( 
.A(n_531),
.B(n_404),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_532),
.B(n_471),
.Y(n_808)
);

BUFx12f_ASAP7_75t_SL g809 ( 
.A(n_567),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_532),
.B(n_468),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_718),
.B(n_576),
.Y(n_811)
);

AOI21xp33_ASAP7_75t_L g812 ( 
.A1(n_677),
.A2(n_629),
.B(n_631),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_764),
.A2(n_552),
.B(n_526),
.Y(n_813)
);

OAI21xp5_ASAP7_75t_L g814 ( 
.A1(n_657),
.A2(n_636),
.B(n_633),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_664),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_677),
.B(n_576),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_667),
.B(n_408),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_L g818 ( 
.A1(n_661),
.A2(n_637),
.B(n_636),
.Y(n_818)
);

AOI21x1_ASAP7_75t_L g819 ( 
.A1(n_666),
.A2(n_639),
.B(n_637),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_668),
.B(n_570),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_752),
.A2(n_576),
.B1(n_588),
.B2(n_647),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_722),
.B(n_751),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_652),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_682),
.A2(n_631),
.B(n_629),
.C(n_605),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_770),
.A2(n_544),
.B(n_526),
.Y(n_825)
);

A2O1A1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_682),
.A2(n_605),
.B(n_640),
.C(n_561),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_681),
.B(n_706),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_654),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_654),
.Y(n_829)
);

NAND2x1p5_ASAP7_75t_L g830 ( 
.A(n_681),
.B(n_588),
.Y(n_830)
);

O2A1O1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_655),
.A2(n_639),
.B(n_468),
.C(n_539),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_727),
.A2(n_586),
.B(n_643),
.Y(n_832)
);

OAI21xp33_ASAP7_75t_L g833 ( 
.A1(n_768),
.A2(n_411),
.B(n_421),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_730),
.A2(n_585),
.B(n_643),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_746),
.A2(n_586),
.B(n_642),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_651),
.A2(n_753),
.B1(n_758),
.B2(n_663),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_737),
.B(n_753),
.Y(n_837)
);

O2A1O1Ixp33_ASAP7_75t_SL g838 ( 
.A1(n_734),
.A2(n_561),
.B(n_601),
.C(n_640),
.Y(n_838)
);

OR2x2_ASAP7_75t_L g839 ( 
.A(n_728),
.B(n_9),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_650),
.A2(n_561),
.B1(n_640),
.B2(n_601),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_702),
.B(n_795),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_765),
.A2(n_585),
.B(n_642),
.Y(n_842)
);

OAI21xp5_ASAP7_75t_L g843 ( 
.A1(n_672),
.A2(n_601),
.B(n_576),
.Y(n_843)
);

AOI21x1_ASAP7_75t_L g844 ( 
.A1(n_669),
.A2(n_647),
.B(n_607),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_707),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_681),
.B(n_567),
.Y(n_846)
);

NAND2x1p5_ASAP7_75t_L g847 ( 
.A(n_681),
.B(n_620),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_687),
.A2(n_614),
.B(n_613),
.Y(n_848)
);

AO21x1_ASAP7_75t_L g849 ( 
.A1(n_749),
.A2(n_613),
.B(n_614),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_725),
.B(n_607),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_760),
.B(n_620),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_782),
.A2(n_535),
.B(n_589),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_710),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_678),
.B(n_622),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_706),
.B(n_589),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_658),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_663),
.A2(n_622),
.B(n_589),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_766),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_771),
.A2(n_622),
.B(n_572),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_673),
.A2(n_724),
.B(n_781),
.Y(n_860)
);

BUFx8_ASAP7_75t_L g861 ( 
.A(n_691),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_693),
.B(n_713),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_714),
.B(n_622),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_774),
.A2(n_698),
.B(n_686),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_656),
.Y(n_865)
);

AO21x1_ASAP7_75t_L g866 ( 
.A1(n_786),
.A2(n_10),
.B(n_11),
.Y(n_866)
);

AO22x1_ASAP7_75t_L g867 ( 
.A1(n_768),
.A2(n_12),
.B1(n_13),
.B2(n_16),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_717),
.B(n_554),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_705),
.A2(n_582),
.B(n_545),
.Y(n_869)
);

NAND3xp33_ASAP7_75t_L g870 ( 
.A(n_708),
.B(n_697),
.C(n_692),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_748),
.B(n_582),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_709),
.A2(n_582),
.B(n_545),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_704),
.B(n_16),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_694),
.B(n_582),
.Y(n_874)
);

O2A1O1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_786),
.A2(n_18),
.B(n_22),
.C(n_24),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_679),
.Y(n_876)
);

INVx1_ASAP7_75t_SL g877 ( 
.A(n_649),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_694),
.B(n_545),
.Y(n_878)
);

NAND2x1_ASAP7_75t_L g879 ( 
.A(n_766),
.B(n_545),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_766),
.A2(n_545),
.B(n_540),
.Y(n_880)
);

INVxp67_ASAP7_75t_L g881 ( 
.A(n_692),
.Y(n_881)
);

OAI21xp33_ASAP7_75t_L g882 ( 
.A1(n_697),
.A2(n_18),
.B(n_22),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_810),
.A2(n_540),
.B(n_87),
.Y(n_883)
);

BUFx3_ASAP7_75t_L g884 ( 
.A(n_671),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_699),
.B(n_540),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_779),
.B(n_540),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_743),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_784),
.A2(n_540),
.B(n_90),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_699),
.B(n_77),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_688),
.B(n_28),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_690),
.Y(n_891)
);

AOI21x1_ASAP7_75t_L g892 ( 
.A1(n_808),
.A2(n_75),
.B(n_158),
.Y(n_892)
);

NOR3xp33_ASAP7_75t_L g893 ( 
.A(n_680),
.B(n_28),
.C(n_31),
.Y(n_893)
);

AOI22xp5_ASAP7_75t_L g894 ( 
.A1(n_763),
.A2(n_93),
.B1(n_153),
.B2(n_151),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_688),
.A2(n_72),
.B1(n_145),
.B2(n_144),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_779),
.B(n_35),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_688),
.B(n_36),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_756),
.A2(n_98),
.B(n_138),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_653),
.B(n_40),
.Y(n_899)
);

NAND2x1p5_ASAP7_75t_L g900 ( 
.A(n_742),
.B(n_64),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_711),
.B(n_40),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_716),
.B(n_100),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_750),
.A2(n_60),
.B(n_132),
.Y(n_903)
);

BUFx12f_ASAP7_75t_L g904 ( 
.A(n_798),
.Y(n_904)
);

CKINVDCx10_ASAP7_75t_R g905 ( 
.A(n_691),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_662),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_775),
.A2(n_127),
.B(n_119),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_729),
.A2(n_117),
.B1(n_106),
.B2(n_104),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_777),
.A2(n_42),
.B(n_43),
.Y(n_909)
);

BUFx4f_ASAP7_75t_L g910 ( 
.A(n_671),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_785),
.A2(n_793),
.B(n_797),
.Y(n_911)
);

AO22x1_ASAP7_75t_L g912 ( 
.A1(n_800),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_912)
);

AND2x2_ASAP7_75t_SL g913 ( 
.A(n_712),
.B(n_46),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_679),
.A2(n_47),
.B(n_52),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_689),
.A2(n_52),
.B(n_56),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_729),
.A2(n_739),
.B1(n_762),
.B2(n_761),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_739),
.B(n_761),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_762),
.A2(n_740),
.B1(n_715),
.B2(n_683),
.Y(n_918)
);

OAI22xp33_ASAP7_75t_L g919 ( 
.A1(n_741),
.A2(n_733),
.B1(n_675),
.B2(n_674),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_742),
.A2(n_721),
.B1(n_700),
.B2(n_656),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_700),
.B(n_721),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_703),
.A2(n_755),
.B(n_806),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_723),
.B(n_755),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_723),
.B(n_757),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_726),
.A2(n_757),
.B(n_806),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_731),
.B(n_759),
.Y(n_926)
);

CKINVDCx10_ASAP7_75t_R g927 ( 
.A(n_720),
.Y(n_927)
);

INVx4_ASAP7_75t_L g928 ( 
.A(n_659),
.Y(n_928)
);

A2O1A1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_800),
.A2(n_805),
.B(n_738),
.C(n_736),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_659),
.B(n_796),
.Y(n_930)
);

O2A1O1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_805),
.A2(n_665),
.B(n_747),
.C(n_744),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_732),
.B(n_773),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_732),
.B(n_773),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_789),
.A2(n_769),
.B(n_759),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_791),
.B(n_787),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_695),
.B(n_701),
.Y(n_936)
);

BUFx3_ASAP7_75t_L g937 ( 
.A(n_696),
.Y(n_937)
);

AOI22xp5_ASAP7_75t_L g938 ( 
.A1(n_780),
.A2(n_803),
.B1(n_684),
.B2(n_720),
.Y(n_938)
);

O2A1O1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_788),
.A2(n_776),
.B(n_802),
.C(n_801),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_735),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_675),
.A2(n_783),
.B1(n_790),
.B2(n_792),
.Y(n_941)
);

BUFx4f_ASAP7_75t_L g942 ( 
.A(n_675),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_799),
.B(n_794),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_745),
.B(n_754),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_792),
.A2(n_790),
.B(n_660),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_670),
.B(n_807),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_809),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_804),
.B(n_674),
.Y(n_948)
);

AND2x6_ASAP7_75t_L g949 ( 
.A(n_719),
.B(n_674),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_676),
.B(n_685),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_778),
.A2(n_632),
.B(n_625),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_778),
.A2(n_632),
.B(n_625),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_767),
.A2(n_632),
.B(n_625),
.Y(n_953)
);

OAI321xp33_ASAP7_75t_L g954 ( 
.A1(n_655),
.A2(n_343),
.A3(n_509),
.B1(n_768),
.B2(n_800),
.C(n_786),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_718),
.B(n_677),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_718),
.B(n_677),
.Y(n_956)
);

INVx4_ASAP7_75t_L g957 ( 
.A(n_681),
.Y(n_957)
);

O2A1O1Ixp33_ASAP7_75t_SL g958 ( 
.A1(n_734),
.A2(n_772),
.B(n_724),
.C(n_673),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_681),
.B(n_706),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_767),
.A2(n_632),
.B(n_625),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_668),
.A2(n_677),
.B1(n_651),
.B2(n_718),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_667),
.B(n_677),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_652),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_677),
.A2(n_668),
.B1(n_511),
.B2(n_752),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_667),
.B(n_557),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_718),
.B(n_677),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_767),
.A2(n_632),
.B(n_625),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_718),
.B(n_677),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_718),
.B(n_677),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_677),
.A2(n_511),
.B(n_668),
.C(n_682),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_681),
.B(n_706),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_677),
.A2(n_668),
.B1(n_511),
.B2(n_752),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_654),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_681),
.B(n_706),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_865),
.B(n_928),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_955),
.B(n_956),
.Y(n_976)
);

AOI21x1_ASAP7_75t_L g977 ( 
.A1(n_885),
.A2(n_886),
.B(n_857),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_823),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_966),
.B(n_968),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_969),
.A2(n_964),
.B1(n_972),
.B2(n_916),
.Y(n_980)
);

AND3x4_ASAP7_75t_L g981 ( 
.A(n_937),
.B(n_893),
.C(n_884),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_L g982 ( 
.A1(n_970),
.A2(n_921),
.B1(n_917),
.B2(n_870),
.Y(n_982)
);

INVxp67_ASAP7_75t_L g983 ( 
.A(n_965),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_954),
.A2(n_931),
.B(n_896),
.C(n_962),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_865),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_961),
.B(n_837),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_811),
.A2(n_836),
.B(n_834),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_901),
.A2(n_899),
.B(n_812),
.C(n_929),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_881),
.A2(n_824),
.B(n_820),
.C(n_918),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_832),
.A2(n_835),
.B(n_958),
.Y(n_990)
);

AOI22xp33_ASAP7_75t_SL g991 ( 
.A1(n_913),
.A2(n_841),
.B1(n_949),
.B2(n_935),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_828),
.Y(n_992)
);

INVx4_ASAP7_75t_SL g993 ( 
.A(n_949),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_816),
.B(n_817),
.Y(n_994)
);

AOI221x1_ASAP7_75t_L g995 ( 
.A1(n_860),
.A2(n_882),
.B1(n_864),
.B2(n_946),
.C(n_941),
.Y(n_995)
);

INVx1_ASAP7_75t_SL g996 ( 
.A(n_815),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_891),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_851),
.B(n_963),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_845),
.Y(n_999)
);

OAI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_843),
.A2(n_814),
.B(n_818),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_862),
.B(n_853),
.Y(n_1001)
);

OAI21x1_ASAP7_75t_SL g1002 ( 
.A1(n_951),
.A2(n_952),
.B(n_866),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_887),
.B(n_920),
.Y(n_1003)
);

INVx2_ASAP7_75t_SL g1004 ( 
.A(n_839),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_865),
.B(n_919),
.Y(n_1005)
);

AOI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_936),
.A2(n_930),
.B1(n_938),
.B2(n_943),
.Y(n_1006)
);

BUFx12f_ASAP7_75t_L g1007 ( 
.A(n_861),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_873),
.B(n_850),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_942),
.Y(n_1009)
);

INVx1_ASAP7_75t_SL g1010 ( 
.A(n_877),
.Y(n_1010)
);

INVxp67_ASAP7_75t_L g1011 ( 
.A(n_947),
.Y(n_1011)
);

A2O1A1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_945),
.A2(n_821),
.B(n_875),
.C(n_826),
.Y(n_1012)
);

NAND2xp33_ASAP7_75t_L g1013 ( 
.A(n_830),
.B(n_847),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_957),
.B(n_928),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_854),
.B(n_833),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_957),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_890),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_942),
.A2(n_900),
.B1(n_908),
.B2(n_878),
.Y(n_1018)
);

AO31x2_ASAP7_75t_L g1019 ( 
.A1(n_849),
.A2(n_840),
.A3(n_859),
.B(n_911),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_L g1020 ( 
.A1(n_922),
.A2(n_925),
.B(n_842),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_SL g1021 ( 
.A1(n_909),
.A2(n_907),
.B(n_892),
.Y(n_1021)
);

AND3x2_ASAP7_75t_L g1022 ( 
.A(n_950),
.B(n_897),
.C(n_912),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_858),
.Y(n_1023)
);

OAI21x1_ASAP7_75t_L g1024 ( 
.A1(n_859),
.A2(n_813),
.B(n_848),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_869),
.A2(n_872),
.B(n_939),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_906),
.B(n_910),
.Y(n_1026)
);

NOR2x1_ASAP7_75t_L g1027 ( 
.A(n_827),
.B(n_974),
.Y(n_1027)
);

AOI21xp33_ASAP7_75t_L g1028 ( 
.A1(n_889),
.A2(n_902),
.B(n_948),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_829),
.B(n_973),
.Y(n_1029)
);

AOI21xp33_ASAP7_75t_L g1030 ( 
.A1(n_831),
.A2(n_863),
.B(n_868),
.Y(n_1030)
);

OAI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_923),
.A2(n_924),
.B(n_926),
.Y(n_1031)
);

OAI21xp33_ASAP7_75t_SL g1032 ( 
.A1(n_874),
.A2(n_971),
.B(n_959),
.Y(n_1032)
);

NAND3x1_ASAP7_75t_L g1033 ( 
.A(n_905),
.B(n_927),
.C(n_861),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_932),
.A2(n_944),
.B(n_933),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_910),
.B(n_900),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_856),
.B(n_876),
.Y(n_1036)
);

AO31x2_ASAP7_75t_L g1037 ( 
.A1(n_914),
.A2(n_915),
.A3(n_855),
.B(n_883),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_825),
.A2(n_852),
.B(n_846),
.Y(n_1038)
);

AO31x2_ASAP7_75t_L g1039 ( 
.A1(n_888),
.A2(n_940),
.A3(n_895),
.B(n_903),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_871),
.A2(n_838),
.B(n_830),
.Y(n_1040)
);

INVx4_ASAP7_75t_L g1041 ( 
.A(n_858),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_847),
.A2(n_879),
.B(n_880),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_898),
.A2(n_894),
.B(n_867),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_904),
.B(n_949),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_949),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_955),
.A2(n_966),
.B1(n_968),
.B2(n_956),
.Y(n_1046)
);

O2A1O1Ixp5_ASAP7_75t_L g1047 ( 
.A1(n_970),
.A2(n_917),
.B(n_677),
.C(n_822),
.Y(n_1047)
);

NOR2x1_ASAP7_75t_L g1048 ( 
.A(n_957),
.B(n_937),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_955),
.B(n_956),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_955),
.A2(n_966),
.B1(n_968),
.B2(n_956),
.Y(n_1050)
);

AOI21x1_ASAP7_75t_SL g1051 ( 
.A1(n_896),
.A2(n_901),
.B(n_816),
.Y(n_1051)
);

O2A1O1Ixp5_ASAP7_75t_L g1052 ( 
.A1(n_970),
.A2(n_917),
.B(n_677),
.C(n_822),
.Y(n_1052)
);

AOI21xp33_ASAP7_75t_L g1053 ( 
.A1(n_870),
.A2(n_917),
.B(n_916),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_955),
.B(n_956),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_953),
.A2(n_967),
.B(n_960),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_937),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_865),
.B(n_928),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_962),
.B(n_955),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_965),
.B(n_962),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_957),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_934),
.A2(n_819),
.B(n_844),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_934),
.A2(n_819),
.B(n_844),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_955),
.B(n_956),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_965),
.B(n_962),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_865),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_823),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_934),
.A2(n_819),
.B(n_844),
.Y(n_1067)
);

NOR2x1_ASAP7_75t_L g1068 ( 
.A(n_957),
.B(n_937),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_934),
.A2(n_819),
.B(n_844),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_865),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_962),
.B(n_955),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_964),
.B(n_972),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_955),
.B(n_956),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_955),
.B(n_956),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_962),
.B(n_955),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_865),
.B(n_928),
.Y(n_1076)
);

AOI21xp33_ASAP7_75t_L g1077 ( 
.A1(n_870),
.A2(n_917),
.B(n_916),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_955),
.A2(n_966),
.B1(n_968),
.B2(n_956),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_934),
.A2(n_819),
.B(n_844),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_865),
.B(n_928),
.Y(n_1080)
);

AOI221xp5_ASAP7_75t_L g1081 ( 
.A1(n_954),
.A2(n_708),
.B1(n_655),
.B2(n_962),
.C(n_870),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_965),
.B(n_962),
.Y(n_1082)
);

AOI21x1_ASAP7_75t_L g1083 ( 
.A1(n_885),
.A2(n_844),
.B(n_886),
.Y(n_1083)
);

NAND2x1_ASAP7_75t_L g1084 ( 
.A(n_957),
.B(n_687),
.Y(n_1084)
);

O2A1O1Ixp5_ASAP7_75t_L g1085 ( 
.A1(n_970),
.A2(n_917),
.B(n_677),
.C(n_822),
.Y(n_1085)
);

OAI22x1_ASAP7_75t_L g1086 ( 
.A1(n_964),
.A2(n_972),
.B1(n_962),
.B2(n_916),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_953),
.A2(n_967),
.B(n_960),
.Y(n_1087)
);

OAI21xp33_ASAP7_75t_L g1088 ( 
.A1(n_962),
.A2(n_677),
.B(n_964),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_962),
.B(n_955),
.Y(n_1089)
);

OAI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_953),
.A2(n_967),
.B(n_960),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_955),
.A2(n_966),
.B1(n_968),
.B2(n_956),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_934),
.A2(n_819),
.B(n_844),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_957),
.Y(n_1093)
);

NAND3xp33_ASAP7_75t_L g1094 ( 
.A(n_964),
.B(n_972),
.C(n_970),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_955),
.B(n_956),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_965),
.B(n_962),
.Y(n_1096)
);

NOR2x1_ASAP7_75t_L g1097 ( 
.A(n_957),
.B(n_937),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_953),
.A2(n_967),
.B(n_960),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_965),
.B(n_962),
.Y(n_1099)
);

BUFx10_ASAP7_75t_L g1100 ( 
.A(n_930),
.Y(n_1100)
);

AOI21xp33_ASAP7_75t_L g1101 ( 
.A1(n_870),
.A2(n_917),
.B(n_916),
.Y(n_1101)
);

O2A1O1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_984),
.A2(n_1088),
.B(n_988),
.C(n_1101),
.Y(n_1102)
);

INVx1_ASAP7_75t_SL g1103 ( 
.A(n_996),
.Y(n_1103)
);

A2O1A1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_1053),
.A2(n_1077),
.B(n_1101),
.C(n_1081),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_1059),
.B(n_1064),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_1053),
.A2(n_1077),
.B1(n_1086),
.B2(n_980),
.Y(n_1106)
);

INVxp67_ASAP7_75t_L g1107 ( 
.A(n_996),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_1058),
.B(n_1071),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_1056),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_1075),
.B(n_1089),
.Y(n_1110)
);

OR2x2_ASAP7_75t_L g1111 ( 
.A(n_1049),
.B(n_1054),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1049),
.B(n_1054),
.Y(n_1112)
);

NAND2x1_ASAP7_75t_L g1113 ( 
.A(n_1016),
.B(n_1060),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_978),
.Y(n_1114)
);

NAND3xp33_ASAP7_75t_L g1115 ( 
.A(n_1094),
.B(n_980),
.C(n_1006),
.Y(n_1115)
);

INVx3_ASAP7_75t_SL g1116 ( 
.A(n_1010),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_1010),
.B(n_976),
.Y(n_1117)
);

BUFx2_ASAP7_75t_SL g1118 ( 
.A(n_1009),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_999),
.Y(n_1119)
);

O2A1O1Ixp5_ASAP7_75t_L g1120 ( 
.A1(n_1072),
.A2(n_1052),
.B(n_1085),
.C(n_1047),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_1009),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_1082),
.B(n_1096),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_1009),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1099),
.B(n_1017),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_979),
.B(n_1074),
.Y(n_1125)
);

INVx1_ASAP7_75t_SL g1126 ( 
.A(n_975),
.Y(n_1126)
);

OR2x2_ASAP7_75t_L g1127 ( 
.A(n_1063),
.B(n_1073),
.Y(n_1127)
);

INVx5_ASAP7_75t_L g1128 ( 
.A(n_1016),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1063),
.B(n_1073),
.Y(n_1129)
);

AOI21x1_ASAP7_75t_SL g1130 ( 
.A1(n_986),
.A2(n_994),
.B(n_1095),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_982),
.A2(n_1012),
.B(n_989),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1066),
.Y(n_1132)
);

INVx3_ASAP7_75t_SL g1133 ( 
.A(n_997),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_975),
.B(n_1057),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_1046),
.B(n_1050),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_SL g1136 ( 
.A(n_1035),
.B(n_1022),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_992),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_983),
.B(n_991),
.Y(n_1138)
);

BUFx3_ASAP7_75t_L g1139 ( 
.A(n_985),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_SL g1140 ( 
.A1(n_1055),
.A2(n_1087),
.B(n_1098),
.C(n_1090),
.Y(n_1140)
);

NAND2x1_ASAP7_75t_L g1141 ( 
.A(n_1060),
.B(n_1093),
.Y(n_1141)
);

AND2x4_ASAP7_75t_L g1142 ( 
.A(n_1057),
.B(n_1076),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1046),
.B(n_1050),
.Y(n_1143)
);

BUFx3_ASAP7_75t_L g1144 ( 
.A(n_985),
.Y(n_1144)
);

AND2x2_ASAP7_75t_SL g1145 ( 
.A(n_1045),
.B(n_986),
.Y(n_1145)
);

AOI222xp33_ASAP7_75t_L g1146 ( 
.A1(n_1078),
.A2(n_1091),
.B1(n_982),
.B2(n_1001),
.C1(n_1003),
.C2(n_994),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_985),
.Y(n_1147)
);

AND3x1_ASAP7_75t_SL g1148 ( 
.A(n_981),
.B(n_1033),
.C(n_1100),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1004),
.B(n_998),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_SL g1150 ( 
.A(n_1078),
.B(n_1091),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1008),
.B(n_995),
.Y(n_1151)
);

NAND2x1p5_ASAP7_75t_L g1152 ( 
.A(n_1093),
.B(n_1076),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_1065),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1031),
.B(n_1034),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1100),
.B(n_1080),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1080),
.B(n_1026),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_1007),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_990),
.A2(n_987),
.B(n_1000),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_1065),
.Y(n_1159)
);

INVx1_ASAP7_75t_SL g1160 ( 
.A(n_1070),
.Y(n_1160)
);

AND2x6_ASAP7_75t_L g1161 ( 
.A(n_1027),
.B(n_1048),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1055),
.A2(n_1090),
.B(n_1087),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1038),
.A2(n_1040),
.B(n_1030),
.Y(n_1163)
);

HB1xp67_ASAP7_75t_L g1164 ( 
.A(n_1070),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1068),
.B(n_1097),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1030),
.A2(n_1024),
.B(n_1020),
.Y(n_1166)
);

AOI221xp5_ASAP7_75t_L g1167 ( 
.A1(n_1028),
.A2(n_1005),
.B1(n_1018),
.B2(n_1002),
.C(n_1044),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1031),
.B(n_1034),
.Y(n_1168)
);

OAI31xp33_ASAP7_75t_L g1169 ( 
.A1(n_1018),
.A2(n_1028),
.A3(n_1015),
.B(n_1011),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_1070),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_993),
.B(n_1023),
.Y(n_1171)
);

INVxp67_ASAP7_75t_SL g1172 ( 
.A(n_1013),
.Y(n_1172)
);

INVx4_ASAP7_75t_L g1173 ( 
.A(n_1023),
.Y(n_1173)
);

AND2x2_ASAP7_75t_SL g1174 ( 
.A(n_1041),
.B(n_993),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1036),
.B(n_1029),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1041),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_993),
.B(n_1014),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1042),
.B(n_1043),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_1084),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1032),
.B(n_1037),
.Y(n_1180)
);

OAI321xp33_ASAP7_75t_L g1181 ( 
.A1(n_977),
.A2(n_1083),
.A3(n_1051),
.B1(n_1021),
.B2(n_1037),
.C(n_1019),
.Y(n_1181)
);

BUFx12f_ASAP7_75t_L g1182 ( 
.A(n_1039),
.Y(n_1182)
);

BUFx12f_ASAP7_75t_L g1183 ( 
.A(n_1039),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_1039),
.B(n_1025),
.Y(n_1184)
);

BUFx12f_ASAP7_75t_L g1185 ( 
.A(n_1019),
.Y(n_1185)
);

OAI21xp33_ASAP7_75t_L g1186 ( 
.A1(n_1061),
.A2(n_1092),
.B(n_1067),
.Y(n_1186)
);

OR2x2_ASAP7_75t_L g1187 ( 
.A(n_1062),
.B(n_1069),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1079),
.B(n_1059),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1058),
.B(n_955),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1058),
.B(n_955),
.Y(n_1190)
);

NAND2x1p5_ASAP7_75t_L g1191 ( 
.A(n_1016),
.B(n_957),
.Y(n_1191)
);

INVx3_ASAP7_75t_SL g1192 ( 
.A(n_1010),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_1056),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1049),
.A2(n_955),
.B1(n_966),
.B2(n_956),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1088),
.B(n_964),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_975),
.B(n_1057),
.Y(n_1196)
);

NAND2x1p5_ASAP7_75t_L g1197 ( 
.A(n_1016),
.B(n_957),
.Y(n_1197)
);

OR2x2_ASAP7_75t_L g1198 ( 
.A(n_1049),
.B(n_1054),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_975),
.B(n_1057),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_978),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_975),
.B(n_1057),
.Y(n_1201)
);

INVx1_ASAP7_75t_SL g1202 ( 
.A(n_996),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_978),
.Y(n_1203)
);

A2O1A1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_1088),
.A2(n_970),
.B(n_916),
.C(n_964),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_1009),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1058),
.B(n_955),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1049),
.A2(n_955),
.B1(n_966),
.B2(n_956),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1058),
.B(n_955),
.Y(n_1208)
);

INVx1_ASAP7_75t_SL g1209 ( 
.A(n_996),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1049),
.A2(n_955),
.B1(n_966),
.B2(n_956),
.Y(n_1210)
);

BUFx8_ASAP7_75t_L g1211 ( 
.A(n_1007),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_978),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1056),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_1009),
.Y(n_1214)
);

INVx2_ASAP7_75t_SL g1215 ( 
.A(n_1056),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_1056),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_978),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_1009),
.Y(n_1218)
);

INVx2_ASAP7_75t_SL g1219 ( 
.A(n_1056),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_1056),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1059),
.B(n_1064),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_1007),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1058),
.B(n_955),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_L g1224 ( 
.A(n_1009),
.Y(n_1224)
);

O2A1O1Ixp5_ASAP7_75t_L g1225 ( 
.A1(n_988),
.A2(n_970),
.B(n_677),
.C(n_917),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_1009),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_996),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_978),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_975),
.B(n_1057),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_978),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1058),
.B(n_955),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_984),
.A2(n_970),
.B(n_1088),
.C(n_962),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_1009),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1009),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1114),
.Y(n_1235)
);

INVx4_ASAP7_75t_L g1236 ( 
.A(n_1121),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1132),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1112),
.B(n_1129),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1108),
.A2(n_1110),
.B1(n_1115),
.B2(n_1195),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1143),
.Y(n_1240)
);

OR2x6_ASAP7_75t_L g1241 ( 
.A(n_1131),
.B(n_1162),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_1220),
.Y(n_1242)
);

OR2x6_ASAP7_75t_L g1243 ( 
.A(n_1131),
.B(n_1162),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1189),
.B(n_1190),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1200),
.Y(n_1245)
);

INVxp67_ASAP7_75t_L g1246 ( 
.A(n_1227),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1143),
.Y(n_1247)
);

OAI22xp33_ASAP7_75t_SL g1248 ( 
.A1(n_1150),
.A2(n_1135),
.B1(n_1136),
.B2(n_1190),
.Y(n_1248)
);

OA21x2_ASAP7_75t_L g1249 ( 
.A1(n_1163),
.A2(n_1120),
.B(n_1158),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1203),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_1211),
.Y(n_1251)
);

INVx6_ASAP7_75t_L g1252 ( 
.A(n_1128),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1189),
.A2(n_1231),
.B1(n_1206),
.B2(n_1223),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1174),
.Y(n_1254)
);

INVx6_ASAP7_75t_L g1255 ( 
.A(n_1128),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1230),
.Y(n_1256)
);

OA21x2_ASAP7_75t_L g1257 ( 
.A1(n_1163),
.A2(n_1158),
.B(n_1166),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1119),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1178),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1188),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_1185),
.Y(n_1261)
);

INVx6_ASAP7_75t_L g1262 ( 
.A(n_1128),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1182),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1151),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_1103),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1112),
.B(n_1129),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1151),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1206),
.A2(n_1223),
.B1(n_1231),
.B2(n_1208),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1212),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1217),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1171),
.B(n_1134),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1109),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1208),
.A2(n_1127),
.B1(n_1198),
.B2(n_1111),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1194),
.A2(n_1207),
.B1(n_1210),
.B2(n_1106),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1228),
.Y(n_1275)
);

BUFx3_ASAP7_75t_L g1276 ( 
.A(n_1213),
.Y(n_1276)
);

BUFx8_ASAP7_75t_SL g1277 ( 
.A(n_1157),
.Y(n_1277)
);

OAI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1136),
.A2(n_1150),
.B1(n_1192),
.B2(n_1116),
.Y(n_1278)
);

CKINVDCx8_ASAP7_75t_R g1279 ( 
.A(n_1118),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1134),
.B(n_1142),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1202),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1137),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1194),
.B(n_1207),
.Y(n_1283)
);

BUFx4f_ASAP7_75t_SL g1284 ( 
.A(n_1211),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_SL g1285 ( 
.A1(n_1138),
.A2(n_1145),
.B1(n_1210),
.B2(n_1172),
.Y(n_1285)
);

BUFx12f_ASAP7_75t_L g1286 ( 
.A(n_1222),
.Y(n_1286)
);

AOI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1180),
.A2(n_1184),
.B(n_1154),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1175),
.Y(n_1288)
);

BUFx12f_ASAP7_75t_L g1289 ( 
.A(n_1121),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1175),
.Y(n_1290)
);

BUFx3_ASAP7_75t_L g1291 ( 
.A(n_1216),
.Y(n_1291)
);

OA21x2_ASAP7_75t_L g1292 ( 
.A1(n_1181),
.A2(n_1186),
.B(n_1104),
.Y(n_1292)
);

INVxp67_ASAP7_75t_L g1293 ( 
.A(n_1202),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1117),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1183),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1234),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1146),
.A2(n_1167),
.B1(n_1105),
.B2(n_1221),
.Y(n_1297)
);

OA21x2_ASAP7_75t_L g1298 ( 
.A1(n_1181),
.A2(n_1225),
.B(n_1167),
.Y(n_1298)
);

AOI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1122),
.A2(n_1125),
.B1(n_1124),
.B2(n_1156),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1107),
.B(n_1209),
.Y(n_1300)
);

INVx2_ASAP7_75t_SL g1301 ( 
.A(n_1139),
.Y(n_1301)
);

CKINVDCx6p67_ASAP7_75t_R g1302 ( 
.A(n_1133),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1187),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1204),
.A2(n_1209),
.B1(n_1126),
.B2(n_1149),
.Y(n_1304)
);

INVx2_ASAP7_75t_SL g1305 ( 
.A(n_1144),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_SL g1306 ( 
.A1(n_1155),
.A2(n_1215),
.B1(n_1193),
.B2(n_1219),
.Y(n_1306)
);

BUFx2_ASAP7_75t_L g1307 ( 
.A(n_1126),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1168),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1102),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1191),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1146),
.A2(n_1169),
.B1(n_1161),
.B2(n_1201),
.Y(n_1311)
);

INVx4_ASAP7_75t_L g1312 ( 
.A(n_1121),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1232),
.A2(n_1152),
.B1(n_1199),
.B2(n_1201),
.Y(n_1313)
);

AO21x2_ASAP7_75t_L g1314 ( 
.A1(n_1140),
.A2(n_1176),
.B(n_1130),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1142),
.B(n_1199),
.Y(n_1315)
);

INVx8_ASAP7_75t_L g1316 ( 
.A(n_1196),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1161),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1153),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1113),
.A2(n_1141),
.B(n_1197),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1161),
.A2(n_1229),
.B1(n_1196),
.B2(n_1177),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1164),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_1170),
.Y(n_1322)
);

OR2x2_ASAP7_75t_L g1323 ( 
.A(n_1229),
.B(n_1152),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1147),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1161),
.Y(n_1325)
);

BUFx8_ASAP7_75t_L g1326 ( 
.A(n_1123),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1165),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1123),
.A2(n_1234),
.B1(n_1205),
.B2(n_1214),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1160),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1179),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1173),
.Y(n_1331)
);

BUFx2_ASAP7_75t_SL g1332 ( 
.A(n_1123),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1159),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1205),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1205),
.Y(n_1335)
);

BUFx2_ASAP7_75t_R g1336 ( 
.A(n_1148),
.Y(n_1336)
);

OAI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1214),
.A2(n_1218),
.B(n_1224),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1214),
.A2(n_1218),
.B1(n_1224),
.B2(n_1226),
.Y(n_1338)
);

BUFx2_ASAP7_75t_SL g1339 ( 
.A(n_1226),
.Y(n_1339)
);

INVxp67_ASAP7_75t_L g1340 ( 
.A(n_1226),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1233),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1233),
.Y(n_1342)
);

AOI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1233),
.A2(n_677),
.B1(n_1110),
.B2(n_1108),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1227),
.Y(n_1344)
);

AO21x1_ASAP7_75t_L g1345 ( 
.A1(n_1274),
.A2(n_1283),
.B(n_1248),
.Y(n_1345)
);

BUFx2_ASAP7_75t_SL g1346 ( 
.A(n_1279),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1344),
.Y(n_1347)
);

AO21x1_ASAP7_75t_SL g1348 ( 
.A1(n_1311),
.A2(n_1325),
.B(n_1317),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1239),
.A2(n_1343),
.B(n_1268),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1264),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1267),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1267),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1254),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1260),
.B(n_1241),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1303),
.Y(n_1355)
);

INVx4_ASAP7_75t_L g1356 ( 
.A(n_1252),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1241),
.B(n_1243),
.Y(n_1357)
);

INVx1_ASAP7_75t_SL g1358 ( 
.A(n_1272),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1287),
.Y(n_1359)
);

AND2x4_ASAP7_75t_L g1360 ( 
.A(n_1259),
.B(n_1317),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1287),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1241),
.Y(n_1362)
);

AND2x4_ASAP7_75t_L g1363 ( 
.A(n_1259),
.B(n_1325),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1243),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1243),
.B(n_1238),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1238),
.B(n_1266),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1243),
.B(n_1266),
.Y(n_1367)
);

INVx2_ASAP7_75t_SL g1368 ( 
.A(n_1344),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1308),
.B(n_1240),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1247),
.B(n_1258),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1273),
.B(n_1253),
.Y(n_1371)
);

BUFx3_ASAP7_75t_L g1372 ( 
.A(n_1254),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1315),
.B(n_1299),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1278),
.B(n_1285),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1269),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1270),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1270),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_SL g1378 ( 
.A1(n_1309),
.A2(n_1254),
.B(n_1313),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1314),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1244),
.B(n_1288),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_L g1381 ( 
.A(n_1272),
.B(n_1276),
.Y(n_1381)
);

BUFx3_ASAP7_75t_L g1382 ( 
.A(n_1254),
.Y(n_1382)
);

INVxp67_ASAP7_75t_SL g1383 ( 
.A(n_1265),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1275),
.Y(n_1384)
);

OA21x2_ASAP7_75t_L g1385 ( 
.A1(n_1290),
.A2(n_1297),
.B(n_1327),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1292),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1249),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1327),
.B(n_1237),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1276),
.B(n_1291),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1257),
.B(n_1304),
.Y(n_1390)
);

INVx2_ASAP7_75t_SL g1391 ( 
.A(n_1252),
.Y(n_1391)
);

NAND2x1_ASAP7_75t_L g1392 ( 
.A(n_1255),
.B(n_1262),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1281),
.Y(n_1393)
);

INVx2_ASAP7_75t_SL g1394 ( 
.A(n_1255),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1245),
.Y(n_1395)
);

OR2x6_ASAP7_75t_L g1396 ( 
.A(n_1263),
.B(n_1295),
.Y(n_1396)
);

BUFx6f_ASAP7_75t_L g1397 ( 
.A(n_1319),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1371),
.B(n_1298),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1354),
.B(n_1257),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1387),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1387),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1354),
.B(n_1257),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1365),
.B(n_1298),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1369),
.B(n_1294),
.Y(n_1404)
);

AND2x4_ASAP7_75t_L g1405 ( 
.A(n_1362),
.B(n_1263),
.Y(n_1405)
);

INVxp67_ASAP7_75t_SL g1406 ( 
.A(n_1359),
.Y(n_1406)
);

INVx4_ASAP7_75t_L g1407 ( 
.A(n_1356),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1365),
.B(n_1261),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1396),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1396),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1390),
.B(n_1261),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1359),
.Y(n_1412)
);

NOR2x1_ASAP7_75t_L g1413 ( 
.A(n_1378),
.B(n_1295),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1390),
.B(n_1307),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1367),
.B(n_1235),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1367),
.B(n_1250),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1362),
.B(n_1307),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1349),
.A2(n_1246),
.B1(n_1300),
.B2(n_1280),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1357),
.B(n_1256),
.Y(n_1419)
);

OAI21xp33_ASAP7_75t_L g1420 ( 
.A1(n_1374),
.A2(n_1293),
.B(n_1306),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1357),
.B(n_1329),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1364),
.B(n_1329),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_1360),
.B(n_1310),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1396),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1369),
.B(n_1282),
.Y(n_1425)
);

OAI33xp33_ASAP7_75t_L g1426 ( 
.A1(n_1380),
.A2(n_1321),
.A3(n_1330),
.B1(n_1334),
.B2(n_1335),
.B3(n_1341),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1397),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1361),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1361),
.B(n_1318),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1386),
.B(n_1291),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1345),
.B(n_1330),
.Y(n_1431)
);

OAI221xp5_ASAP7_75t_L g1432 ( 
.A1(n_1373),
.A2(n_1320),
.B1(n_1279),
.B2(n_1322),
.C(n_1323),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1415),
.B(n_1383),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1403),
.B(n_1379),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1403),
.B(n_1379),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1400),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1415),
.B(n_1347),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_L g1438 ( 
.A(n_1420),
.B(n_1381),
.Y(n_1438)
);

OAI21xp33_ASAP7_75t_L g1439 ( 
.A1(n_1420),
.A2(n_1378),
.B(n_1366),
.Y(n_1439)
);

NAND3xp33_ASAP7_75t_L g1440 ( 
.A(n_1431),
.B(n_1393),
.C(n_1368),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_SL g1441 ( 
.A1(n_1418),
.A2(n_1280),
.B(n_1389),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_SL g1442 ( 
.A(n_1413),
.B(n_1345),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1416),
.B(n_1419),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_SL g1444 ( 
.A(n_1413),
.B(n_1284),
.Y(n_1444)
);

AOI211xp5_ASAP7_75t_L g1445 ( 
.A1(n_1432),
.A2(n_1431),
.B(n_1398),
.C(n_1426),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1416),
.B(n_1368),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1416),
.B(n_1384),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1404),
.B(n_1358),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1404),
.B(n_1408),
.Y(n_1449)
);

OAI221xp5_ASAP7_75t_SL g1450 ( 
.A1(n_1418),
.A2(n_1396),
.B1(n_1338),
.B2(n_1302),
.C(n_1323),
.Y(n_1450)
);

AOI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1432),
.A2(n_1385),
.B1(n_1396),
.B2(n_1346),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1419),
.B(n_1370),
.Y(n_1452)
);

OAI21xp5_ASAP7_75t_SL g1453 ( 
.A1(n_1398),
.A2(n_1280),
.B(n_1271),
.Y(n_1453)
);

OAI21xp5_ASAP7_75t_SL g1454 ( 
.A1(n_1408),
.A2(n_1271),
.B(n_1328),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1421),
.B(n_1408),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1405),
.A2(n_1348),
.B1(n_1385),
.B2(n_1382),
.Y(n_1456)
);

OAI21xp5_ASAP7_75t_SL g1457 ( 
.A1(n_1405),
.A2(n_1271),
.B(n_1337),
.Y(n_1457)
);

OAI221xp5_ASAP7_75t_L g1458 ( 
.A1(n_1411),
.A2(n_1346),
.B1(n_1392),
.B2(n_1242),
.C(n_1394),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1399),
.B(n_1360),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_SL g1460 ( 
.A1(n_1409),
.A2(n_1382),
.B1(n_1372),
.B2(n_1353),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_SL g1461 ( 
.A1(n_1409),
.A2(n_1382),
.B1(n_1372),
.B2(n_1353),
.Y(n_1461)
);

NAND3xp33_ASAP7_75t_L g1462 ( 
.A(n_1429),
.B(n_1385),
.C(n_1388),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1422),
.B(n_1355),
.Y(n_1463)
);

AOI221xp5_ASAP7_75t_L g1464 ( 
.A1(n_1426),
.A2(n_1388),
.B1(n_1350),
.B2(n_1351),
.C(n_1352),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1399),
.B(n_1360),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1402),
.B(n_1363),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1422),
.B(n_1355),
.Y(n_1467)
);

OAI221xp5_ASAP7_75t_L g1468 ( 
.A1(n_1411),
.A2(n_1392),
.B1(n_1242),
.B2(n_1394),
.C(n_1391),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1422),
.B(n_1375),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_SL g1470 ( 
.A(n_1407),
.B(n_1251),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1425),
.B(n_1375),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_SL g1472 ( 
.A(n_1405),
.B(n_1356),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1425),
.B(n_1376),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1423),
.B(n_1376),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1423),
.B(n_1377),
.Y(n_1475)
);

NAND3xp33_ASAP7_75t_L g1476 ( 
.A(n_1429),
.B(n_1385),
.C(n_1395),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1443),
.B(n_1414),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1459),
.B(n_1402),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1438),
.B(n_1302),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1459),
.B(n_1465),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1436),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1437),
.B(n_1414),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1436),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1434),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1465),
.B(n_1466),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1434),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1435),
.B(n_1414),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1435),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1449),
.B(n_1412),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1469),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1466),
.B(n_1402),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1455),
.B(n_1405),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1474),
.B(n_1411),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1463),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1455),
.B(n_1400),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1467),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1440),
.B(n_1412),
.Y(n_1497)
);

INVxp67_ASAP7_75t_L g1498 ( 
.A(n_1440),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1447),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1475),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1462),
.B(n_1427),
.Y(n_1501)
);

INVxp67_ASAP7_75t_L g1502 ( 
.A(n_1442),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1471),
.B(n_1428),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1473),
.B(n_1428),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1445),
.B(n_1406),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1448),
.B(n_1423),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1462),
.B(n_1427),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1452),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1445),
.B(n_1406),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1456),
.B(n_1401),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1446),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1501),
.B(n_1409),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1488),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1483),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1484),
.B(n_1410),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1497),
.B(n_1433),
.Y(n_1516)
);

OAI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1505),
.A2(n_1451),
.B1(n_1444),
.B2(n_1470),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_1505),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1484),
.B(n_1410),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1498),
.B(n_1476),
.Y(n_1520)
);

INVx2_ASAP7_75t_SL g1521 ( 
.A(n_1501),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1483),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_R g1523 ( 
.A(n_1479),
.B(n_1251),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1486),
.B(n_1410),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1488),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1481),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1498),
.B(n_1476),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1483),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1481),
.Y(n_1529)
);

INVxp67_ASAP7_75t_SL g1530 ( 
.A(n_1497),
.Y(n_1530)
);

OAI21xp33_ASAP7_75t_L g1531 ( 
.A1(n_1509),
.A2(n_1439),
.B(n_1502),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1486),
.B(n_1410),
.Y(n_1532)
);

AND2x2_ASAP7_75t_SL g1533 ( 
.A(n_1509),
.B(n_1451),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1502),
.B(n_1464),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1487),
.B(n_1430),
.Y(n_1535)
);

NOR3xp33_ASAP7_75t_SL g1536 ( 
.A(n_1489),
.B(n_1439),
.C(n_1450),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1478),
.B(n_1424),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1487),
.B(n_1430),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1478),
.B(n_1424),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1495),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1493),
.B(n_1430),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1493),
.B(n_1417),
.Y(n_1542)
);

INVxp67_ASAP7_75t_SL g1543 ( 
.A(n_1503),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1477),
.B(n_1417),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1495),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1510),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1491),
.B(n_1424),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1501),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1495),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1491),
.B(n_1424),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1500),
.Y(n_1551)
);

NOR2x1p5_ASAP7_75t_L g1552 ( 
.A(n_1518),
.B(n_1286),
.Y(n_1552)
);

AOI21xp33_ASAP7_75t_L g1553 ( 
.A1(n_1517),
.A2(n_1468),
.B(n_1458),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1551),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1546),
.B(n_1480),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1551),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1531),
.B(n_1534),
.Y(n_1557)
);

NOR2x1_ASAP7_75t_L g1558 ( 
.A(n_1518),
.B(n_1520),
.Y(n_1558)
);

INVx1_ASAP7_75t_SL g1559 ( 
.A(n_1523),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1513),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1546),
.B(n_1480),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1531),
.B(n_1534),
.Y(n_1562)
);

NAND2x1_ASAP7_75t_SL g1563 ( 
.A(n_1512),
.B(n_1501),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1518),
.B(n_1499),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1513),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1520),
.B(n_1482),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1512),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1525),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1514),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1533),
.A2(n_1441),
.B1(n_1453),
.B2(n_1461),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1512),
.B(n_1521),
.Y(n_1571)
);

NAND3xp33_ASAP7_75t_SL g1572 ( 
.A(n_1527),
.B(n_1441),
.C(n_1460),
.Y(n_1572)
);

AOI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1533),
.A2(n_1472),
.B(n_1453),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1536),
.B(n_1499),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1512),
.B(n_1485),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1525),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1536),
.B(n_1500),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1516),
.B(n_1286),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1533),
.B(n_1511),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1527),
.B(n_1482),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1521),
.B(n_1515),
.Y(n_1581)
);

AOI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1530),
.A2(n_1457),
.B(n_1503),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1521),
.B(n_1507),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1515),
.B(n_1485),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1535),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1535),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1544),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1543),
.B(n_1477),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1519),
.B(n_1492),
.Y(n_1589)
);

AOI221xp5_ASAP7_75t_L g1590 ( 
.A1(n_1530),
.A2(n_1511),
.B1(n_1507),
.B2(n_1510),
.C(n_1508),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1548),
.B(n_1507),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1514),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1516),
.B(n_1490),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1519),
.B(n_1492),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1554),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1556),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1575),
.B(n_1543),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1566),
.B(n_1544),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1558),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1566),
.B(n_1541),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1560),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_L g1602 ( 
.A(n_1559),
.B(n_1541),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1580),
.B(n_1538),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1575),
.B(n_1548),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1560),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1574),
.B(n_1524),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1580),
.B(n_1579),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1565),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1563),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1557),
.A2(n_1507),
.B1(n_1510),
.B2(n_1348),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1565),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1562),
.A2(n_1548),
.B1(n_1532),
.B2(n_1524),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1571),
.B(n_1532),
.Y(n_1613)
);

NOR2x1_ASAP7_75t_L g1614 ( 
.A(n_1552),
.B(n_1526),
.Y(n_1614)
);

INVx1_ASAP7_75t_SL g1615 ( 
.A(n_1563),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1578),
.B(n_1542),
.Y(n_1616)
);

INVx3_ASAP7_75t_L g1617 ( 
.A(n_1583),
.Y(n_1617)
);

INVx1_ASAP7_75t_SL g1618 ( 
.A(n_1571),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1568),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1568),
.Y(n_1620)
);

AND3x2_ASAP7_75t_L g1621 ( 
.A(n_1581),
.B(n_1529),
.C(n_1526),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1576),
.Y(n_1622)
);

INVx1_ASAP7_75t_SL g1623 ( 
.A(n_1581),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1576),
.Y(n_1624)
);

INVxp67_ASAP7_75t_SL g1625 ( 
.A(n_1567),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1564),
.B(n_1538),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1555),
.B(n_1529),
.Y(n_1627)
);

OAI221xp5_ASAP7_75t_L g1628 ( 
.A1(n_1553),
.A2(n_1457),
.B1(n_1454),
.B2(n_1489),
.C(n_1504),
.Y(n_1628)
);

NOR2x1p5_ASAP7_75t_L g1629 ( 
.A(n_1572),
.B(n_1542),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1577),
.B(n_1540),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1617),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1623),
.Y(n_1632)
);

AOI221xp5_ASAP7_75t_L g1633 ( 
.A1(n_1599),
.A2(n_1602),
.B1(n_1606),
.B2(n_1628),
.C(n_1590),
.Y(n_1633)
);

INVx1_ASAP7_75t_SL g1634 ( 
.A(n_1609),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1601),
.Y(n_1635)
);

OAI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1629),
.A2(n_1570),
.B1(n_1573),
.B2(n_1582),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_L g1637 ( 
.A(n_1602),
.B(n_1277),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1618),
.B(n_1584),
.Y(n_1638)
);

O2A1O1Ixp33_ASAP7_75t_L g1639 ( 
.A1(n_1615),
.A2(n_1588),
.B(n_1593),
.C(n_1587),
.Y(n_1639)
);

AOI211xp5_ASAP7_75t_SL g1640 ( 
.A1(n_1625),
.A2(n_1567),
.B(n_1583),
.C(n_1588),
.Y(n_1640)
);

OR3x1_ASAP7_75t_L g1641 ( 
.A(n_1616),
.B(n_1586),
.C(n_1585),
.Y(n_1641)
);

OAI21xp33_ASAP7_75t_SL g1642 ( 
.A1(n_1614),
.A2(n_1561),
.B(n_1555),
.Y(n_1642)
);

A2O1A1Ixp33_ASAP7_75t_L g1643 ( 
.A1(n_1610),
.A2(n_1561),
.B(n_1583),
.C(n_1567),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1607),
.B(n_1616),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1605),
.Y(n_1645)
);

INVx2_ASAP7_75t_SL g1646 ( 
.A(n_1617),
.Y(n_1646)
);

AOI221xp5_ASAP7_75t_L g1647 ( 
.A1(n_1610),
.A2(n_1586),
.B1(n_1585),
.B2(n_1569),
.C(n_1592),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1617),
.B(n_1584),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1597),
.B(n_1589),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1608),
.Y(n_1650)
);

INVx2_ASAP7_75t_SL g1651 ( 
.A(n_1621),
.Y(n_1651)
);

OAI22xp33_ASAP7_75t_SL g1652 ( 
.A1(n_1630),
.A2(n_1591),
.B1(n_1540),
.B2(n_1545),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1611),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1613),
.Y(n_1654)
);

A2O1A1Ixp33_ASAP7_75t_SL g1655 ( 
.A1(n_1612),
.A2(n_1569),
.B(n_1592),
.C(n_1528),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_SL g1656 ( 
.A(n_1597),
.B(n_1336),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1635),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1645),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1634),
.B(n_1613),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1651),
.B(n_1627),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1648),
.Y(n_1661)
);

OAI21xp5_ASAP7_75t_SL g1662 ( 
.A1(n_1636),
.A2(n_1612),
.B(n_1604),
.Y(n_1662)
);

INVx1_ASAP7_75t_SL g1663 ( 
.A(n_1632),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_SL g1664 ( 
.A(n_1633),
.B(n_1627),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1644),
.B(n_1633),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1648),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1646),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1631),
.B(n_1627),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1650),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1653),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1641),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1644),
.B(n_1604),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1649),
.B(n_1598),
.Y(n_1673)
);

NOR2x1_ASAP7_75t_L g1674 ( 
.A(n_1637),
.B(n_1619),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1654),
.B(n_1595),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1640),
.B(n_1596),
.Y(n_1676)
);

OA22x2_ASAP7_75t_L g1677 ( 
.A1(n_1671),
.A2(n_1638),
.B1(n_1620),
.B2(n_1622),
.Y(n_1677)
);

AOI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1665),
.A2(n_1639),
.B(n_1655),
.Y(n_1678)
);

OAI221xp5_ASAP7_75t_L g1679 ( 
.A1(n_1662),
.A2(n_1642),
.B1(n_1647),
.B2(n_1643),
.C(n_1639),
.Y(n_1679)
);

NOR3xp33_ASAP7_75t_L g1680 ( 
.A(n_1663),
.B(n_1647),
.C(n_1652),
.Y(n_1680)
);

OAI211xp5_ASAP7_75t_L g1681 ( 
.A1(n_1664),
.A2(n_1671),
.B(n_1676),
.C(n_1674),
.Y(n_1681)
);

AOI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1664),
.A2(n_1656),
.B(n_1624),
.Y(n_1682)
);

OAI21xp33_ASAP7_75t_L g1683 ( 
.A1(n_1659),
.A2(n_1660),
.B(n_1672),
.Y(n_1683)
);

AOI222xp33_ASAP7_75t_L g1684 ( 
.A1(n_1657),
.A2(n_1591),
.B1(n_1589),
.B2(n_1594),
.C1(n_1545),
.C2(n_1549),
.Y(n_1684)
);

OAI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1660),
.A2(n_1626),
.B(n_1600),
.Y(n_1685)
);

AOI211xp5_ASAP7_75t_L g1686 ( 
.A1(n_1661),
.A2(n_1603),
.B(n_1626),
.C(n_1591),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1661),
.B(n_1594),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1666),
.B(n_1603),
.Y(n_1688)
);

NAND2x1_ASAP7_75t_SL g1689 ( 
.A(n_1677),
.B(n_1668),
.Y(n_1689)
);

OA211x2_ASAP7_75t_L g1690 ( 
.A1(n_1683),
.A2(n_1675),
.B(n_1667),
.C(n_1666),
.Y(n_1690)
);

AND5x1_ASAP7_75t_L g1691 ( 
.A(n_1686),
.B(n_1673),
.C(n_1668),
.D(n_1667),
.E(n_1670),
.Y(n_1691)
);

NAND5xp2_ASAP7_75t_L g1692 ( 
.A(n_1679),
.B(n_1669),
.C(n_1658),
.D(n_1673),
.E(n_1668),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_SL g1693 ( 
.A(n_1678),
.B(n_1514),
.Y(n_1693)
);

NOR2xp67_ASAP7_75t_L g1694 ( 
.A(n_1681),
.B(n_1522),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1688),
.Y(n_1695)
);

NAND3xp33_ASAP7_75t_L g1696 ( 
.A(n_1680),
.B(n_1326),
.C(n_1324),
.Y(n_1696)
);

NAND4xp25_ASAP7_75t_L g1697 ( 
.A(n_1682),
.B(n_1454),
.C(n_1506),
.D(n_1324),
.Y(n_1697)
);

AOI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1687),
.A2(n_1522),
.B1(n_1528),
.B2(n_1549),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_L g1699 ( 
.A(n_1685),
.B(n_1277),
.Y(n_1699)
);

AOI221xp5_ASAP7_75t_L g1700 ( 
.A1(n_1692),
.A2(n_1684),
.B1(n_1522),
.B2(n_1528),
.C(n_1504),
.Y(n_1700)
);

NAND4xp25_ASAP7_75t_L g1701 ( 
.A(n_1696),
.B(n_1550),
.C(n_1547),
.D(n_1539),
.Y(n_1701)
);

NOR3x1_ASAP7_75t_L g1702 ( 
.A(n_1695),
.B(n_1305),
.C(n_1301),
.Y(n_1702)
);

NOR3xp33_ASAP7_75t_L g1703 ( 
.A(n_1699),
.B(n_1305),
.C(n_1301),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1689),
.Y(n_1704)
);

A2O1A1Ixp33_ASAP7_75t_L g1705 ( 
.A1(n_1694),
.A2(n_1550),
.B(n_1547),
.C(n_1539),
.Y(n_1705)
);

AOI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1704),
.A2(n_1690),
.B1(n_1697),
.B2(n_1693),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1702),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1701),
.Y(n_1708)
);

INVxp67_ASAP7_75t_L g1709 ( 
.A(n_1703),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1705),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1700),
.Y(n_1711)
);

AND4x1_ASAP7_75t_L g1712 ( 
.A(n_1706),
.B(n_1691),
.C(n_1698),
.D(n_1326),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1707),
.B(n_1537),
.Y(n_1713)
);

NAND3x1_ASAP7_75t_SL g1714 ( 
.A(n_1709),
.B(n_1326),
.C(n_1289),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1710),
.B(n_1537),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1708),
.B(n_1490),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1715),
.Y(n_1717)
);

XNOR2xp5_ASAP7_75t_L g1718 ( 
.A(n_1712),
.B(n_1714),
.Y(n_1718)
);

OAI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1716),
.A2(n_1711),
.B1(n_1709),
.B2(n_1289),
.Y(n_1719)
);

AO22x1_ASAP7_75t_L g1720 ( 
.A1(n_1717),
.A2(n_1713),
.B1(n_1296),
.B2(n_1236),
.Y(n_1720)
);

NOR3xp33_ASAP7_75t_L g1721 ( 
.A(n_1720),
.B(n_1719),
.C(n_1718),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1721),
.B(n_1508),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1721),
.Y(n_1723)
);

OAI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1723),
.A2(n_1340),
.B1(n_1494),
.B2(n_1496),
.Y(n_1724)
);

OAI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1722),
.A2(n_1333),
.B(n_1494),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1724),
.B(n_1496),
.Y(n_1726)
);

OAI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1725),
.A2(n_1333),
.B(n_1312),
.Y(n_1727)
);

AOI22x1_ASAP7_75t_L g1728 ( 
.A1(n_1726),
.A2(n_1236),
.B1(n_1312),
.B2(n_1339),
.Y(n_1728)
);

OAI221xp5_ASAP7_75t_R g1729 ( 
.A1(n_1728),
.A2(n_1727),
.B1(n_1316),
.B2(n_1332),
.C(n_1339),
.Y(n_1729)
);

OAI221xp5_ASAP7_75t_R g1730 ( 
.A1(n_1729),
.A2(n_1316),
.B1(n_1332),
.B2(n_1296),
.C(n_1312),
.Y(n_1730)
);

AOI211xp5_ASAP7_75t_L g1731 ( 
.A1(n_1730),
.A2(n_1334),
.B(n_1331),
.C(n_1342),
.Y(n_1731)
);


endmodule