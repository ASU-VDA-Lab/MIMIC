module fake_netlist_6_2271_n_1270 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1270);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1270;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_188;
wire n_509;
wire n_245;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_873;
wire n_461;
wire n_383;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_713;
wire n_976;
wire n_224;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_277;
wire n_618;
wire n_199;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_210;
wire n_1069;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_1052;
wire n_462;
wire n_1033;
wire n_304;
wire n_694;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_615;
wire n_1249;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_797;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1035;
wire n_294;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_272;
wire n_526;
wire n_1183;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_184;
wire n_552;
wire n_216;
wire n_912;
wire n_745;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_474;
wire n_312;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_819;
wire n_767;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_211;
wire n_231;
wire n_505;
wire n_319;
wire n_537;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1267;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_259;
wire n_385;
wire n_858;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_238;
wire n_1095;
wire n_202;
wire n_597;
wire n_280;
wire n_1187;
wire n_610;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_183;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_302;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_239;
wire n_782;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_258;
wire n_456;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_548;
wire n_282;
wire n_833;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_273;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1241;
wire n_569;
wire n_737;
wire n_1235;
wire n_1229;
wire n_306;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_299;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_1098;
wire n_391;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_855;
wire n_591;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_969;
wire n_988;
wire n_1065;
wire n_1255;
wire n_568;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_214;
wire n_246;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1147;
wire n_763;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1205;
wire n_1258;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_911;
wire n_653;
wire n_236;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_802;
wire n_561;
wire n_980;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_257;
wire n_730;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_412;
wire n_640;
wire n_965;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_167),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_106),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_110),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_23),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_143),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_31),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_104),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_81),
.Y(n_188)
);

BUFx10_ASAP7_75t_L g189 ( 
.A(n_112),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_105),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_133),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_37),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_152),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_2),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_109),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_116),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_28),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_139),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_61),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_127),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_140),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_76),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_78),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_43),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_154),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_118),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_124),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_119),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_136),
.Y(n_210)
);

INVxp67_ASAP7_75t_SL g211 ( 
.A(n_30),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_51),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_155),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_44),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_54),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_95),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_157),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_120),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_89),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_174),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_169),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_27),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_13),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_159),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_80),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_35),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_111),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_100),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_6),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_117),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_131),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_62),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_53),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_1),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_60),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_141),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_223),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_183),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_183),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_229),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_186),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_186),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_179),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_180),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_192),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_202),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_193),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_195),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_202),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_196),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_198),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_181),
.Y(n_252)
);

BUFx10_ASAP7_75t_L g253 ( 
.A(n_194),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_234),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_182),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_200),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_184),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_205),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_234),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_222),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_231),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_231),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_190),
.Y(n_263)
);

BUFx8_ASAP7_75t_SL g264 ( 
.A(n_214),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_188),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_185),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_263),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_260),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_263),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_260),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_243),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_244),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_261),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_266),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_253),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_263),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_262),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_245),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_266),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_247),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_248),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_240),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_250),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_252),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_251),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_255),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_256),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_258),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_264),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_257),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_237),
.Y(n_293)
);

NOR2xp67_ASAP7_75t_L g294 ( 
.A(n_238),
.B(n_219),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_265),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_238),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_246),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_249),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_241),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_253),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_241),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_239),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_242),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_242),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_254),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_254),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_253),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_259),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_259),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_260),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_260),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_261),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_263),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_243),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_243),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_238),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_243),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_243),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_298),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_273),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_271),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_272),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_278),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_276),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_298),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_293),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_277),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_316),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_280),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_316),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_285),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_299),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_286),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_286),
.Y(n_334)
);

INVxp33_ASAP7_75t_SL g335 ( 
.A(n_287),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_292),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_292),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_295),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_267),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_295),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_289),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_276),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_288),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_288),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_283),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_281),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_290),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_267),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_281),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_282),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_314),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_282),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_297),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_276),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_296),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_297),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_315),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_317),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_318),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_284),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_284),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_269),
.Y(n_362)
);

INVxp33_ASAP7_75t_L g363 ( 
.A(n_305),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_269),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_291),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_306),
.Y(n_366)
);

BUFx8_ASAP7_75t_SL g367 ( 
.A(n_327),
.Y(n_367)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_339),
.Y(n_368)
);

BUFx12f_ASAP7_75t_L g369 ( 
.A(n_321),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_348),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_343),
.Y(n_371)
);

CKINVDCx11_ASAP7_75t_R g372 ( 
.A(n_345),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_328),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_333),
.B(n_309),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_348),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_333),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_334),
.B(n_309),
.Y(n_377)
);

AND2x4_ASAP7_75t_L g378 ( 
.A(n_334),
.B(n_191),
.Y(n_378)
);

BUFx8_ASAP7_75t_SL g379 ( 
.A(n_355),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_343),
.Y(n_380)
);

INVx5_ASAP7_75t_L g381 ( 
.A(n_362),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_338),
.B(n_275),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_338),
.B(n_201),
.Y(n_383)
);

INVx5_ASAP7_75t_L g384 ( 
.A(n_324),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_326),
.B(n_301),
.Y(n_385)
);

AND2x4_ASAP7_75t_L g386 ( 
.A(n_340),
.B(n_203),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_322),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_364),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_364),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_340),
.B(n_275),
.Y(n_390)
);

INVx5_ASAP7_75t_L g391 ( 
.A(n_342),
.Y(n_391)
);

BUFx12f_ASAP7_75t_L g392 ( 
.A(n_323),
.Y(n_392)
);

INVx6_ASAP7_75t_L g393 ( 
.A(n_320),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_360),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_360),
.B(n_204),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_361),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_361),
.B(n_300),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_336),
.B(n_209),
.Y(n_398)
);

INVx5_ASAP7_75t_L g399 ( 
.A(n_354),
.Y(n_399)
);

BUFx12f_ASAP7_75t_L g400 ( 
.A(n_329),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_355),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_330),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_346),
.Y(n_403)
);

INVx5_ASAP7_75t_L g404 ( 
.A(n_346),
.Y(n_404)
);

BUFx8_ASAP7_75t_SL g405 ( 
.A(n_366),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_337),
.B(n_294),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_353),
.B(n_300),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_349),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_332),
.B(n_303),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_363),
.B(n_304),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_376),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_373),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_376),
.B(n_353),
.Y(n_413)
);

BUFx12f_ASAP7_75t_L g414 ( 
.A(n_372),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_382),
.B(n_302),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_382),
.B(n_356),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_403),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_403),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_390),
.B(n_302),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_390),
.B(n_274),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_376),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_376),
.B(n_356),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_376),
.B(n_349),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_376),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_387),
.Y(n_425)
);

OA21x2_ASAP7_75t_L g426 ( 
.A1(n_403),
.A2(n_352),
.B(n_350),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_371),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_393),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_367),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_394),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_394),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_371),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_394),
.B(n_350),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_388),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_400),
.Y(n_435)
);

OAI22x1_ASAP7_75t_L g436 ( 
.A1(n_385),
.A2(n_366),
.B1(n_312),
.B2(n_359),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_397),
.B(n_344),
.Y(n_437)
);

OA21x2_ASAP7_75t_L g438 ( 
.A1(n_388),
.A2(n_380),
.B(n_370),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_370),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_393),
.Y(n_440)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_394),
.Y(n_441)
);

OAI21x1_ASAP7_75t_L g442 ( 
.A1(n_389),
.A2(n_352),
.B(n_344),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_393),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_394),
.B(n_319),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_394),
.B(n_319),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_374),
.A2(n_194),
.B1(n_197),
.B2(n_211),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_397),
.A2(n_308),
.B1(n_335),
.B2(n_279),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_370),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_380),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_407),
.A2(n_347),
.B1(n_358),
.B2(n_357),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_396),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_388),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_389),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_407),
.B(n_409),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_398),
.B(n_325),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_396),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_396),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_396),
.Y(n_458)
);

AND2x6_ASAP7_75t_L g459 ( 
.A(n_396),
.B(n_199),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_396),
.Y(n_460)
);

OAI21x1_ASAP7_75t_L g461 ( 
.A1(n_389),
.A2(n_325),
.B(n_313),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_393),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_377),
.B(n_307),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_402),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_389),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_401),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_408),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_408),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_400),
.Y(n_469)
);

NOR2x1_ASAP7_75t_L g470 ( 
.A(n_410),
.B(n_307),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_408),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_408),
.B(n_331),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_408),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_408),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_375),
.Y(n_475)
);

OAI21x1_ASAP7_75t_L g476 ( 
.A1(n_375),
.A2(n_313),
.B(n_199),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_401),
.B(n_341),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_375),
.Y(n_478)
);

BUFx8_ASAP7_75t_L g479 ( 
.A(n_369),
.Y(n_479)
);

OAI22x1_ASAP7_75t_L g480 ( 
.A1(n_379),
.A2(n_351),
.B1(n_365),
.B2(n_273),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_375),
.Y(n_481)
);

AND2x6_ASAP7_75t_L g482 ( 
.A(n_378),
.B(n_210),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_378),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_406),
.A2(n_187),
.B1(n_228),
.B2(n_220),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_400),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_378),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_368),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_368),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_404),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_378),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_368),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_383),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_383),
.Y(n_493)
);

INVx6_ASAP7_75t_L g494 ( 
.A(n_369),
.Y(n_494)
);

OAI21x1_ASAP7_75t_L g495 ( 
.A1(n_404),
.A2(n_218),
.B(n_215),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_383),
.Y(n_496)
);

AND2x6_ASAP7_75t_L g497 ( 
.A(n_383),
.B(n_225),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_386),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_368),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_386),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_386),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_392),
.B(n_268),
.Y(n_502)
);

CKINVDCx11_ASAP7_75t_R g503 ( 
.A(n_392),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_386),
.B(n_268),
.Y(n_504)
);

NOR2x1_ASAP7_75t_L g505 ( 
.A(n_395),
.B(n_398),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_454),
.B(n_398),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_412),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_438),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_488),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_R g510 ( 
.A(n_425),
.B(n_405),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_463),
.B(n_395),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_485),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_427),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_438),
.Y(n_514)
);

CKINVDCx16_ASAP7_75t_R g515 ( 
.A(n_414),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_429),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_432),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_503),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_411),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_438),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_503),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_434),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_480),
.B(n_477),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_449),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_434),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_452),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_435),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_452),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_469),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_466),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_417),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_418),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_450),
.B(n_398),
.Y(n_533)
);

CKINVDCx16_ASAP7_75t_R g534 ( 
.A(n_462),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_504),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_479),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_439),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_488),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_415),
.B(n_395),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_479),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_494),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_412),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_494),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_463),
.B(n_395),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_494),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_448),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_462),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_437),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_443),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_436),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_441),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_437),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_475),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_426),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_426),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_447),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_481),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_416),
.B(n_381),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_413),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_411),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_413),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_422),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_422),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_416),
.B(n_404),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_SL g565 ( 
.A(n_411),
.B(n_197),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_486),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_411),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_R g568 ( 
.A(n_428),
.B(n_185),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_420),
.B(n_404),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_441),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_426),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_421),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_534),
.B(n_419),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_542),
.B(n_472),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_508),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_569),
.B(n_472),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_559),
.B(n_470),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_522),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_508),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_519),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_507),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_514),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_514),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_522),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_519),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_520),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_525),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_569),
.B(n_464),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_539),
.B(n_464),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_520),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_556),
.B(n_440),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_561),
.B(n_486),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_554),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_525),
.Y(n_594)
);

NAND3xp33_ASAP7_75t_L g595 ( 
.A(n_506),
.B(n_484),
.C(n_446),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_562),
.B(n_500),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_526),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_556),
.B(n_502),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_519),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_563),
.B(n_500),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_526),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_528),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_528),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_533),
.B(n_421),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_554),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_555),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_547),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_555),
.Y(n_608)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_519),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_571),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_571),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_509),
.Y(n_612)
);

AND2x6_ASAP7_75t_L g613 ( 
.A(n_612),
.B(n_551),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_598),
.B(n_530),
.Y(n_614)
);

AND2x6_ASAP7_75t_L g615 ( 
.A(n_612),
.B(n_551),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_578),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_607),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_578),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_577),
.B(n_511),
.Y(n_619)
);

BUFx10_ASAP7_75t_L g620 ( 
.A(n_591),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_592),
.B(n_548),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_595),
.A2(n_550),
.B1(n_604),
.B2(n_446),
.Y(n_622)
);

OR2x6_ASAP7_75t_L g623 ( 
.A(n_576),
.B(n_588),
.Y(n_623)
);

NAND3xp33_ASAP7_75t_L g624 ( 
.A(n_574),
.B(n_550),
.C(n_544),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_596),
.A2(n_535),
.B1(n_566),
.B2(n_523),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_584),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_589),
.B(n_558),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_596),
.A2(n_517),
.B1(n_524),
.B2(n_513),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_592),
.B(n_552),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_584),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_587),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_594),
.Y(n_632)
);

BUFx2_ASAP7_75t_L g633 ( 
.A(n_607),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_580),
.Y(n_634)
);

BUFx4f_ASAP7_75t_L g635 ( 
.A(n_580),
.Y(n_635)
);

INVx5_ASAP7_75t_L g636 ( 
.A(n_580),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_607),
.B(n_573),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_594),
.Y(n_638)
);

BUFx10_ASAP7_75t_L g639 ( 
.A(n_581),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_587),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_600),
.B(n_531),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_597),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_581),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_600),
.A2(n_530),
.B1(n_490),
.B2(n_492),
.Y(n_644)
);

OR2x6_ASAP7_75t_L g645 ( 
.A(n_612),
.B(n_505),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_597),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_601),
.B(n_549),
.Y(n_647)
);

INVx2_ASAP7_75t_SL g648 ( 
.A(n_580),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_601),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_609),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_602),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_603),
.Y(n_652)
);

OR2x6_ASAP7_75t_L g653 ( 
.A(n_609),
.B(n_444),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_580),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_602),
.B(n_541),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_580),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_609),
.B(n_549),
.Y(n_657)
);

NAND3xp33_ASAP7_75t_L g658 ( 
.A(n_603),
.B(n_493),
.C(n_483),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_609),
.Y(n_659)
);

INVx4_ASAP7_75t_L g660 ( 
.A(n_585),
.Y(n_660)
);

NAND2xp33_ASAP7_75t_L g661 ( 
.A(n_585),
.B(n_541),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_585),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_585),
.Y(n_663)
);

BUFx10_ASAP7_75t_L g664 ( 
.A(n_585),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_608),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_585),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_599),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_605),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_599),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_608),
.B(n_532),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_579),
.B(n_553),
.Y(n_671)
);

INVxp67_ASAP7_75t_SL g672 ( 
.A(n_575),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_605),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_579),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_593),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_599),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_599),
.B(n_543),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_575),
.B(n_557),
.Y(n_678)
);

INVx4_ASAP7_75t_L g679 ( 
.A(n_599),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_610),
.Y(n_680)
);

INVx5_ASAP7_75t_L g681 ( 
.A(n_599),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_610),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_593),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_575),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_593),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_582),
.B(n_537),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_606),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_582),
.B(n_423),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_606),
.A2(n_222),
.B1(n_497),
.B2(n_482),
.Y(n_689)
);

XOR2xp5_ASAP7_75t_L g690 ( 
.A(n_606),
.B(n_516),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_611),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_611),
.Y(n_692)
);

OAI21xp33_ASAP7_75t_SL g693 ( 
.A1(n_611),
.A2(n_433),
.B(n_423),
.Y(n_693)
);

AO21x2_ASAP7_75t_L g694 ( 
.A1(n_582),
.A2(n_433),
.B(n_476),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_583),
.A2(n_482),
.B1(n_497),
.B2(n_496),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_583),
.Y(n_696)
);

AND2x6_ASAP7_75t_L g697 ( 
.A(n_590),
.B(n_551),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_583),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_672),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_672),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_665),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_680),
.Y(n_702)
);

INVxp67_ASAP7_75t_SL g703 ( 
.A(n_641),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_682),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_639),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_633),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_632),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_635),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_616),
.Y(n_709)
);

XOR2xp5_ASAP7_75t_L g710 ( 
.A(n_690),
.B(n_516),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_618),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_626),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_629),
.B(n_232),
.Y(n_713)
);

INVx4_ASAP7_75t_SL g714 ( 
.A(n_613),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_637),
.B(n_586),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_614),
.B(n_527),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_630),
.Y(n_717)
);

NAND2x1p5_ASAP7_75t_L g718 ( 
.A(n_635),
.B(n_570),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_631),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_620),
.B(n_617),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_640),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_649),
.Y(n_722)
);

INVx4_ASAP7_75t_SL g723 ( 
.A(n_613),
.Y(n_723)
);

INVx5_ASAP7_75t_L g724 ( 
.A(n_613),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_638),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_651),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_687),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_642),
.Y(n_728)
);

INVxp33_ASAP7_75t_L g729 ( 
.A(n_647),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_698),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_670),
.Y(n_731)
);

OAI21xp5_ASAP7_75t_L g732 ( 
.A1(n_624),
.A2(n_497),
.B(n_482),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_621),
.B(n_189),
.Y(n_733)
);

XNOR2x2_ASAP7_75t_L g734 ( 
.A(n_624),
.B(n_189),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_675),
.Y(n_735)
);

BUFx2_ASAP7_75t_L g736 ( 
.A(n_662),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_634),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_683),
.Y(n_738)
);

INVxp67_ASAP7_75t_L g739 ( 
.A(n_643),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_620),
.B(n_527),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_669),
.B(n_547),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_621),
.B(n_189),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_685),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_691),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_655),
.B(n_529),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_692),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_646),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_657),
.B(n_529),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_696),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_634),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_668),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_673),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_674),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_677),
.B(n_586),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_678),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_623),
.B(n_586),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_678),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_652),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_686),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_671),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_671),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_684),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_684),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_625),
.B(n_512),
.Y(n_764)
);

BUFx6f_ASAP7_75t_SL g765 ( 
.A(n_639),
.Y(n_765)
);

NAND2x1p5_ASAP7_75t_L g766 ( 
.A(n_636),
.B(n_681),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_625),
.B(n_512),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_693),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_693),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_622),
.B(n_546),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_688),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_622),
.B(n_543),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_641),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_688),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_623),
.B(n_590),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_623),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_658),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_658),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_666),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_697),
.Y(n_780)
);

CKINVDCx20_ASAP7_75t_R g781 ( 
.A(n_663),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_650),
.B(n_590),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_697),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_697),
.Y(n_784)
);

XOR2xp5_ASAP7_75t_L g785 ( 
.A(n_644),
.B(n_536),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_703),
.B(n_619),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_772),
.A2(n_644),
.B1(n_661),
.B2(n_627),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_741),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_732),
.A2(n_689),
.B(n_695),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_720),
.B(n_628),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_731),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_729),
.B(n_628),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_781),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_745),
.B(n_636),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_716),
.B(n_515),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_773),
.B(n_666),
.Y(n_796)
);

NAND2xp33_ASAP7_75t_SL g797 ( 
.A(n_765),
.B(n_536),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_764),
.A2(n_565),
.B1(n_482),
.B2(n_497),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_740),
.Y(n_799)
);

NOR3xp33_ASAP7_75t_L g800 ( 
.A(n_767),
.B(n_565),
.C(n_501),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_759),
.B(n_774),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_741),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_709),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_760),
.B(n_653),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_734),
.A2(n_776),
.B1(n_785),
.B2(n_770),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_748),
.B(n_705),
.Y(n_806)
);

NAND2xp33_ASAP7_75t_SL g807 ( 
.A(n_765),
.B(n_540),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_701),
.Y(n_808)
);

AND2x6_ASAP7_75t_SL g809 ( 
.A(n_733),
.B(n_540),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_761),
.B(n_653),
.Y(n_810)
);

NAND2x1_ASAP7_75t_L g811 ( 
.A(n_699),
.B(n_700),
.Y(n_811)
);

OAI22xp5_ASAP7_75t_L g812 ( 
.A1(n_724),
.A2(n_689),
.B1(n_695),
.B2(n_681),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_701),
.Y(n_813)
);

INVx4_ASAP7_75t_L g814 ( 
.A(n_737),
.Y(n_814)
);

NAND2xp33_ASAP7_75t_SL g815 ( 
.A(n_708),
.B(n_510),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_715),
.B(n_653),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_702),
.Y(n_817)
);

INVx2_ASAP7_75t_SL g818 ( 
.A(n_737),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_736),
.B(n_518),
.Y(n_819)
);

BUFx12f_ASAP7_75t_L g820 ( 
.A(n_742),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_710),
.B(n_518),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_771),
.B(n_755),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_706),
.B(n_645),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_702),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_771),
.B(n_697),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_739),
.B(n_521),
.Y(n_826)
);

INVxp67_ASAP7_75t_L g827 ( 
.A(n_713),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_704),
.B(n_656),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_757),
.B(n_645),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_708),
.B(n_521),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_724),
.B(n_636),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_711),
.B(n_645),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_712),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_717),
.B(n_648),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_704),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_756),
.B(n_656),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_719),
.B(n_654),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_721),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_737),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_722),
.B(n_650),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_777),
.A2(n_482),
.B1(n_497),
.B2(n_498),
.Y(n_841)
);

BUFx5_ASAP7_75t_L g842 ( 
.A(n_768),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_708),
.B(n_545),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_726),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_751),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_752),
.B(n_659),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_753),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_727),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_699),
.B(n_613),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_SL g850 ( 
.A(n_778),
.B(n_545),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_754),
.B(n_659),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_754),
.B(n_707),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_750),
.B(n_208),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_750),
.B(n_208),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_730),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_735),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_725),
.B(n_615),
.Y(n_857)
);

NOR2xp67_ASAP7_75t_L g858 ( 
.A(n_724),
.B(n_660),
.Y(n_858)
);

BUFx2_ASAP7_75t_L g859 ( 
.A(n_750),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_700),
.B(n_615),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_786),
.B(n_768),
.Y(n_861)
);

AND2x6_ASAP7_75t_SL g862 ( 
.A(n_821),
.B(n_270),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_808),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_799),
.B(n_775),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_822),
.B(n_769),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_822),
.B(n_769),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_803),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_839),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_818),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_833),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_811),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_SL g872 ( 
.A1(n_789),
.A2(n_766),
.B1(n_783),
.B2(n_780),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_806),
.B(n_779),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_813),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_820),
.Y(n_875)
);

NOR3x1_ASAP7_75t_L g876 ( 
.A(n_790),
.B(n_784),
.C(n_310),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_791),
.B(n_738),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_852),
.B(n_743),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_859),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_801),
.B(n_744),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_788),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_838),
.Y(n_882)
);

AND2x6_ASAP7_75t_L g883 ( 
.A(n_787),
.B(n_714),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_828),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_800),
.A2(n_723),
.B1(n_714),
.B2(n_455),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_845),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_804),
.B(n_746),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_805),
.A2(n_226),
.B1(n_227),
.B2(n_190),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_827),
.B(n_728),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_823),
.B(n_749),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_831),
.A2(n_681),
.B(n_718),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_802),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_844),
.B(n_762),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_795),
.B(n_747),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_850),
.B(n_723),
.Y(n_895)
);

AND2x4_ASAP7_75t_SL g896 ( 
.A(n_836),
.B(n_664),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_792),
.B(n_758),
.Y(n_897)
);

NAND2x1_ASAP7_75t_L g898 ( 
.A(n_828),
.B(n_615),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_814),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_836),
.B(n_782),
.Y(n_900)
);

INVxp67_ASAP7_75t_SL g901 ( 
.A(n_849),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_816),
.B(n_782),
.Y(n_902)
);

BUFx8_ASAP7_75t_L g903 ( 
.A(n_815),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_798),
.A2(n_226),
.B1(n_227),
.B2(n_190),
.Y(n_904)
);

A2O1A1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_797),
.A2(n_235),
.B(n_226),
.C(n_227),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_810),
.B(n_763),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_817),
.Y(n_907)
);

INVx8_ASAP7_75t_L g908 ( 
.A(n_793),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_809),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_847),
.B(n_615),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_856),
.B(n_634),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_794),
.A2(n_226),
.B1(n_227),
.B2(n_190),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_832),
.Y(n_913)
);

NOR2xp67_ASAP7_75t_L g914 ( 
.A(n_848),
.B(n_660),
.Y(n_914)
);

INVx2_ASAP7_75t_SL g915 ( 
.A(n_814),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_829),
.B(n_855),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_807),
.B(n_667),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_819),
.B(n_0),
.Y(n_918)
);

NAND2x1p5_ASAP7_75t_L g919 ( 
.A(n_858),
.B(n_679),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_851),
.B(n_679),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_842),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_857),
.B(n_667),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_796),
.B(n_667),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_824),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_835),
.B(n_676),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_834),
.Y(n_926)
);

OAI22xp33_ASAP7_75t_L g927 ( 
.A1(n_789),
.A2(n_676),
.B1(n_570),
.B2(n_560),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_842),
.B(n_676),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_812),
.A2(n_455),
.B1(n_459),
.B2(n_564),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_842),
.B(n_0),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_826),
.B(n_664),
.Y(n_931)
);

OR2x2_ASAP7_75t_L g932 ( 
.A(n_849),
.B(n_860),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_842),
.Y(n_933)
);

O2A1O1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_812),
.A2(n_270),
.B(n_310),
.C(n_311),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_842),
.B(n_1),
.Y(n_935)
);

A2O1A1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_853),
.A2(n_854),
.B(n_843),
.C(n_830),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_860),
.B(n_2),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_825),
.B(n_3),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_840),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_825),
.B(n_568),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_863),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_874),
.Y(n_942)
);

INVx5_ASAP7_75t_L g943 ( 
.A(n_883),
.Y(n_943)
);

INVx2_ASAP7_75t_SL g944 ( 
.A(n_908),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_939),
.B(n_901),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_907),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_932),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_865),
.B(n_837),
.Y(n_948)
);

NAND2xp33_ASAP7_75t_L g949 ( 
.A(n_883),
.B(n_846),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_883),
.A2(n_841),
.B1(n_459),
.B2(n_235),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_926),
.B(n_311),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_884),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_924),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_871),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_867),
.Y(n_955)
);

OAI21xp5_ASAP7_75t_L g956 ( 
.A1(n_905),
.A2(n_207),
.B(n_206),
.Y(n_956)
);

NAND2x1p5_ASAP7_75t_L g957 ( 
.A(n_895),
.B(n_560),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_908),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_908),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_861),
.B(n_3),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_913),
.B(n_884),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_870),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_916),
.B(n_4),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_865),
.B(n_4),
.Y(n_964)
);

BUFx12f_ASAP7_75t_L g965 ( 
.A(n_903),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_866),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_897),
.A2(n_445),
.B(n_444),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_882),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_903),
.Y(n_969)
);

BUFx4f_ASAP7_75t_L g970 ( 
.A(n_883),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_887),
.B(n_878),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_886),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_866),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_893),
.Y(n_974)
);

BUFx3_ASAP7_75t_L g975 ( 
.A(n_875),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_893),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_879),
.B(n_694),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_909),
.B(n_560),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_880),
.B(n_5),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_899),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_877),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_925),
.B(n_864),
.Y(n_982)
);

NOR2x1_ASAP7_75t_L g983 ( 
.A(n_914),
.B(n_694),
.Y(n_983)
);

INVx4_ASAP7_75t_L g984 ( 
.A(n_862),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_890),
.Y(n_985)
);

NOR2x2_ASAP7_75t_L g986 ( 
.A(n_868),
.B(n_468),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_906),
.B(n_5),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_940),
.B(n_6),
.Y(n_988)
);

INVx1_ASAP7_75t_SL g989 ( 
.A(n_937),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_902),
.B(n_920),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_923),
.B(n_7),
.Y(n_991)
);

INVxp67_ASAP7_75t_L g992 ( 
.A(n_889),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_925),
.Y(n_993)
);

AOI22xp33_ASAP7_75t_L g994 ( 
.A1(n_888),
.A2(n_459),
.B1(n_564),
.B2(n_471),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_868),
.Y(n_995)
);

AO22x1_ASAP7_75t_L g996 ( 
.A1(n_876),
.A2(n_570),
.B1(n_8),
.B2(n_9),
.Y(n_996)
);

OR2x6_ASAP7_75t_L g997 ( 
.A(n_891),
.B(n_560),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_873),
.B(n_572),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_921),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_954),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_970),
.A2(n_917),
.B(n_930),
.Y(n_1001)
);

O2A1O1Ixp33_ASAP7_75t_SL g1002 ( 
.A1(n_944),
.A2(n_936),
.B(n_898),
.C(n_918),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_961),
.B(n_900),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_970),
.A2(n_885),
.B1(n_872),
.B2(n_904),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_989),
.B(n_937),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_941),
.Y(n_1006)
);

O2A1O1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_964),
.A2(n_960),
.B(n_989),
.C(n_988),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_984),
.A2(n_935),
.B(n_930),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_949),
.A2(n_935),
.B(n_927),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_984),
.A2(n_938),
.B(n_894),
.Y(n_1010)
);

BUFx4f_ASAP7_75t_L g1011 ( 
.A(n_965),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_956),
.A2(n_938),
.B(n_912),
.Y(n_1012)
);

BUFx2_ASAP7_75t_L g1013 ( 
.A(n_997),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_975),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_956),
.A2(n_929),
.B(n_931),
.C(n_922),
.Y(n_1015)
);

NAND2xp33_ASAP7_75t_L g1016 ( 
.A(n_969),
.B(n_881),
.Y(n_1016)
);

NAND3xp33_ASAP7_75t_L g1017 ( 
.A(n_964),
.B(n_910),
.C(n_911),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_996),
.A2(n_934),
.B(n_928),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_952),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_943),
.A2(n_892),
.B1(n_915),
.B2(n_869),
.Y(n_1020)
);

AOI21x1_ASAP7_75t_L g1021 ( 
.A1(n_951),
.A2(n_933),
.B(n_928),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_995),
.B(n_896),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_945),
.B(n_919),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_945),
.B(n_919),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_993),
.B(n_7),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_950),
.A2(n_212),
.B1(n_213),
.B2(n_216),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_947),
.B(n_8),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_963),
.A2(n_221),
.B(n_217),
.Y(n_1028)
);

OAI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_987),
.A2(n_230),
.B(n_224),
.Y(n_1029)
);

INVx5_ASAP7_75t_L g1030 ( 
.A(n_943),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_SL g1031 ( 
.A1(n_943),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_981),
.B(n_10),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_943),
.A2(n_445),
.B(n_236),
.Y(n_1033)
);

NAND2xp33_ASAP7_75t_L g1034 ( 
.A(n_957),
.B(n_459),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_999),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_958),
.B(n_11),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_948),
.B(n_12),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_959),
.B(n_12),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_957),
.A2(n_572),
.B1(n_567),
.B2(n_233),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_952),
.B(n_13),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_974),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_976),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_992),
.B(n_14),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_997),
.A2(n_474),
.B(n_458),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_997),
.A2(n_468),
.B(n_495),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_948),
.A2(n_538),
.B(n_509),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_942),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_985),
.B(n_14),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_973),
.B(n_15),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_979),
.B(n_15),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_971),
.B(n_16),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_946),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_979),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_982),
.B(n_567),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_998),
.A2(n_538),
.B(n_509),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_978),
.A2(n_538),
.B(n_442),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_980),
.B(n_17),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_967),
.A2(n_491),
.B(n_487),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_991),
.A2(n_499),
.B(n_478),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_980),
.Y(n_1060)
);

HB1xp67_ASAP7_75t_L g1061 ( 
.A(n_966),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_953),
.Y(n_1062)
);

OAI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_982),
.A2(n_459),
.B(n_461),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_955),
.B(n_18),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_994),
.A2(n_572),
.B(n_567),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_977),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1021),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1007),
.B(n_972),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_1060),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1006),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_1003),
.B(n_990),
.Y(n_1071)
);

AOI221xp5_ASAP7_75t_L g1072 ( 
.A1(n_1053),
.A2(n_962),
.B1(n_968),
.B2(n_977),
.C(n_22),
.Y(n_1072)
);

HB1xp67_ASAP7_75t_L g1073 ( 
.A(n_1061),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1008),
.B(n_983),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1062),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1047),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1005),
.B(n_986),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1037),
.B(n_19),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_1030),
.B(n_567),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1010),
.B(n_19),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_1030),
.B(n_20),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1025),
.B(n_20),
.Y(n_1082)
);

AND3x1_ASAP7_75t_L g1083 ( 
.A(n_1050),
.B(n_21),
.C(n_22),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1032),
.B(n_21),
.Y(n_1084)
);

AOI21x1_ASAP7_75t_SL g1085 ( 
.A1(n_1081),
.A2(n_1049),
.B(n_1064),
.Y(n_1085)
);

OR2x2_ASAP7_75t_L g1086 ( 
.A(n_1077),
.B(n_1023),
.Y(n_1086)
);

OA21x2_ASAP7_75t_L g1087 ( 
.A1(n_1067),
.A2(n_1013),
.B(n_1024),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_1067),
.A2(n_1019),
.B(n_1020),
.Y(n_1088)
);

AO21x2_ASAP7_75t_L g1089 ( 
.A1(n_1074),
.A2(n_1051),
.B(n_1027),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_1068),
.A2(n_1019),
.B(n_1035),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1073),
.B(n_1041),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_1080),
.A2(n_1002),
.B(n_1012),
.C(n_1043),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_1073),
.A2(n_1001),
.B(n_1000),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_1076),
.A2(n_1042),
.B(n_1052),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1069),
.B(n_1060),
.Y(n_1095)
);

INVx1_ASAP7_75t_SL g1096 ( 
.A(n_1081),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_1072),
.A2(n_1031),
.B(n_1004),
.Y(n_1097)
);

INVx2_ASAP7_75t_SL g1098 ( 
.A(n_1076),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1070),
.B(n_1075),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_1079),
.A2(n_1009),
.B(n_1044),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_1079),
.A2(n_1054),
.B(n_1017),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1082),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_1084),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_SL g1104 ( 
.A1(n_1078),
.A2(n_1026),
.B(n_1028),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_SL g1105 ( 
.A1(n_1083),
.A2(n_1018),
.B(n_1016),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1071),
.A2(n_1026),
.B(n_1029),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_SL g1107 ( 
.A(n_1081),
.B(n_1031),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_1067),
.A2(n_1040),
.B(n_1045),
.Y(n_1108)
);

AOI21xp33_ASAP7_75t_L g1109 ( 
.A1(n_1080),
.A2(n_1038),
.B(n_1036),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1099),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_1096),
.Y(n_1111)
);

INVx4_ASAP7_75t_L g1112 ( 
.A(n_1103),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1097),
.A2(n_1030),
.B1(n_1011),
.B2(n_1014),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1099),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_1097),
.A2(n_1015),
.B1(n_1014),
.B2(n_1060),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1091),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_1111),
.B(n_1096),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1112),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1117),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_1117),
.B(n_1112),
.Y(n_1120)
);

INVx6_ASAP7_75t_L g1121 ( 
.A(n_1120),
.Y(n_1121)
);

CKINVDCx11_ASAP7_75t_R g1122 ( 
.A(n_1120),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1121),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1122),
.B(n_1119),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1124),
.B(n_1118),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1124),
.B(n_1113),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1123),
.A2(n_1115),
.B(n_1093),
.Y(n_1127)
);

OAI221xp5_ASAP7_75t_L g1128 ( 
.A1(n_1126),
.A2(n_1107),
.B1(n_1116),
.B2(n_1110),
.C(n_1114),
.Y(n_1128)
);

INVxp67_ASAP7_75t_L g1129 ( 
.A(n_1125),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1127),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1129),
.B(n_1103),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1130),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_1131),
.Y(n_1133)
);

A2O1A1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_1132),
.A2(n_1128),
.B(n_1011),
.C(n_1092),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_1134),
.B(n_1103),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1133),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1136),
.B(n_1102),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1135),
.Y(n_1138)
);

NOR3xp33_ASAP7_75t_L g1139 ( 
.A(n_1138),
.B(n_1104),
.C(n_1109),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1137),
.B(n_1089),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1140),
.A2(n_1109),
.B(n_1105),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1139),
.B(n_1095),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1142),
.B(n_1090),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1141),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_1142),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1145),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1143),
.B(n_1144),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_1145),
.B(n_1089),
.Y(n_1148)
);

OR2x2_ASAP7_75t_L g1149 ( 
.A(n_1146),
.B(n_1087),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1148),
.B(n_1088),
.Y(n_1150)
);

XNOR2xp5_ASAP7_75t_L g1151 ( 
.A(n_1149),
.B(n_1147),
.Y(n_1151)
);

INVx2_ASAP7_75t_SL g1152 ( 
.A(n_1150),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_1152),
.Y(n_1153)
);

AOI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1151),
.A2(n_1087),
.B(n_1091),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1153),
.B(n_1014),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1154),
.B(n_1098),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1155),
.B(n_1100),
.Y(n_1157)
);

NAND2x1p5_ASAP7_75t_L g1158 ( 
.A(n_1156),
.B(n_1108),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1157),
.B(n_23),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1158),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_1159),
.Y(n_1161)
);

O2A1O1Ixp5_ASAP7_75t_L g1162 ( 
.A1(n_1160),
.A2(n_1106),
.B(n_1086),
.C(n_26),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1159),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1161),
.B(n_1094),
.Y(n_1164)
);

INVxp67_ASAP7_75t_SL g1165 ( 
.A(n_1163),
.Y(n_1165)
);

OAI221xp5_ASAP7_75t_L g1166 ( 
.A1(n_1162),
.A2(n_1107),
.B1(n_1106),
.B2(n_26),
.C(n_27),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1164),
.B(n_24),
.Y(n_1167)
);

HB1xp67_ASAP7_75t_L g1168 ( 
.A(n_1165),
.Y(n_1168)
);

OAI211xp5_ASAP7_75t_L g1169 ( 
.A1(n_1168),
.A2(n_1166),
.B(n_25),
.C(n_28),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1167),
.B(n_24),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1170),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1169),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1172),
.Y(n_1173)
);

AOI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1171),
.A2(n_1101),
.B1(n_1057),
.B2(n_30),
.Y(n_1174)
);

AOI221xp5_ASAP7_75t_L g1175 ( 
.A1(n_1173),
.A2(n_25),
.B1(n_29),
.B2(n_31),
.C(n_32),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1174),
.A2(n_29),
.B(n_32),
.Y(n_1176)
);

AOI211xp5_ASAP7_75t_L g1177 ( 
.A1(n_1176),
.A2(n_33),
.B(n_34),
.C(n_1033),
.Y(n_1177)
);

OA22x2_ASAP7_75t_L g1178 ( 
.A1(n_1175),
.A2(n_33),
.B1(n_34),
.B2(n_1085),
.Y(n_1178)
);

AOI221xp5_ASAP7_75t_L g1179 ( 
.A1(n_1177),
.A2(n_1022),
.B1(n_1048),
.B2(n_39),
.C(n_40),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1178),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1178),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1180),
.B(n_36),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1181),
.A2(n_38),
.B(n_41),
.Y(n_1183)
);

NOR2x1_ASAP7_75t_L g1184 ( 
.A(n_1179),
.B(n_42),
.Y(n_1184)
);

NAND3xp33_ASAP7_75t_L g1185 ( 
.A(n_1184),
.B(n_404),
.C(n_46),
.Y(n_1185)
);

NOR3x1_ASAP7_75t_L g1186 ( 
.A(n_1182),
.B(n_45),
.C(n_47),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1185),
.A2(n_1183),
.B1(n_49),
.B2(n_50),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1186),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1188),
.B(n_48),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1187),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1190),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1189),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1192),
.B(n_52),
.Y(n_1193)
);

INVx2_ASAP7_75t_SL g1194 ( 
.A(n_1191),
.Y(n_1194)
);

BUFx12f_ASAP7_75t_L g1195 ( 
.A(n_1194),
.Y(n_1195)
);

AOI221xp5_ASAP7_75t_L g1196 ( 
.A1(n_1193),
.A2(n_1039),
.B1(n_56),
.B2(n_57),
.C(n_58),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1195),
.A2(n_55),
.B1(n_59),
.B2(n_63),
.Y(n_1197)
);

NAND4xp25_ASAP7_75t_L g1198 ( 
.A(n_1196),
.B(n_64),
.C(n_65),
.D(n_66),
.Y(n_1198)
);

AOI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1195),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_1199)
);

NAND3xp33_ASAP7_75t_SL g1200 ( 
.A(n_1198),
.B(n_70),
.C(n_71),
.Y(n_1200)
);

NOR3xp33_ASAP7_75t_SL g1201 ( 
.A(n_1197),
.B(n_72),
.C(n_73),
.Y(n_1201)
);

AOI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1199),
.A2(n_74),
.B1(n_75),
.B2(n_77),
.Y(n_1202)
);

NOR4xp25_ASAP7_75t_L g1203 ( 
.A(n_1200),
.B(n_79),
.C(n_82),
.D(n_83),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_1202),
.B(n_84),
.Y(n_1204)
);

AOI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1204),
.A2(n_1201),
.B1(n_86),
.B2(n_87),
.Y(n_1205)
);

AOI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1203),
.A2(n_85),
.B1(n_88),
.B2(n_90),
.Y(n_1206)
);

XNOR2xp5_ASAP7_75t_L g1207 ( 
.A(n_1205),
.B(n_91),
.Y(n_1207)
);

XNOR2xp5_ASAP7_75t_L g1208 ( 
.A(n_1206),
.B(n_92),
.Y(n_1208)
);

AOI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1208),
.A2(n_93),
.B1(n_94),
.B2(n_96),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1207),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1210),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1209),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1211),
.B(n_97),
.Y(n_1213)
);

NOR2x1p5_ASAP7_75t_L g1214 ( 
.A(n_1212),
.B(n_98),
.Y(n_1214)
);

NOR2xp67_ASAP7_75t_L g1215 ( 
.A(n_1214),
.B(n_99),
.Y(n_1215)
);

NOR3xp33_ASAP7_75t_SL g1216 ( 
.A(n_1213),
.B(n_101),
.C(n_102),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1214),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1217),
.A2(n_103),
.B1(n_107),
.B2(n_108),
.Y(n_1218)
);

OAI22xp33_ASAP7_75t_SL g1219 ( 
.A1(n_1215),
.A2(n_1216),
.B1(n_115),
.B2(n_121),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1217),
.A2(n_113),
.B1(n_122),
.B2(n_123),
.Y(n_1220)
);

OAI321xp33_ASAP7_75t_L g1221 ( 
.A1(n_1219),
.A2(n_125),
.A3(n_126),
.B1(n_128),
.B2(n_129),
.C(n_130),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1218),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_SL g1223 ( 
.A1(n_1222),
.A2(n_1220),
.B(n_134),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_1221),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1224),
.A2(n_572),
.B1(n_1034),
.B2(n_137),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1223),
.A2(n_132),
.B(n_135),
.Y(n_1226)
);

OAI22xp33_ASAP7_75t_SL g1227 ( 
.A1(n_1224),
.A2(n_138),
.B1(n_142),
.B2(n_144),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_1226),
.B(n_145),
.Y(n_1228)
);

OA22x2_ASAP7_75t_L g1229 ( 
.A1(n_1227),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1225),
.A2(n_149),
.B(n_150),
.Y(n_1230)
);

NOR2x1p5_ASAP7_75t_L g1231 ( 
.A(n_1228),
.B(n_1230),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1229),
.A2(n_151),
.B(n_153),
.Y(n_1232)
);

NAND3xp33_ASAP7_75t_L g1233 ( 
.A(n_1228),
.B(n_156),
.C(n_160),
.Y(n_1233)
);

AOI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1231),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_1234)
);

OAI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1232),
.A2(n_164),
.B1(n_166),
.B2(n_168),
.Y(n_1235)
);

OAI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1233),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_1236)
);

OAI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1231),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_1237)
);

AO22x2_ASAP7_75t_L g1238 ( 
.A1(n_1231),
.A2(n_177),
.B1(n_178),
.B2(n_456),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_SL g1239 ( 
.A1(n_1231),
.A2(n_421),
.B1(n_460),
.B2(n_467),
.Y(n_1239)
);

OA22x2_ASAP7_75t_L g1240 ( 
.A1(n_1231),
.A2(n_456),
.B1(n_430),
.B2(n_465),
.Y(n_1240)
);

AO22x2_ASAP7_75t_L g1241 ( 
.A1(n_1231),
.A2(n_430),
.B1(n_1065),
.B2(n_1059),
.Y(n_1241)
);

AO22x2_ASAP7_75t_L g1242 ( 
.A1(n_1231),
.A2(n_1055),
.B1(n_453),
.B2(n_1056),
.Y(n_1242)
);

OAI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1231),
.A2(n_431),
.B1(n_473),
.B2(n_467),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1231),
.A2(n_404),
.B1(n_421),
.B2(n_424),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1231),
.A2(n_451),
.B1(n_473),
.B2(n_467),
.Y(n_1245)
);

AOI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1231),
.A2(n_451),
.B1(n_473),
.B2(n_467),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1235),
.A2(n_391),
.B(n_384),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1236),
.B(n_399),
.Y(n_1248)
);

NAND3xp33_ASAP7_75t_L g1249 ( 
.A(n_1238),
.B(n_399),
.C(n_391),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_SL g1250 ( 
.A1(n_1237),
.A2(n_1243),
.B(n_1240),
.Y(n_1250)
);

AO21x2_ASAP7_75t_L g1251 ( 
.A1(n_1244),
.A2(n_1063),
.B(n_1046),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1234),
.B(n_399),
.Y(n_1252)
);

AO21x2_ASAP7_75t_L g1253 ( 
.A1(n_1245),
.A2(n_1058),
.B(n_384),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1242),
.B(n_399),
.Y(n_1254)
);

OA21x2_ASAP7_75t_L g1255 ( 
.A1(n_1241),
.A2(n_1246),
.B(n_1239),
.Y(n_1255)
);

OR2x6_ASAP7_75t_L g1256 ( 
.A(n_1250),
.B(n_1066),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1255),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1254),
.B(n_399),
.Y(n_1258)
);

OR2x2_ASAP7_75t_L g1259 ( 
.A(n_1248),
.B(n_424),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1252),
.A2(n_1247),
.B(n_1249),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1253),
.B(n_399),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1257),
.A2(n_1251),
.B1(n_431),
.B2(n_451),
.Y(n_1262)
);

NAND3xp33_ASAP7_75t_L g1263 ( 
.A(n_1260),
.B(n_431),
.C(n_473),
.Y(n_1263)
);

AOI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1261),
.A2(n_1066),
.B1(n_424),
.B2(n_431),
.Y(n_1264)
);

OAI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1262),
.A2(n_1259),
.B(n_1258),
.Y(n_1265)
);

AOI221xp5_ASAP7_75t_L g1266 ( 
.A1(n_1265),
.A2(n_1264),
.B1(n_1263),
.B2(n_1256),
.C(n_1066),
.Y(n_1266)
);

AOI221xp5_ASAP7_75t_L g1267 ( 
.A1(n_1266),
.A2(n_460),
.B1(n_457),
.B2(n_451),
.C(n_424),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1267),
.A2(n_460),
.B1(n_457),
.B2(n_489),
.Y(n_1268)
);

AOI211xp5_ASAP7_75t_L g1269 ( 
.A1(n_1268),
.A2(n_489),
.B(n_460),
.C(n_457),
.Y(n_1269)
);

AOI211xp5_ASAP7_75t_L g1270 ( 
.A1(n_1269),
.A2(n_489),
.B(n_457),
.C(n_384),
.Y(n_1270)
);


endmodule