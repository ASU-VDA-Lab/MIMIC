module fake_ariane_1411_n_1686 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1686);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1686;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_68),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_81),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_15),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_16),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_56),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_115),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_15),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_125),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_113),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_4),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_34),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_9),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_102),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_23),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_32),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_90),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_120),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_18),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_74),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_153),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_91),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_72),
.Y(n_185)
);

INVxp67_ASAP7_75t_SL g186 ( 
.A(n_13),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_121),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_158),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_60),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_31),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_20),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_130),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_47),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_33),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_140),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_26),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_76),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_108),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_109),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_96),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_40),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_105),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_124),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_1),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_67),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_142),
.Y(n_207)
);

BUFx10_ASAP7_75t_L g208 ( 
.A(n_157),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_22),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_97),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_46),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_156),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_151),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_92),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_51),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_40),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_2),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_160),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_41),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_36),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_110),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_12),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_87),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_35),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_119),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_133),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_57),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_63),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_135),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_69),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_150),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_10),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_88),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_25),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_59),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_111),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_10),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_84),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_149),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_14),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_50),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_2),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_41),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_61),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_101),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_6),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_16),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_21),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_95),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_54),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_44),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_46),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_58),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_29),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_89),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_11),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_127),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_79),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_152),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_82),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_129),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_14),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_24),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_86),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_28),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_52),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_112),
.Y(n_267)
);

BUFx8_ASAP7_75t_SL g268 ( 
.A(n_23),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_44),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_148),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_53),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_144),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_116),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_34),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_143),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_106),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_100),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_139),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_18),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_32),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_64),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_66),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_31),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_13),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_62),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_9),
.Y(n_286)
);

INVxp33_ASAP7_75t_SL g287 ( 
.A(n_27),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_5),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_147),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_159),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_99),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_19),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_39),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_27),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_3),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_55),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_107),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_136),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_12),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_71),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_8),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_26),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_3),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_161),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_114),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_19),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_70),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_20),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_11),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_80),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_85),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_75),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_37),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_126),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_93),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_22),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_103),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_141),
.Y(n_318)
);

BUFx5_ASAP7_75t_L g319 ( 
.A(n_118),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_0),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_50),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_33),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_122),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_132),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_98),
.Y(n_325)
);

BUFx10_ASAP7_75t_L g326 ( 
.A(n_128),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_268),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_256),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_166),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_194),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_194),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_242),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_216),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_191),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_194),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_201),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_194),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_191),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_206),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_194),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_216),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_246),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_246),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_246),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_246),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_225),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_246),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_257),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_174),
.Y(n_349)
);

INVxp33_ASAP7_75t_L g350 ( 
.A(n_168),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_174),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_260),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_211),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_164),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_211),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_267),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_293),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_293),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_171),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_214),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_171),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_214),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_164),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_315),
.Y(n_364)
);

INVxp33_ASAP7_75t_SL g365 ( 
.A(n_165),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_237),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_274),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_169),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_302),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_190),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_177),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_195),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_181),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_197),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_240),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_202),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_191),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_167),
.Y(n_378)
);

INVxp33_ASAP7_75t_L g379 ( 
.A(n_205),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_217),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_180),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_196),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_219),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_241),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_262),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_279),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_165),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_280),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_286),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_295),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_184),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_303),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_252),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_208),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_252),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_316),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_208),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_193),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_200),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_175),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_207),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_210),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_212),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_221),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_227),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_230),
.Y(n_406)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_265),
.Y(n_407)
);

CKINVDCx14_ASAP7_75t_R g408 ( 
.A(n_208),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_333),
.B(n_326),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_335),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_397),
.B(n_341),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_330),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_330),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_335),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_331),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_331),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_337),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_337),
.Y(n_418)
);

NOR2x1_ASAP7_75t_L g419 ( 
.A(n_359),
.B(n_188),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_340),
.Y(n_420)
);

CKINVDCx8_ASAP7_75t_R g421 ( 
.A(n_336),
.Y(n_421)
);

OAI21x1_ASAP7_75t_L g422 ( 
.A1(n_368),
.A2(n_250),
.B(n_249),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_391),
.B(n_231),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_375),
.A2(n_287),
.B1(n_254),
.B2(n_288),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_378),
.B(n_326),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_340),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_342),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_342),
.Y(n_428)
);

INVx5_ASAP7_75t_L g429 ( 
.A(n_368),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_332),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_350),
.B(n_326),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_343),
.Y(n_432)
);

INVx4_ASAP7_75t_L g433 ( 
.A(n_391),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_382),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_379),
.B(n_173),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_343),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_398),
.B(n_231),
.Y(n_437)
);

AND2x6_ASAP7_75t_L g438 ( 
.A(n_398),
.B(n_192),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_344),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_344),
.Y(n_440)
);

OA21x2_ASAP7_75t_L g441 ( 
.A1(n_359),
.A2(n_271),
.B(n_258),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_346),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_352),
.Y(n_443)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_370),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_345),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_345),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_334),
.A2(n_287),
.B1(n_322),
.B2(n_321),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_360),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_347),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_347),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_365),
.A2(n_173),
.B1(n_322),
.B2(n_321),
.Y(n_451)
);

AND2x6_ASAP7_75t_L g452 ( 
.A(n_399),
.B(n_192),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_361),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_393),
.B(n_178),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_361),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_360),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_399),
.B(n_281),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_395),
.B(n_178),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_381),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_381),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_408),
.B(n_289),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_338),
.A2(n_313),
.B1(n_320),
.B2(n_309),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_372),
.Y(n_463)
);

CKINVDCx16_ASAP7_75t_R g464 ( 
.A(n_394),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_349),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_401),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_366),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_377),
.A2(n_313),
.B1(n_320),
.B2(n_222),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_362),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_401),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_362),
.B(n_290),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_402),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_402),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_403),
.B(n_310),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_328),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_403),
.B(n_312),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_404),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_404),
.Y(n_478)
);

BUFx8_ASAP7_75t_L g479 ( 
.A(n_405),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_405),
.B(n_314),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_406),
.B(n_209),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_400),
.A2(n_186),
.B1(n_251),
.B2(n_220),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_444),
.B(n_374),
.Y(n_483)
);

BUFx4f_ASAP7_75t_L g484 ( 
.A(n_460),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_451),
.A2(n_224),
.B1(n_299),
.B2(n_306),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_412),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_412),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_442),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_444),
.B(n_376),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_467),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_440),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_413),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_431),
.B(n_354),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_413),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_431),
.B(n_406),
.Y(n_495)
);

AOI22xp33_ASAP7_75t_L g496 ( 
.A1(n_437),
.A2(n_363),
.B1(n_387),
.B2(n_407),
.Y(n_496)
);

AO21x2_ASAP7_75t_L g497 ( 
.A1(n_422),
.A2(n_373),
.B(n_371),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_440),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_479),
.Y(n_499)
);

NOR3xp33_ASAP7_75t_L g500 ( 
.A(n_447),
.B(n_234),
.C(n_232),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_440),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_440),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_445),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_415),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_479),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_445),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_448),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_433),
.B(n_371),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_435),
.B(n_163),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_435),
.B(n_163),
.Y(n_510)
);

BUFx10_ASAP7_75t_L g511 ( 
.A(n_463),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_L g512 ( 
.A1(n_437),
.A2(n_396),
.B1(n_392),
.B2(n_390),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_481),
.B(n_170),
.Y(n_513)
);

BUFx6f_ASAP7_75t_SL g514 ( 
.A(n_423),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_433),
.B(n_373),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_460),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_416),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_445),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_SL g519 ( 
.A1(n_479),
.A2(n_348),
.B1(n_339),
.B2(n_329),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_445),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_481),
.B(n_170),
.Y(n_521)
);

INVx8_ASAP7_75t_L g522 ( 
.A(n_438),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_416),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_409),
.B(n_172),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_433),
.B(n_380),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_432),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_448),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_443),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_415),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_461),
.B(n_380),
.Y(n_530)
);

AND2x2_ASAP7_75t_SL g531 ( 
.A(n_441),
.B(n_192),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_432),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_433),
.B(n_383),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_409),
.B(n_383),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_460),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_479),
.B(n_172),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_414),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_423),
.B(n_384),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_437),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_437),
.Y(n_540)
);

AOI21x1_ASAP7_75t_L g541 ( 
.A1(n_422),
.A2(n_385),
.B(n_384),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_451),
.A2(n_283),
.B1(n_243),
.B2(n_247),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_416),
.Y(n_543)
);

BUFx4f_ASAP7_75t_L g544 ( 
.A(n_460),
.Y(n_544)
);

NOR2x1p5_ASAP7_75t_L g545 ( 
.A(n_454),
.B(n_327),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_477),
.B(n_385),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_421),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_423),
.B(n_386),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_417),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_417),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_454),
.B(n_176),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_458),
.B(n_176),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_418),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_432),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_416),
.Y(n_555)
);

INVxp33_ASAP7_75t_SL g556 ( 
.A(n_430),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_418),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_427),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g559 ( 
.A1(n_457),
.A2(n_392),
.B1(n_390),
.B2(n_389),
.Y(n_559)
);

CKINVDCx6p67_ASAP7_75t_R g560 ( 
.A(n_464),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_446),
.Y(n_561)
);

INVxp67_ASAP7_75t_SL g562 ( 
.A(n_448),
.Y(n_562)
);

NAND2x1p5_ASAP7_75t_L g563 ( 
.A(n_441),
.B(n_457),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_477),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_416),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_460),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_446),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_446),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_414),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_414),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_477),
.B(n_386),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_416),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_466),
.B(n_388),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_420),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_428),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_423),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_428),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_421),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_449),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_466),
.B(n_388),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_458),
.B(n_179),
.Y(n_581)
);

BUFx8_ASAP7_75t_SL g582 ( 
.A(n_434),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_420),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_449),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_450),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_450),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_459),
.Y(n_587)
);

NOR2x1p5_ASAP7_75t_L g588 ( 
.A(n_411),
.B(n_389),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_420),
.Y(n_589)
);

NAND2xp33_ASAP7_75t_L g590 ( 
.A(n_470),
.B(n_179),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_457),
.B(n_182),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_425),
.B(n_305),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_434),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_459),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_420),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_457),
.B(n_182),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_478),
.Y(n_597)
);

INVxp33_ASAP7_75t_L g598 ( 
.A(n_424),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_420),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_459),
.Y(n_600)
);

OAI21xp33_ASAP7_75t_L g601 ( 
.A1(n_470),
.A2(n_248),
.B(n_292),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_420),
.Y(n_602)
);

NAND3xp33_ASAP7_75t_L g603 ( 
.A(n_478),
.B(n_311),
.C(n_317),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_426),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_478),
.B(n_218),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_478),
.B(n_235),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_480),
.B(n_311),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_456),
.B(n_317),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_472),
.B(n_349),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_472),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_426),
.Y(n_611)
);

CKINVDCx6p67_ASAP7_75t_R g612 ( 
.A(n_475),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_426),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_426),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_473),
.B(n_351),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_473),
.Y(n_616)
);

BUFx4f_ASAP7_75t_L g617 ( 
.A(n_460),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_480),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_453),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_480),
.B(n_318),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_453),
.Y(n_621)
);

BUFx2_ASAP7_75t_L g622 ( 
.A(n_424),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_455),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_456),
.B(n_318),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_426),
.Y(n_625)
);

INVx1_ASAP7_75t_SL g626 ( 
.A(n_475),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_SL g627 ( 
.A1(n_482),
.A2(n_364),
.B1(n_356),
.B2(n_369),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_426),
.Y(n_628)
);

BUFx10_ASAP7_75t_L g629 ( 
.A(n_480),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_436),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_456),
.Y(n_631)
);

AND2x6_ASAP7_75t_L g632 ( 
.A(n_610),
.B(n_419),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_629),
.B(n_447),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_486),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_524),
.B(n_530),
.Y(n_635)
);

A2O1A1Ixp33_ASAP7_75t_L g636 ( 
.A1(n_618),
.A2(n_476),
.B(n_474),
.C(n_419),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_507),
.Y(n_637)
);

NOR2xp67_ASAP7_75t_L g638 ( 
.A(n_488),
.B(n_469),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_539),
.B(n_469),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_539),
.B(n_469),
.Y(n_640)
);

O2A1O1Ixp33_ASAP7_75t_L g641 ( 
.A1(n_534),
.A2(n_482),
.B(n_462),
.C(n_468),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_540),
.B(n_469),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_495),
.B(n_471),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_540),
.B(n_465),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_626),
.B(n_612),
.Y(n_645)
);

BUFx8_ASAP7_75t_L g646 ( 
.A(n_514),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_629),
.B(n_323),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_593),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_576),
.B(n_546),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_493),
.B(n_263),
.Y(n_650)
);

OR2x6_ASAP7_75t_L g651 ( 
.A(n_499),
.B(n_465),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_509),
.B(n_269),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_510),
.B(n_284),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_576),
.B(n_465),
.Y(n_654)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_490),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_629),
.B(n_324),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_629),
.B(n_324),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_597),
.B(n_325),
.Y(n_658)
);

NOR3xp33_ASAP7_75t_L g659 ( 
.A(n_483),
.B(n_294),
.C(n_308),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_592),
.A2(n_203),
.B1(n_185),
.B2(n_307),
.Y(n_660)
);

NOR2xp67_ASAP7_75t_L g661 ( 
.A(n_488),
.B(n_528),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_546),
.B(n_429),
.Y(n_662)
);

OAI221xp5_ASAP7_75t_L g663 ( 
.A1(n_485),
.A2(n_301),
.B1(n_355),
.B2(n_351),
.C(n_353),
.Y(n_663)
);

INVx1_ASAP7_75t_SL g664 ( 
.A(n_612),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_507),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_571),
.B(n_429),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_573),
.B(n_429),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_514),
.A2(n_199),
.B1(n_162),
.B2(n_304),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_622),
.B(n_367),
.Y(n_669)
);

INVxp33_ASAP7_75t_L g670 ( 
.A(n_582),
.Y(n_670)
);

NOR3xp33_ASAP7_75t_L g671 ( 
.A(n_489),
.B(n_353),
.C(n_358),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_573),
.B(n_429),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_499),
.B(n_505),
.Y(n_673)
);

OAI21xp33_ASAP7_75t_L g674 ( 
.A1(n_485),
.A2(n_355),
.B(n_357),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_505),
.B(n_183),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_580),
.B(n_441),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_527),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_527),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_597),
.B(n_319),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_580),
.B(n_410),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_597),
.B(n_319),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_527),
.Y(n_682)
);

OR2x6_ASAP7_75t_L g683 ( 
.A(n_622),
.B(n_545),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_564),
.B(n_319),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_564),
.B(n_319),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_631),
.Y(n_686)
);

OAI22xp33_ASAP7_75t_L g687 ( 
.A1(n_598),
.A2(n_358),
.B1(n_410),
.B2(n_436),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_511),
.B(n_410),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_528),
.B(n_410),
.Y(n_689)
);

NAND3xp33_ASAP7_75t_L g690 ( 
.A(n_542),
.B(n_436),
.C(n_439),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_588),
.B(n_610),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_513),
.B(n_0),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_588),
.B(n_187),
.Y(n_693)
);

NOR2x1p5_ASAP7_75t_L g694 ( 
.A(n_560),
.B(n_189),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_537),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_521),
.B(n_1),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_560),
.B(n_4),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_516),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_511),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_616),
.B(n_605),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_563),
.B(n_319),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_551),
.B(n_5),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_606),
.B(n_198),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_552),
.B(n_6),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_L g705 ( 
.A(n_501),
.B(n_438),
.Y(n_705)
);

CKINVDCx11_ASAP7_75t_R g706 ( 
.A(n_511),
.Y(n_706)
);

INVxp67_ASAP7_75t_L g707 ( 
.A(n_547),
.Y(n_707)
);

NAND3xp33_ASAP7_75t_L g708 ( 
.A(n_603),
.B(n_436),
.C(n_439),
.Y(n_708)
);

NOR2xp67_ASAP7_75t_L g709 ( 
.A(n_547),
.B(n_436),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_556),
.B(n_204),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_508),
.B(n_213),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_578),
.B(n_436),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_487),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_515),
.B(n_215),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_487),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_525),
.B(n_223),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_533),
.B(n_226),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_563),
.B(n_319),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_559),
.B(n_228),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_538),
.B(n_229),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_492),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_537),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_492),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_531),
.A2(n_438),
.B1(n_452),
.B2(n_439),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_548),
.B(n_233),
.Y(n_725)
);

OAI22xp5_ASAP7_75t_L g726 ( 
.A1(n_619),
.A2(n_296),
.B1(n_259),
.B2(n_255),
.Y(n_726)
);

BUFx10_ASAP7_75t_L g727 ( 
.A(n_545),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_494),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_581),
.B(n_7),
.Y(n_729)
);

INVx8_ASAP7_75t_L g730 ( 
.A(n_522),
.Y(n_730)
);

BUFx6f_ASAP7_75t_SL g731 ( 
.A(n_519),
.Y(n_731)
);

HB1xp67_ASAP7_75t_L g732 ( 
.A(n_514),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_621),
.B(n_236),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_569),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_496),
.B(n_439),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_531),
.A2(n_438),
.B1(n_452),
.B2(n_439),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_536),
.B(n_7),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_512),
.B(n_8),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_621),
.B(n_277),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_623),
.B(n_275),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_623),
.B(n_278),
.Y(n_741)
);

BUFx12f_ASAP7_75t_L g742 ( 
.A(n_609),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_627),
.B(n_17),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_500),
.A2(n_238),
.B1(n_245),
.B2(n_253),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_562),
.B(n_609),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_615),
.B(n_282),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_494),
.A2(n_239),
.B(n_244),
.Y(n_747)
);

HB1xp67_ASAP7_75t_L g748 ( 
.A(n_497),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_570),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_601),
.B(n_291),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_501),
.B(n_319),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_504),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_608),
.Y(n_753)
);

NOR2xp67_ASAP7_75t_L g754 ( 
.A(n_603),
.B(n_261),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_601),
.B(n_297),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_624),
.B(n_285),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_491),
.B(n_319),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_491),
.B(n_273),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_498),
.B(n_273),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_498),
.B(n_502),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_502),
.B(n_272),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_591),
.B(n_17),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_596),
.B(n_21),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_503),
.B(n_300),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_607),
.B(n_24),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_506),
.B(n_298),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_504),
.Y(n_767)
);

OR2x2_ASAP7_75t_L g768 ( 
.A(n_620),
.B(n_25),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_SL g769 ( 
.A(n_522),
.B(n_270),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_506),
.B(n_266),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_590),
.B(n_518),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_518),
.B(n_264),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_520),
.B(n_452),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_517),
.Y(n_774)
);

OR2x6_ASAP7_75t_L g775 ( 
.A(n_522),
.B(n_276),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_526),
.Y(n_776)
);

HB1xp67_ASAP7_75t_L g777 ( 
.A(n_497),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_516),
.B(n_276),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_532),
.Y(n_779)
);

NAND2xp33_ASAP7_75t_L g780 ( 
.A(n_529),
.B(n_452),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_484),
.B(n_192),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_683),
.B(n_529),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_645),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_643),
.B(n_587),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_682),
.B(n_516),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_634),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_648),
.Y(n_787)
);

NOR3xp33_ASAP7_75t_SL g788 ( 
.A(n_710),
.B(n_575),
.C(n_549),
.Y(n_788)
);

AND2x6_ASAP7_75t_L g789 ( 
.A(n_730),
.B(n_549),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_713),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_715),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_706),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_SL g793 ( 
.A(n_691),
.B(n_550),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_648),
.B(n_531),
.Y(n_794)
);

OR2x2_ASAP7_75t_SL g795 ( 
.A(n_697),
.B(n_550),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_655),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_730),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_721),
.Y(n_798)
);

NAND3xp33_ASAP7_75t_SL g799 ( 
.A(n_744),
.B(n_579),
.C(n_557),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_643),
.B(n_635),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_723),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_635),
.A2(n_579),
.B1(n_553),
.B2(n_557),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_649),
.B(n_745),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_679),
.A2(n_484),
.B(n_544),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_SL g805 ( 
.A1(n_663),
.A2(n_575),
.B1(n_586),
.B2(n_585),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_728),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_633),
.B(n_553),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_752),
.Y(n_808)
);

AOI22xp5_ASAP7_75t_L g809 ( 
.A1(n_762),
.A2(n_577),
.B1(n_584),
.B2(n_585),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_682),
.B(n_516),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_700),
.B(n_594),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_767),
.Y(n_812)
);

NOR2x1_ASAP7_75t_L g813 ( 
.A(n_661),
.B(n_517),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_743),
.A2(n_594),
.B1(n_600),
.B2(n_577),
.Y(n_814)
);

NAND3xp33_ASAP7_75t_L g815 ( 
.A(n_692),
.B(n_586),
.C(n_558),
.Y(n_815)
);

NOR2x2_ASAP7_75t_L g816 ( 
.A(n_683),
.B(n_630),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_646),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_753),
.B(n_600),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_712),
.B(n_558),
.Y(n_819)
);

INVx5_ASAP7_75t_L g820 ( 
.A(n_730),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_680),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_639),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_640),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_642),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_760),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_695),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_682),
.B(n_535),
.Y(n_827)
);

AND3x1_ASAP7_75t_L g828 ( 
.A(n_659),
.B(n_583),
.C(n_628),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_776),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_632),
.B(n_554),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_738),
.A2(n_567),
.B1(n_554),
.B2(n_561),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_722),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_698),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_664),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_676),
.A2(n_568),
.B1(n_561),
.B2(n_567),
.Y(n_835)
);

INVx2_ASAP7_75t_SL g836 ( 
.A(n_655),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_779),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_762),
.A2(n_543),
.B1(n_628),
.B2(n_625),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_632),
.B(n_568),
.Y(n_839)
);

O2A1O1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_641),
.A2(n_589),
.B(n_628),
.C(n_625),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_683),
.B(n_555),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_734),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_742),
.B(n_689),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_698),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_749),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_746),
.B(n_674),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_637),
.Y(n_847)
);

BUFx2_ASAP7_75t_SL g848 ( 
.A(n_732),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_698),
.Y(n_849)
);

INVx4_ASAP7_75t_L g850 ( 
.A(n_775),
.Y(n_850)
);

INVx4_ASAP7_75t_L g851 ( 
.A(n_775),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_698),
.B(n_566),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_654),
.Y(n_853)
);

AND2x2_ASAP7_75t_SL g854 ( 
.A(n_737),
.B(n_617),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_665),
.Y(n_855)
);

AND2x6_ASAP7_75t_L g856 ( 
.A(n_737),
.B(n_735),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_688),
.B(n_595),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_763),
.A2(n_765),
.B1(n_692),
.B2(n_696),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_707),
.B(n_555),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_677),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_678),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_652),
.B(n_555),
.Y(n_862)
);

BUFx8_ASAP7_75t_L g863 ( 
.A(n_731),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_644),
.Y(n_864)
);

OR2x6_ASAP7_75t_L g865 ( 
.A(n_732),
.B(n_522),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_686),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_763),
.A2(n_497),
.B1(n_522),
.B2(n_452),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_771),
.B(n_566),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_667),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_731),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_727),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_765),
.A2(n_438),
.B1(n_452),
.B2(n_611),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_651),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_771),
.B(n_566),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_699),
.B(n_555),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_652),
.B(n_583),
.Y(n_876)
);

INVx8_ASAP7_75t_L g877 ( 
.A(n_775),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_650),
.B(n_541),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_702),
.B(n_565),
.Y(n_879)
);

AND2x6_ASAP7_75t_SL g880 ( 
.A(n_702),
.B(n_28),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_653),
.B(n_583),
.Y(n_881)
);

OR2x2_ASAP7_75t_SL g882 ( 
.A(n_669),
.B(n_630),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_774),
.Y(n_883)
);

OR2x6_ASAP7_75t_L g884 ( 
.A(n_694),
.B(n_613),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_704),
.B(n_729),
.Y(n_885)
);

AND2x6_ASAP7_75t_SL g886 ( 
.A(n_704),
.B(n_29),
.Y(n_886)
);

NOR2xp67_ASAP7_75t_L g887 ( 
.A(n_668),
.B(n_517),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_729),
.B(n_565),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_651),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_696),
.B(n_565),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_638),
.B(n_565),
.Y(n_891)
);

CKINVDCx20_ASAP7_75t_R g892 ( 
.A(n_727),
.Y(n_892)
);

BUFx4f_ASAP7_75t_SL g893 ( 
.A(n_675),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_672),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_653),
.B(n_589),
.Y(n_895)
);

AOI21xp33_ASAP7_75t_L g896 ( 
.A1(n_650),
.A2(n_574),
.B(n_572),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_651),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_687),
.B(n_543),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_687),
.B(n_543),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_748),
.B(n_535),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_748),
.B(n_535),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_662),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_751),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_777),
.B(n_535),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_660),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_768),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_773),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_751),
.Y(n_908)
);

A2O1A1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_636),
.A2(n_523),
.B(n_630),
.C(n_614),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_757),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_777),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_757),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_709),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_666),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_L g915 ( 
.A1(n_750),
.A2(n_755),
.B1(n_690),
.B2(n_719),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_733),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_754),
.A2(n_572),
.B(n_614),
.C(n_613),
.Y(n_917)
);

CKINVDCx20_ASAP7_75t_R g918 ( 
.A(n_670),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_658),
.B(n_535),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_739),
.Y(n_920)
);

NOR3xp33_ASAP7_75t_SL g921 ( 
.A(n_658),
.B(n_647),
.C(n_656),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_720),
.B(n_574),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_673),
.Y(n_923)
);

INVx4_ASAP7_75t_L g924 ( 
.A(n_769),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_671),
.B(n_541),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_701),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_758),
.Y(n_927)
);

INVxp67_ASAP7_75t_SL g928 ( 
.A(n_780),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_701),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_725),
.B(n_599),
.Y(n_930)
);

AND2x6_ASAP7_75t_L g931 ( 
.A(n_724),
.B(n_611),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_740),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_761),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_759),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_764),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_741),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_703),
.B(n_604),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_766),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_L g939 ( 
.A1(n_656),
.A2(n_438),
.B1(n_604),
.B2(n_602),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_SL g940 ( 
.A(n_693),
.B(n_599),
.Y(n_940)
);

INVx4_ASAP7_75t_L g941 ( 
.A(n_705),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_770),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_786),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_800),
.A2(n_681),
.B(n_679),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_803),
.B(n_657),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_844),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_885),
.B(n_726),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_826),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_817),
.Y(n_949)
);

O2A1O1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_916),
.A2(n_756),
.B(n_714),
.C(n_717),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_858),
.A2(n_708),
.B1(n_716),
.B2(n_711),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_807),
.A2(n_685),
.B(n_684),
.C(n_718),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_905),
.B(n_718),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_SL g954 ( 
.A1(n_859),
.A2(n_747),
.B(n_772),
.C(n_736),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_787),
.B(n_724),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_787),
.B(n_684),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_790),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_782),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_834),
.Y(n_959)
);

OAI21x1_ASAP7_75t_L g960 ( 
.A1(n_868),
.A2(n_778),
.B(n_781),
.Y(n_960)
);

INVx6_ASAP7_75t_SL g961 ( 
.A(n_884),
.Y(n_961)
);

INVx5_ASAP7_75t_L g962 ( 
.A(n_865),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_791),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_920),
.A2(n_778),
.B(n_736),
.C(n_36),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_798),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_801),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_806),
.Y(n_967)
);

OAI21x1_ASAP7_75t_L g968 ( 
.A1(n_868),
.A2(n_566),
.B(n_438),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_782),
.B(n_30),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_796),
.B(n_30),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_819),
.A2(n_566),
.B(n_276),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_932),
.A2(n_35),
.B(n_37),
.C(n_38),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_832),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_836),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_936),
.B(n_38),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_808),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_L g977 ( 
.A1(n_802),
.A2(n_809),
.B1(n_805),
.B2(n_812),
.Y(n_977)
);

INVx4_ASAP7_75t_L g978 ( 
.A(n_797),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_841),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_794),
.B(n_795),
.Y(n_980)
);

INVx1_ASAP7_75t_SL g981 ( 
.A(n_911),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_844),
.Y(n_982)
);

NAND2xp33_ASAP7_75t_L g983 ( 
.A(n_789),
.B(n_192),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_938),
.B(n_39),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_841),
.B(n_42),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_942),
.B(n_42),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_811),
.A2(n_876),
.B(n_862),
.Y(n_987)
);

AO32x1_ASAP7_75t_L g988 ( 
.A1(n_878),
.A2(n_43),
.A3(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_799),
.A2(n_43),
.B(n_45),
.C(n_48),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_846),
.A2(n_273),
.B1(n_49),
.B2(n_65),
.Y(n_990)
);

BUFx6f_ASAP7_75t_SL g991 ( 
.A(n_884),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_842),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_792),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_854),
.B(n_49),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_843),
.B(n_73),
.Y(n_995)
);

A2O1A1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_876),
.A2(n_77),
.B(n_78),
.C(n_83),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_821),
.B(n_94),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_829),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_788),
.A2(n_104),
.B(n_131),
.C(n_134),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_881),
.A2(n_137),
.B(n_138),
.C(n_146),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_845),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_SL g1002 ( 
.A(n_924),
.B(n_154),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_881),
.A2(n_155),
.B(n_895),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_837),
.Y(n_1004)
);

CKINVDCx12_ASAP7_75t_R g1005 ( 
.A(n_884),
.Y(n_1005)
);

AOI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_856),
.A2(n_854),
.B1(n_793),
.B2(n_889),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_844),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_906),
.B(n_893),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_853),
.B(n_864),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_R g1010 ( 
.A(n_871),
.B(n_892),
.Y(n_1010)
);

BUFx4f_ASAP7_75t_L g1011 ( 
.A(n_897),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_844),
.Y(n_1012)
);

AOI22x1_ASAP7_75t_L g1013 ( 
.A1(n_804),
.A2(n_933),
.B1(n_894),
.B2(n_869),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_825),
.B(n_911),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_895),
.A2(n_928),
.B(n_922),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_SL g1016 ( 
.A(n_924),
.B(n_877),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_788),
.A2(n_840),
.B(n_888),
.C(n_879),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_793),
.A2(n_921),
.B(n_815),
.C(n_935),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_928),
.A2(n_930),
.B(n_937),
.Y(n_1019)
);

NOR2xp67_ASAP7_75t_L g1020 ( 
.A(n_870),
.B(n_783),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_897),
.B(n_820),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_863),
.Y(n_1022)
);

BUFx2_ASAP7_75t_L g1023 ( 
.A(n_882),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_822),
.B(n_823),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_866),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_909),
.A2(n_925),
.B(n_899),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_893),
.B(n_933),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_859),
.B(n_935),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_923),
.B(n_873),
.Y(n_1029)
);

NAND2xp33_ASAP7_75t_L g1030 ( 
.A(n_789),
.B(n_797),
.Y(n_1030)
);

O2A1O1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_890),
.A2(n_921),
.B(n_857),
.C(n_919),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_852),
.A2(n_874),
.B(n_891),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_873),
.B(n_889),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_856),
.A2(n_897),
.B1(n_814),
.B2(n_828),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_818),
.B(n_883),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_824),
.B(n_856),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_814),
.A2(n_898),
.B1(n_867),
.B2(n_831),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_856),
.B(n_848),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_847),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_918),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_852),
.A2(n_785),
.B(n_827),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_820),
.B(n_797),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_860),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_785),
.A2(n_827),
.B(n_810),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_887),
.A2(n_896),
.B(n_926),
.C(n_929),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_SL g1046 ( 
.A1(n_856),
.A2(n_877),
.B1(n_880),
.B2(n_886),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_820),
.B(n_875),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_910),
.A2(n_912),
.B(n_903),
.C(n_908),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_867),
.A2(n_831),
.B1(n_941),
.B2(n_838),
.Y(n_1049)
);

INVx4_ASAP7_75t_L g1050 ( 
.A(n_877),
.Y(n_1050)
);

A2O1A1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_915),
.A2(n_902),
.B(n_914),
.C(n_830),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_865),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_865),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_861),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_833),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_855),
.A2(n_813),
.B(n_902),
.C(n_914),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_833),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_855),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_907),
.A2(n_839),
.B(n_849),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_789),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_900),
.A2(n_904),
.B(n_901),
.Y(n_1061)
);

AOI22xp33_ASAP7_75t_L g1062 ( 
.A1(n_931),
.A2(n_915),
.B1(n_913),
.B2(n_940),
.Y(n_1062)
);

INVxp67_ASAP7_75t_L g1063 ( 
.A(n_931),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_835),
.B(n_931),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_850),
.B(n_851),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_789),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_927),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_1013),
.A2(n_934),
.B(n_939),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_1004),
.Y(n_1069)
);

INVx8_ASAP7_75t_L g1070 ( 
.A(n_962),
.Y(n_1070)
);

OAI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_987),
.A2(n_939),
.B(n_789),
.Y(n_1071)
);

AOI211x1_ASAP7_75t_L g1072 ( 
.A1(n_977),
.A2(n_816),
.B(n_931),
.C(n_872),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_977),
.A2(n_850),
.B1(n_851),
.B2(n_947),
.Y(n_1073)
);

O2A1O1Ixp5_ASAP7_75t_L g1074 ( 
.A1(n_1003),
.A2(n_951),
.B(n_1026),
.C(n_990),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_1015),
.A2(n_983),
.B(n_1019),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_958),
.B(n_969),
.Y(n_1076)
);

AO21x1_ASAP7_75t_L g1077 ( 
.A1(n_990),
.A2(n_1049),
.B(n_951),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_943),
.Y(n_1078)
);

NOR2x1_ASAP7_75t_SL g1079 ( 
.A(n_962),
.B(n_1060),
.Y(n_1079)
);

AOI221x1_ASAP7_75t_L g1080 ( 
.A1(n_1018),
.A2(n_1051),
.B1(n_1045),
.B2(n_1037),
.C(n_1061),
.Y(n_1080)
);

INVx5_ASAP7_75t_L g1081 ( 
.A(n_1052),
.Y(n_1081)
);

OAI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_945),
.A2(n_1028),
.B(n_1017),
.Y(n_1082)
);

NAND3xp33_ASAP7_75t_L g1083 ( 
.A(n_989),
.B(n_972),
.C(n_975),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_1026),
.A2(n_944),
.B(n_952),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1009),
.B(n_1024),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_960),
.A2(n_1041),
.B(n_1044),
.Y(n_1086)
);

NAND3xp33_ASAP7_75t_L g1087 ( 
.A(n_984),
.B(n_986),
.C(n_994),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_1050),
.B(n_979),
.Y(n_1088)
);

BUFx5_ASAP7_75t_L g1089 ( 
.A(n_1067),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_SL g1090 ( 
.A1(n_1049),
.A2(n_1037),
.B(n_995),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_1050),
.B(n_962),
.Y(n_1091)
);

INVxp67_ASAP7_75t_SL g1092 ( 
.A(n_1014),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1009),
.B(n_1024),
.Y(n_1093)
);

AOI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_953),
.A2(n_980),
.B1(n_955),
.B2(n_1006),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1014),
.B(n_1035),
.Y(n_1095)
);

NOR2xp67_ASAP7_75t_SL g1096 ( 
.A(n_993),
.B(n_959),
.Y(n_1096)
);

AO21x2_ASAP7_75t_L g1097 ( 
.A1(n_1064),
.A2(n_1036),
.B(n_971),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_956),
.A2(n_1034),
.B1(n_1062),
.B2(n_985),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_974),
.B(n_981),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_1033),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_1031),
.A2(n_1048),
.B(n_964),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_1010),
.Y(n_1102)
);

HB1xp67_ASAP7_75t_L g1103 ( 
.A(n_1058),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_997),
.A2(n_954),
.B(n_1030),
.Y(n_1104)
);

INVxp67_ASAP7_75t_SL g1105 ( 
.A(n_985),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_1036),
.A2(n_1063),
.B1(n_1027),
.B2(n_976),
.Y(n_1106)
);

OAI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1059),
.A2(n_997),
.B(n_999),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_1040),
.B(n_1008),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_957),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1029),
.B(n_965),
.Y(n_1110)
);

OR2x2_ASAP7_75t_L g1111 ( 
.A(n_963),
.B(n_966),
.Y(n_1111)
);

OR2x6_ASAP7_75t_L g1112 ( 
.A(n_1038),
.B(n_949),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_996),
.A2(n_1000),
.B(n_1002),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_967),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_1066),
.A2(n_1056),
.B(n_1021),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_970),
.A2(n_1047),
.B(n_1042),
.Y(n_1116)
);

INVxp67_ASAP7_75t_L g1117 ( 
.A(n_1025),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_998),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_992),
.Y(n_1119)
);

A2O1A1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_1002),
.A2(n_1046),
.B(n_1023),
.C(n_1020),
.Y(n_1120)
);

AO31x2_ASAP7_75t_L g1121 ( 
.A1(n_948),
.A2(n_973),
.A3(n_1001),
.B(n_1043),
.Y(n_1121)
);

INVxp67_ASAP7_75t_L g1122 ( 
.A(n_1039),
.Y(n_1122)
);

NAND2x1p5_ASAP7_75t_L g1123 ( 
.A(n_1011),
.B(n_962),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1054),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1016),
.B(n_1065),
.Y(n_1125)
);

OR2x6_ASAP7_75t_L g1126 ( 
.A(n_1052),
.B(n_1022),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1011),
.B(n_1053),
.Y(n_1127)
);

AOI21x1_ASAP7_75t_L g1128 ( 
.A1(n_988),
.A2(n_946),
.B(n_1012),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_991),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1055),
.B(n_1057),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_946),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1055),
.B(n_1057),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_1055),
.B(n_982),
.Y(n_1133)
);

O2A1O1Ixp5_ASAP7_75t_SL g1134 ( 
.A1(n_988),
.A2(n_1005),
.B(n_961),
.C(n_982),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_982),
.B(n_1007),
.Y(n_1135)
);

AND2x2_ASAP7_75t_SL g1136 ( 
.A(n_1007),
.B(n_1012),
.Y(n_1136)
);

AOI221x1_ASAP7_75t_L g1137 ( 
.A1(n_1007),
.A2(n_990),
.B1(n_885),
.B2(n_977),
.C(n_1003),
.Y(n_1137)
);

AND3x2_ASAP7_75t_L g1138 ( 
.A(n_988),
.B(n_978),
.C(n_434),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_978),
.A2(n_800),
.B1(n_858),
.B2(n_885),
.Y(n_1139)
);

OAI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_947),
.A2(n_858),
.B1(n_800),
.B2(n_885),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_987),
.A2(n_1003),
.B(n_1015),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_958),
.B(n_787),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1013),
.A2(n_968),
.B(n_1032),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_SL g1144 ( 
.A1(n_977),
.A2(n_1017),
.B(n_945),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_1028),
.B(n_858),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_SL g1146 ( 
.A1(n_950),
.A2(n_784),
.B(n_885),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1009),
.B(n_800),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_943),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1013),
.A2(n_968),
.B(n_1032),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_977),
.A2(n_800),
.B1(n_858),
.B2(n_885),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_947),
.A2(n_858),
.B(n_885),
.C(n_800),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_958),
.B(n_787),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_959),
.Y(n_1153)
);

INVx4_ASAP7_75t_L g1154 ( 
.A(n_959),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_962),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_953),
.B(n_556),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_SL g1157 ( 
.A1(n_950),
.A2(n_784),
.B(n_885),
.Y(n_1157)
);

O2A1O1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_977),
.A2(n_800),
.B(n_885),
.C(n_947),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_943),
.Y(n_1159)
);

OAI22x1_ASAP7_75t_L g1160 ( 
.A1(n_980),
.A2(n_858),
.B1(n_743),
.B2(n_485),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_987),
.A2(n_1003),
.B(n_1015),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_987),
.A2(n_1003),
.B(n_1015),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_953),
.B(n_556),
.Y(n_1163)
);

AO31x2_ASAP7_75t_L g1164 ( 
.A1(n_1037),
.A2(n_917),
.A3(n_1051),
.B(n_1049),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1013),
.A2(n_968),
.B(n_1032),
.Y(n_1165)
);

AOI21x1_ASAP7_75t_L g1166 ( 
.A1(n_987),
.A2(n_1015),
.B(n_1019),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_949),
.Y(n_1167)
);

NAND2xp33_ASAP7_75t_SL g1168 ( 
.A(n_1010),
.B(n_800),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1013),
.A2(n_968),
.B(n_1032),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_987),
.A2(n_800),
.B(n_885),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_987),
.A2(n_1003),
.B(n_1015),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1009),
.B(n_800),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1009),
.B(n_800),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_987),
.A2(n_1003),
.B(n_1015),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1009),
.B(n_800),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1013),
.A2(n_968),
.B(n_1032),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_987),
.A2(n_1003),
.B(n_1015),
.Y(n_1177)
);

INVx1_ASAP7_75t_SL g1178 ( 
.A(n_974),
.Y(n_1178)
);

AO31x2_ASAP7_75t_L g1179 ( 
.A1(n_1037),
.A2(n_917),
.A3(n_1051),
.B(n_1049),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_947),
.A2(n_858),
.B(n_885),
.C(n_800),
.Y(n_1180)
);

NAND3xp33_ASAP7_75t_SL g1181 ( 
.A(n_947),
.B(n_528),
.C(n_488),
.Y(n_1181)
);

NAND2xp33_ASAP7_75t_L g1182 ( 
.A(n_947),
.B(n_800),
.Y(n_1182)
);

AO31x2_ASAP7_75t_L g1183 ( 
.A1(n_1037),
.A2(n_917),
.A3(n_1051),
.B(n_1049),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1009),
.B(n_800),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_977),
.A2(n_800),
.B1(n_858),
.B2(n_885),
.Y(n_1185)
);

OAI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_947),
.A2(n_858),
.B1(n_800),
.B2(n_885),
.Y(n_1186)
);

AO32x2_ASAP7_75t_L g1187 ( 
.A1(n_1037),
.A2(n_990),
.A3(n_977),
.B1(n_1049),
.B2(n_951),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_943),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_953),
.B(n_556),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_943),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1050),
.B(n_841),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_1011),
.Y(n_1192)
);

NAND2x1p5_ASAP7_75t_L g1193 ( 
.A(n_1011),
.B(n_1050),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_1028),
.B(n_858),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_947),
.A2(n_858),
.B(n_885),
.C(n_800),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_SL g1196 ( 
.A1(n_977),
.A2(n_1017),
.B(n_945),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1009),
.B(n_800),
.Y(n_1197)
);

INVx5_ASAP7_75t_L g1198 ( 
.A(n_1052),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_962),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_958),
.B(n_787),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1009),
.B(n_800),
.Y(n_1201)
);

AND2x6_ASAP7_75t_L g1202 ( 
.A(n_1034),
.B(n_1060),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1076),
.B(n_1142),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1152),
.B(n_1200),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_1150),
.B(n_1185),
.Y(n_1205)
);

INVx3_ASAP7_75t_L g1206 ( 
.A(n_1192),
.Y(n_1206)
);

OAI22xp33_ASAP7_75t_SL g1207 ( 
.A1(n_1145),
.A2(n_1194),
.B1(n_1094),
.B2(n_1095),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_1091),
.B(n_1081),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1078),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_SL g1210 ( 
.A1(n_1144),
.A2(n_1196),
.B(n_1077),
.Y(n_1210)
);

AO21x2_ASAP7_75t_L g1211 ( 
.A1(n_1107),
.A2(n_1090),
.B(n_1104),
.Y(n_1211)
);

NAND2x1p5_ASAP7_75t_L g1212 ( 
.A(n_1081),
.B(n_1198),
.Y(n_1212)
);

AOI22x1_ASAP7_75t_L g1213 ( 
.A1(n_1170),
.A2(n_1177),
.B1(n_1171),
.B2(n_1174),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1165),
.A2(n_1176),
.B(n_1169),
.Y(n_1214)
);

OA21x2_ASAP7_75t_L g1215 ( 
.A1(n_1074),
.A2(n_1080),
.B(n_1137),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1087),
.A2(n_1156),
.B1(n_1189),
.B2(n_1163),
.Y(n_1216)
);

INVx2_ASAP7_75t_SL g1217 ( 
.A(n_1167),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1086),
.A2(n_1166),
.B(n_1068),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1113),
.A2(n_1182),
.B(n_1158),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1109),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1114),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1084),
.A2(n_1115),
.B(n_1071),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_1136),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1087),
.A2(n_1151),
.B(n_1180),
.Y(n_1224)
);

NAND2x1p5_ASAP7_75t_L g1225 ( 
.A(n_1081),
.B(n_1198),
.Y(n_1225)
);

AO31x2_ASAP7_75t_L g1226 ( 
.A1(n_1106),
.A2(n_1160),
.A3(n_1098),
.B(n_1195),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_1097),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1140),
.A2(n_1186),
.B1(n_1083),
.B2(n_1184),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1147),
.B(n_1172),
.Y(n_1229)
);

OAI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1094),
.A2(n_1173),
.B1(n_1175),
.B2(n_1197),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1146),
.A2(n_1157),
.B(n_1083),
.Y(n_1231)
);

HB1xp67_ASAP7_75t_L g1232 ( 
.A(n_1097),
.Y(n_1232)
);

AO21x2_ASAP7_75t_L g1233 ( 
.A1(n_1101),
.A2(n_1128),
.B(n_1092),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1085),
.B(n_1093),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1170),
.A2(n_1082),
.B(n_1139),
.C(n_1201),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_1102),
.Y(n_1236)
);

BUFx3_ASAP7_75t_L g1237 ( 
.A(n_1103),
.Y(n_1237)
);

BUFx2_ASAP7_75t_SL g1238 ( 
.A(n_1154),
.Y(n_1238)
);

CKINVDCx16_ASAP7_75t_R g1239 ( 
.A(n_1154),
.Y(n_1239)
);

NAND3xp33_ASAP7_75t_L g1240 ( 
.A(n_1073),
.B(n_1168),
.C(n_1072),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1091),
.B(n_1198),
.Y(n_1241)
);

A2O1A1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1120),
.A2(n_1187),
.B(n_1181),
.C(n_1072),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1148),
.Y(n_1243)
);

OR2x6_ASAP7_75t_L g1244 ( 
.A(n_1070),
.B(n_1125),
.Y(n_1244)
);

OR2x6_ASAP7_75t_L g1245 ( 
.A(n_1070),
.B(n_1112),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1159),
.B(n_1188),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1202),
.A2(n_1117),
.B1(n_1118),
.B2(n_1190),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1155),
.A2(n_1199),
.B(n_1134),
.Y(n_1248)
);

AOI221x1_ASAP7_75t_L g1249 ( 
.A1(n_1116),
.A2(n_1110),
.B1(n_1099),
.B2(n_1124),
.C(n_1129),
.Y(n_1249)
);

HB1xp67_ASAP7_75t_L g1250 ( 
.A(n_1164),
.Y(n_1250)
);

AOI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1135),
.A2(n_1133),
.B(n_1112),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1155),
.A2(n_1199),
.B(n_1132),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1178),
.B(n_1108),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1187),
.A2(n_1183),
.B(n_1179),
.C(n_1164),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1202),
.A2(n_1119),
.B1(n_1187),
.B2(n_1122),
.Y(n_1255)
);

BUFx2_ASAP7_75t_R g1256 ( 
.A(n_1127),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1202),
.B(n_1164),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1202),
.B(n_1179),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1179),
.B(n_1183),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1130),
.A2(n_1123),
.B(n_1193),
.Y(n_1260)
);

INVx6_ASAP7_75t_L g1261 ( 
.A(n_1192),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1126),
.Y(n_1262)
);

AOI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1126),
.A2(n_1112),
.B1(n_1191),
.B2(n_1088),
.Y(n_1263)
);

NOR2x1_ASAP7_75t_L g1264 ( 
.A(n_1126),
.B(n_1088),
.Y(n_1264)
);

OA21x2_ASAP7_75t_L g1265 ( 
.A1(n_1138),
.A2(n_1183),
.B(n_1089),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1089),
.A2(n_1070),
.B(n_1079),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1089),
.B(n_1131),
.Y(n_1267)
);

OAI22x1_ASAP7_75t_L g1268 ( 
.A1(n_1096),
.A2(n_1094),
.B1(n_858),
.B2(n_1105),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1121),
.A2(n_1075),
.B(n_1143),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1121),
.A2(n_1075),
.B(n_1143),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1167),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1111),
.Y(n_1272)
);

NAND2x1_ASAP7_75t_L g1273 ( 
.A(n_1144),
.B(n_1196),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1141),
.A2(n_1162),
.B(n_1161),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1069),
.Y(n_1275)
);

INVx1_ASAP7_75t_SL g1276 ( 
.A(n_1103),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1150),
.B(n_1185),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1076),
.B(n_1142),
.Y(n_1278)
);

NAND2x1p5_ASAP7_75t_L g1279 ( 
.A(n_1081),
.B(n_962),
.Y(n_1279)
);

O2A1O1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_1150),
.A2(n_1185),
.B(n_1158),
.C(n_1180),
.Y(n_1280)
);

OAI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1150),
.A2(n_1185),
.B(n_1158),
.Y(n_1281)
);

INVx4_ASAP7_75t_L g1282 ( 
.A(n_1153),
.Y(n_1282)
);

CKINVDCx20_ASAP7_75t_R g1283 ( 
.A(n_1153),
.Y(n_1283)
);

NAND3xp33_ASAP7_75t_L g1284 ( 
.A(n_1087),
.B(n_858),
.C(n_1150),
.Y(n_1284)
);

OR2x6_ASAP7_75t_L g1285 ( 
.A(n_1090),
.B(n_1070),
.Y(n_1285)
);

INVx4_ASAP7_75t_SL g1286 ( 
.A(n_1202),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_1150),
.B(n_1185),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1167),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1150),
.A2(n_1185),
.B(n_1158),
.Y(n_1289)
);

INVx8_ASAP7_75t_L g1290 ( 
.A(n_1070),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1076),
.B(n_1142),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1150),
.A2(n_1185),
.B(n_1158),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1141),
.A2(n_1162),
.B(n_1161),
.Y(n_1293)
);

INVxp67_ASAP7_75t_L g1294 ( 
.A(n_1100),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1111),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1111),
.Y(n_1296)
);

CKINVDCx20_ASAP7_75t_R g1297 ( 
.A(n_1153),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1075),
.A2(n_1149),
.B(n_1143),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1150),
.A2(n_1185),
.B1(n_885),
.B2(n_858),
.Y(n_1299)
);

INVx1_ASAP7_75t_SL g1300 ( 
.A(n_1103),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1153),
.Y(n_1301)
);

CKINVDCx11_ASAP7_75t_R g1302 ( 
.A(n_1154),
.Y(n_1302)
);

AOI22x1_ASAP7_75t_L g1303 ( 
.A1(n_1170),
.A2(n_488),
.B1(n_528),
.B2(n_1144),
.Y(n_1303)
);

BUFx12f_ASAP7_75t_L g1304 ( 
.A(n_1102),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1141),
.A2(n_1162),
.B(n_1161),
.Y(n_1305)
);

INVx1_ASAP7_75t_SL g1306 ( 
.A(n_1103),
.Y(n_1306)
);

CKINVDCx6p67_ASAP7_75t_R g1307 ( 
.A(n_1154),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1069),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1069),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1069),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_SL g1311 ( 
.A1(n_1150),
.A2(n_1185),
.B1(n_743),
.B2(n_1098),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1069),
.Y(n_1312)
);

A2O1A1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1158),
.A2(n_858),
.B(n_885),
.C(n_1150),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1097),
.Y(n_1314)
);

O2A1O1Ixp33_ASAP7_75t_SL g1315 ( 
.A1(n_1151),
.A2(n_1195),
.B(n_1180),
.C(n_1185),
.Y(n_1315)
);

AO31x2_ASAP7_75t_L g1316 ( 
.A1(n_1077),
.A2(n_1137),
.A3(n_1080),
.B(n_1037),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1150),
.B(n_1185),
.Y(n_1317)
);

CKINVDCx6p67_ASAP7_75t_R g1318 ( 
.A(n_1154),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1092),
.B(n_1085),
.Y(n_1319)
);

CKINVDCx20_ASAP7_75t_R g1320 ( 
.A(n_1236),
.Y(n_1320)
);

CKINVDCx6p67_ASAP7_75t_R g1321 ( 
.A(n_1283),
.Y(n_1321)
);

CKINVDCx6p67_ASAP7_75t_R g1322 ( 
.A(n_1297),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1205),
.B(n_1277),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_SL g1324 ( 
.A1(n_1313),
.A2(n_1280),
.B(n_1281),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1205),
.B(n_1277),
.Y(n_1325)
);

O2A1O1Ixp5_ASAP7_75t_L g1326 ( 
.A1(n_1287),
.A2(n_1317),
.B(n_1289),
.C(n_1292),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1233),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1299),
.A2(n_1287),
.B1(n_1317),
.B2(n_1284),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1299),
.A2(n_1311),
.B1(n_1313),
.B2(n_1216),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_SL g1330 ( 
.A1(n_1280),
.A2(n_1235),
.B(n_1228),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1233),
.Y(n_1331)
);

O2A1O1Ixp5_ASAP7_75t_L g1332 ( 
.A1(n_1231),
.A2(n_1224),
.B(n_1219),
.C(n_1273),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1230),
.B(n_1294),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1209),
.Y(n_1334)
);

O2A1O1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1315),
.A2(n_1235),
.B(n_1207),
.C(n_1230),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1271),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1278),
.B(n_1291),
.Y(n_1337)
);

A2O1A1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1311),
.A2(n_1242),
.B(n_1219),
.C(n_1240),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1319),
.B(n_1272),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_SL g1340 ( 
.A1(n_1242),
.A2(n_1268),
.B(n_1249),
.Y(n_1340)
);

OAI211xp5_ASAP7_75t_L g1341 ( 
.A1(n_1315),
.A2(n_1303),
.B(n_1247),
.C(n_1215),
.Y(n_1341)
);

A2O1A1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1254),
.A2(n_1247),
.B(n_1258),
.C(n_1257),
.Y(n_1342)
);

O2A1O1Ixp33_ASAP7_75t_L g1343 ( 
.A1(n_1210),
.A2(n_1211),
.B(n_1253),
.C(n_1254),
.Y(n_1343)
);

INVxp33_ASAP7_75t_L g1344 ( 
.A(n_1253),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_1286),
.B(n_1285),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1295),
.B(n_1296),
.Y(n_1346)
);

O2A1O1Ixp5_ASAP7_75t_L g1347 ( 
.A1(n_1267),
.A2(n_1251),
.B(n_1259),
.C(n_1258),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1237),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1220),
.B(n_1221),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_1302),
.Y(n_1350)
);

NOR2xp67_ASAP7_75t_L g1351 ( 
.A(n_1282),
.B(n_1217),
.Y(n_1351)
);

O2A1O1Ixp5_ASAP7_75t_L g1352 ( 
.A1(n_1259),
.A2(n_1257),
.B(n_1293),
.C(n_1206),
.Y(n_1352)
);

AOI221x1_ASAP7_75t_SL g1353 ( 
.A1(n_1243),
.A2(n_1246),
.B1(n_1226),
.B2(n_1211),
.C(n_1215),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1276),
.B(n_1300),
.Y(n_1354)
);

A2O1A1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1255),
.A2(n_1250),
.B(n_1222),
.C(n_1226),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1306),
.B(n_1226),
.Y(n_1356)
);

A2O1A1Ixp33_ASAP7_75t_L g1357 ( 
.A1(n_1255),
.A2(n_1250),
.B(n_1226),
.C(n_1293),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1239),
.B(n_1238),
.Y(n_1358)
);

O2A1O1Ixp5_ASAP7_75t_L g1359 ( 
.A1(n_1206),
.A2(n_1208),
.B(n_1241),
.C(n_1282),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1262),
.B(n_1244),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1244),
.B(n_1256),
.Y(n_1361)
);

CKINVDCx16_ASAP7_75t_R g1362 ( 
.A(n_1304),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1256),
.B(n_1288),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1285),
.A2(n_1307),
.B1(n_1318),
.B2(n_1263),
.Y(n_1364)
);

INVx2_ASAP7_75t_SL g1365 ( 
.A(n_1261),
.Y(n_1365)
);

O2A1O1Ixp5_ASAP7_75t_L g1366 ( 
.A1(n_1208),
.A2(n_1241),
.B(n_1314),
.C(n_1232),
.Y(n_1366)
);

O2A1O1Ixp5_ASAP7_75t_L g1367 ( 
.A1(n_1227),
.A2(n_1232),
.B(n_1314),
.C(n_1316),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1285),
.A2(n_1213),
.B1(n_1264),
.B2(n_1261),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1261),
.A2(n_1245),
.B1(n_1223),
.B2(n_1265),
.Y(n_1369)
);

AOI221x1_ASAP7_75t_SL g1370 ( 
.A1(n_1316),
.A2(n_1312),
.B1(n_1308),
.B2(n_1275),
.C(n_1309),
.Y(n_1370)
);

O2A1O1Ixp5_ASAP7_75t_L g1371 ( 
.A1(n_1316),
.A2(n_1310),
.B(n_1248),
.C(n_1286),
.Y(n_1371)
);

O2A1O1Ixp5_ASAP7_75t_L g1372 ( 
.A1(n_1286),
.A2(n_1252),
.B(n_1260),
.C(n_1266),
.Y(n_1372)
);

OA21x2_ASAP7_75t_L g1373 ( 
.A1(n_1298),
.A2(n_1218),
.B(n_1270),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1245),
.B(n_1223),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1245),
.A2(n_1301),
.B1(n_1212),
.B2(n_1225),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1269),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1214),
.A2(n_1279),
.B(n_1290),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1290),
.B(n_1279),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1204),
.B(n_1203),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1229),
.B(n_1234),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1233),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1205),
.A2(n_1090),
.B(n_1277),
.Y(n_1382)
);

O2A1O1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1313),
.A2(n_1185),
.B(n_1150),
.C(n_1205),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1205),
.A2(n_1090),
.B(n_1277),
.Y(n_1384)
);

OA21x2_ASAP7_75t_L g1385 ( 
.A1(n_1274),
.A2(n_1305),
.B(n_1293),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1205),
.A2(n_1090),
.B(n_1277),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1204),
.B(n_1203),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_1302),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1299),
.A2(n_1277),
.B1(n_1287),
.B2(n_1205),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1204),
.B(n_1203),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_SL g1391 ( 
.A1(n_1313),
.A2(n_1280),
.B(n_1158),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1204),
.B(n_1203),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1204),
.B(n_1203),
.Y(n_1393)
);

BUFx2_ASAP7_75t_L g1394 ( 
.A(n_1294),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1229),
.B(n_1234),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_1302),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_SL g1397 ( 
.A1(n_1313),
.A2(n_1280),
.B(n_1158),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1299),
.A2(n_1277),
.B1(n_1287),
.B2(n_1205),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1205),
.A2(n_1090),
.B(n_1277),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1299),
.A2(n_1277),
.B1(n_1287),
.B2(n_1205),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1299),
.A2(n_1277),
.B1(n_1287),
.B2(n_1205),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1204),
.B(n_1203),
.Y(n_1402)
);

OR2x6_ASAP7_75t_L g1403 ( 
.A(n_1345),
.B(n_1357),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1334),
.Y(n_1404)
);

OR2x6_ASAP7_75t_L g1405 ( 
.A(n_1345),
.B(n_1357),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1327),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1356),
.B(n_1333),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_1377),
.Y(n_1408)
);

AO21x2_ASAP7_75t_L g1409 ( 
.A1(n_1355),
.A2(n_1331),
.B(n_1381),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1385),
.B(n_1352),
.Y(n_1410)
);

BUFx3_ASAP7_75t_L g1411 ( 
.A(n_1348),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1349),
.Y(n_1412)
);

BUFx3_ASAP7_75t_L g1413 ( 
.A(n_1377),
.Y(n_1413)
);

OA21x2_ASAP7_75t_L g1414 ( 
.A1(n_1367),
.A2(n_1371),
.B(n_1332),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1385),
.B(n_1342),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1373),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1394),
.B(n_1339),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1353),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1385),
.B(n_1342),
.Y(n_1419)
);

AO21x2_ASAP7_75t_L g1420 ( 
.A1(n_1338),
.A2(n_1376),
.B(n_1340),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1347),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1346),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1389),
.A2(n_1401),
.B1(n_1400),
.B2(n_1398),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1323),
.B(n_1325),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1382),
.B(n_1384),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1379),
.B(n_1387),
.Y(n_1426)
);

OR2x6_ASAP7_75t_L g1427 ( 
.A(n_1324),
.B(n_1369),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1390),
.B(n_1402),
.Y(n_1428)
);

AO21x2_ASAP7_75t_L g1429 ( 
.A1(n_1338),
.A2(n_1399),
.B(n_1386),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1372),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1370),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1366),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1392),
.B(n_1393),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1328),
.B(n_1330),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1343),
.Y(n_1435)
);

AO21x2_ASAP7_75t_L g1436 ( 
.A1(n_1341),
.A2(n_1397),
.B(n_1391),
.Y(n_1436)
);

AO21x2_ASAP7_75t_L g1437 ( 
.A1(n_1329),
.A2(n_1335),
.B(n_1383),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1337),
.B(n_1344),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1344),
.B(n_1326),
.Y(n_1439)
);

AND2x4_ASAP7_75t_L g1440 ( 
.A(n_1413),
.B(n_1415),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1437),
.A2(n_1380),
.B1(n_1395),
.B2(n_1361),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1406),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1416),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1415),
.B(n_1354),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1415),
.B(n_1336),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1404),
.Y(n_1446)
);

AO21x2_ASAP7_75t_L g1447 ( 
.A1(n_1418),
.A2(n_1368),
.B(n_1360),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1418),
.B(n_1336),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1437),
.A2(n_1363),
.B1(n_1374),
.B2(n_1322),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1406),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1437),
.A2(n_1374),
.B1(n_1321),
.B2(n_1322),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1419),
.B(n_1410),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1419),
.B(n_1359),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1439),
.B(n_1358),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1421),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_1408),
.Y(n_1456)
);

AOI221xp5_ASAP7_75t_L g1457 ( 
.A1(n_1423),
.A2(n_1364),
.B1(n_1375),
.B2(n_1358),
.C(n_1388),
.Y(n_1457)
);

INVx1_ASAP7_75t_SL g1458 ( 
.A(n_1408),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1416),
.Y(n_1459)
);

AOI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1425),
.A2(n_1378),
.B(n_1365),
.Y(n_1460)
);

INVxp67_ASAP7_75t_L g1461 ( 
.A(n_1439),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1416),
.Y(n_1462)
);

OAI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1461),
.A2(n_1427),
.B1(n_1425),
.B2(n_1434),
.Y(n_1463)
);

BUFx3_ASAP7_75t_L g1464 ( 
.A(n_1448),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1446),
.Y(n_1465)
);

INVx1_ASAP7_75t_SL g1466 ( 
.A(n_1445),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_SL g1467 ( 
.A(n_1445),
.B(n_1439),
.Y(n_1467)
);

OAI31xp33_ASAP7_75t_L g1468 ( 
.A1(n_1441),
.A2(n_1434),
.A3(n_1423),
.B(n_1435),
.Y(n_1468)
);

BUFx2_ASAP7_75t_L g1469 ( 
.A(n_1453),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1455),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_SL g1471 ( 
.A(n_1445),
.B(n_1424),
.Y(n_1471)
);

AOI221xp5_ASAP7_75t_L g1472 ( 
.A1(n_1441),
.A2(n_1431),
.B1(n_1461),
.B2(n_1435),
.C(n_1455),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_R g1473 ( 
.A(n_1448),
.B(n_1320),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1452),
.B(n_1421),
.Y(n_1474)
);

AOI33xp33_ASAP7_75t_L g1475 ( 
.A1(n_1452),
.A2(n_1431),
.A3(n_1438),
.B1(n_1412),
.B2(n_1428),
.B3(n_1426),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_SL g1476 ( 
.A1(n_1440),
.A2(n_1437),
.B1(n_1429),
.B2(n_1436),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1442),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1444),
.B(n_1424),
.Y(n_1478)
);

OAI211xp5_ASAP7_75t_L g1479 ( 
.A1(n_1457),
.A2(n_1408),
.B(n_1414),
.C(n_1411),
.Y(n_1479)
);

INVx3_ASAP7_75t_L g1480 ( 
.A(n_1456),
.Y(n_1480)
);

AOI221xp5_ASAP7_75t_L g1481 ( 
.A1(n_1452),
.A2(n_1437),
.B1(n_1432),
.B2(n_1422),
.C(n_1407),
.Y(n_1481)
);

NAND4xp25_ASAP7_75t_SL g1482 ( 
.A(n_1457),
.B(n_1433),
.C(n_1426),
.D(n_1428),
.Y(n_1482)
);

OAI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1457),
.A2(n_1427),
.B1(n_1405),
.B2(n_1403),
.Y(n_1483)
);

OAI211xp5_ASAP7_75t_L g1484 ( 
.A1(n_1448),
.A2(n_1414),
.B(n_1411),
.C(n_1430),
.Y(n_1484)
);

OAI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1454),
.A2(n_1427),
.B1(n_1405),
.B2(n_1403),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1440),
.A2(n_1436),
.B1(n_1429),
.B2(n_1420),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1440),
.A2(n_1436),
.B1(n_1429),
.B2(n_1420),
.Y(n_1487)
);

AO21x2_ASAP7_75t_L g1488 ( 
.A1(n_1447),
.A2(n_1430),
.B(n_1432),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1451),
.A2(n_1427),
.B1(n_1433),
.B2(n_1403),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_SL g1490 ( 
.A1(n_1440),
.A2(n_1429),
.B1(n_1436),
.B2(n_1420),
.Y(n_1490)
);

OAI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1454),
.A2(n_1427),
.B1(n_1405),
.B2(n_1403),
.Y(n_1491)
);

OAI221xp5_ASAP7_75t_SL g1492 ( 
.A1(n_1452),
.A2(n_1427),
.B1(n_1407),
.B2(n_1403),
.C(n_1405),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1449),
.A2(n_1427),
.B1(n_1433),
.B2(n_1405),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1454),
.B(n_1417),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1442),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1440),
.A2(n_1436),
.B1(n_1429),
.B2(n_1420),
.Y(n_1496)
);

INVxp67_ASAP7_75t_SL g1497 ( 
.A(n_1453),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1469),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1465),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1465),
.Y(n_1500)
);

OAI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1468),
.A2(n_1460),
.B(n_1449),
.Y(n_1501)
);

NAND3xp33_ASAP7_75t_SL g1502 ( 
.A(n_1468),
.B(n_1458),
.C(n_1460),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1470),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1477),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1475),
.B(n_1444),
.Y(n_1505)
);

INVxp67_ASAP7_75t_L g1506 ( 
.A(n_1464),
.Y(n_1506)
);

OA21x2_ASAP7_75t_L g1507 ( 
.A1(n_1479),
.A2(n_1462),
.B(n_1459),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1495),
.Y(n_1508)
);

BUFx2_ASAP7_75t_L g1509 ( 
.A(n_1469),
.Y(n_1509)
);

AOI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1483),
.A2(n_1460),
.B(n_1405),
.Y(n_1510)
);

OAI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1486),
.A2(n_1443),
.B(n_1459),
.Y(n_1511)
);

OA21x2_ASAP7_75t_L g1512 ( 
.A1(n_1484),
.A2(n_1462),
.B(n_1459),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1497),
.B(n_1453),
.Y(n_1513)
);

INVx4_ASAP7_75t_SL g1514 ( 
.A(n_1464),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1474),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1481),
.B(n_1444),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_1488),
.Y(n_1517)
);

AO21x2_ASAP7_75t_L g1518 ( 
.A1(n_1488),
.A2(n_1409),
.B(n_1447),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1474),
.B(n_1450),
.Y(n_1519)
);

AND2x4_ASAP7_75t_L g1520 ( 
.A(n_1480),
.B(n_1440),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1494),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1499),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1499),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1499),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1521),
.B(n_1478),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1518),
.Y(n_1526)
);

OAI221xp5_ASAP7_75t_L g1527 ( 
.A1(n_1501),
.A2(n_1476),
.B1(n_1472),
.B2(n_1490),
.C(n_1496),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1498),
.Y(n_1528)
);

NOR2xp67_ASAP7_75t_L g1529 ( 
.A(n_1502),
.B(n_1482),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1513),
.B(n_1466),
.Y(n_1530)
);

AOI211xp5_ASAP7_75t_SL g1531 ( 
.A1(n_1502),
.A2(n_1463),
.B(n_1492),
.C(n_1491),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1516),
.A2(n_1487),
.B1(n_1440),
.B2(n_1447),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1500),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1500),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_1506),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_1498),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1513),
.B(n_1473),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1521),
.B(n_1494),
.Y(n_1538)
);

AOI211xp5_ASAP7_75t_SL g1539 ( 
.A1(n_1510),
.A2(n_1485),
.B(n_1493),
.C(n_1489),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1514),
.B(n_1467),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1498),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1505),
.B(n_1417),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1514),
.B(n_1471),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1500),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1506),
.B(n_1350),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1514),
.B(n_1456),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1509),
.Y(n_1547)
);

INVx1_ASAP7_75t_SL g1548 ( 
.A(n_1509),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1507),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1507),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1514),
.B(n_1445),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1505),
.B(n_1417),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1518),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1519),
.B(n_1516),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1549),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1522),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1529),
.B(n_1509),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1522),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1549),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1537),
.B(n_1514),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1549),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1523),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1527),
.A2(n_1501),
.B1(n_1517),
.B2(n_1507),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1523),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1537),
.B(n_1515),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1554),
.B(n_1519),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1529),
.B(n_1525),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1524),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1533),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1543),
.B(n_1520),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1525),
.B(n_1503),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1533),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1554),
.B(n_1519),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1535),
.B(n_1504),
.Y(n_1574)
);

INVx2_ASAP7_75t_SL g1575 ( 
.A(n_1528),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1534),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1543),
.B(n_1551),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1534),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1549),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1540),
.B(n_1546),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1548),
.B(n_1504),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1538),
.B(n_1508),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1544),
.Y(n_1583)
);

INVxp67_ASAP7_75t_L g1584 ( 
.A(n_1545),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1550),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1538),
.B(n_1548),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1528),
.Y(n_1587)
);

AOI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1563),
.A2(n_1527),
.B(n_1557),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1566),
.B(n_1542),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1587),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1580),
.B(n_1536),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1567),
.B(n_1536),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1557),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1567),
.B(n_1541),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1556),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1560),
.B(n_1530),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1556),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1560),
.B(n_1530),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1557),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1566),
.B(n_1542),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1573),
.B(n_1552),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1573),
.B(n_1552),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1558),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1565),
.B(n_1541),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1580),
.B(n_1546),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1577),
.B(n_1546),
.Y(n_1606)
);

INVx3_ASAP7_75t_L g1607 ( 
.A(n_1557),
.Y(n_1607)
);

CKINVDCx16_ASAP7_75t_R g1608 ( 
.A(n_1574),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1558),
.Y(n_1609)
);

BUFx3_ASAP7_75t_L g1610 ( 
.A(n_1575),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1562),
.Y(n_1611)
);

CKINVDCx6p67_ASAP7_75t_R g1612 ( 
.A(n_1586),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1555),
.Y(n_1613)
);

INVxp67_ASAP7_75t_L g1614 ( 
.A(n_1607),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1588),
.A2(n_1532),
.B1(n_1507),
.B2(n_1550),
.Y(n_1615)
);

AO211x2_ASAP7_75t_L g1616 ( 
.A1(n_1592),
.A2(n_1586),
.B(n_1510),
.C(n_1531),
.Y(n_1616)
);

INVxp67_ASAP7_75t_L g1617 ( 
.A(n_1607),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1595),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1595),
.Y(n_1619)
);

AOI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1608),
.A2(n_1507),
.B1(n_1550),
.B2(n_1518),
.Y(n_1620)
);

INVx1_ASAP7_75t_SL g1621 ( 
.A(n_1612),
.Y(n_1621)
);

AOI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1608),
.A2(n_1507),
.B1(n_1550),
.B2(n_1518),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1597),
.Y(n_1623)
);

O2A1O1Ixp33_ASAP7_75t_SL g1624 ( 
.A1(n_1604),
.A2(n_1584),
.B(n_1571),
.C(n_1547),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1596),
.B(n_1565),
.Y(n_1625)
);

OAI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1594),
.A2(n_1531),
.B(n_1539),
.Y(n_1626)
);

A2O1A1Ixp33_ASAP7_75t_L g1627 ( 
.A1(n_1589),
.A2(n_1539),
.B(n_1511),
.C(n_1517),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1612),
.B(n_1575),
.Y(n_1628)
);

OAI322xp33_ASAP7_75t_L g1629 ( 
.A1(n_1590),
.A2(n_1582),
.A3(n_1571),
.B1(n_1581),
.B2(n_1559),
.C1(n_1555),
.C2(n_1561),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1597),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_SL g1631 ( 
.A1(n_1593),
.A2(n_1512),
.B(n_1396),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1590),
.B(n_1582),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1625),
.B(n_1610),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1627),
.A2(n_1626),
.B1(n_1615),
.B2(n_1620),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1621),
.B(n_1607),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1618),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1619),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1628),
.B(n_1593),
.Y(n_1638)
);

INVxp67_ASAP7_75t_L g1639 ( 
.A(n_1632),
.Y(n_1639)
);

INVx3_ASAP7_75t_L g1640 ( 
.A(n_1623),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1630),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1624),
.B(n_1599),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1614),
.B(n_1610),
.Y(n_1643)
);

A2O1A1Ixp33_ASAP7_75t_L g1644 ( 
.A1(n_1634),
.A2(n_1622),
.B(n_1616),
.C(n_1632),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1639),
.B(n_1617),
.Y(n_1645)
);

NOR2x1_ASAP7_75t_L g1646 ( 
.A(n_1640),
.B(n_1599),
.Y(n_1646)
);

AOI221xp5_ASAP7_75t_L g1647 ( 
.A1(n_1642),
.A2(n_1629),
.B1(n_1631),
.B2(n_1638),
.C(n_1641),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1635),
.B(n_1596),
.Y(n_1648)
);

AOI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1633),
.A2(n_1598),
.B1(n_1613),
.B2(n_1606),
.Y(n_1649)
);

AOI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1643),
.A2(n_1598),
.B1(n_1613),
.B2(n_1606),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1640),
.A2(n_1591),
.B(n_1547),
.Y(n_1651)
);

AOI211xp5_ASAP7_75t_L g1652 ( 
.A1(n_1636),
.A2(n_1611),
.B(n_1603),
.C(n_1609),
.Y(n_1652)
);

NAND3xp33_ASAP7_75t_L g1653 ( 
.A(n_1637),
.B(n_1591),
.C(n_1603),
.Y(n_1653)
);

OAI21xp33_ASAP7_75t_L g1654 ( 
.A1(n_1648),
.A2(n_1591),
.B(n_1605),
.Y(n_1654)
);

OAI211xp5_ASAP7_75t_L g1655 ( 
.A1(n_1647),
.A2(n_1611),
.B(n_1609),
.C(n_1605),
.Y(n_1655)
);

OAI22xp5_ASAP7_75t_L g1656 ( 
.A1(n_1649),
.A2(n_1644),
.B1(n_1650),
.B2(n_1601),
.Y(n_1656)
);

OAI221xp5_ASAP7_75t_SL g1657 ( 
.A1(n_1645),
.A2(n_1602),
.B1(n_1589),
.B2(n_1601),
.C(n_1600),
.Y(n_1657)
);

OAI21xp5_ASAP7_75t_L g1658 ( 
.A1(n_1651),
.A2(n_1591),
.B(n_1602),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1658),
.Y(n_1659)
);

NOR2x1_ASAP7_75t_L g1660 ( 
.A(n_1656),
.B(n_1646),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1657),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1654),
.B(n_1577),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1655),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1658),
.Y(n_1664)
);

NOR2x1_ASAP7_75t_L g1665 ( 
.A(n_1660),
.B(n_1653),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_R g1666 ( 
.A(n_1659),
.B(n_1320),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1664),
.Y(n_1667)
);

OAI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1663),
.A2(n_1600),
.B1(n_1652),
.B2(n_1585),
.Y(n_1668)
);

INVx2_ASAP7_75t_SL g1669 ( 
.A(n_1662),
.Y(n_1669)
);

OAI211xp5_ASAP7_75t_L g1670 ( 
.A1(n_1665),
.A2(n_1661),
.B(n_1555),
.C(n_1585),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1667),
.Y(n_1671)
);

NOR3xp33_ASAP7_75t_L g1672 ( 
.A(n_1668),
.B(n_1661),
.C(n_1362),
.Y(n_1672)
);

NAND4xp75_ASAP7_75t_L g1673 ( 
.A(n_1671),
.B(n_1669),
.C(n_1666),
.D(n_1559),
.Y(n_1673)
);

AOI322xp5_ASAP7_75t_L g1674 ( 
.A1(n_1673),
.A2(n_1672),
.A3(n_1670),
.B1(n_1585),
.B2(n_1579),
.C1(n_1561),
.C2(n_1559),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1674),
.B(n_1570),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1674),
.Y(n_1676)
);

OAI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1676),
.A2(n_1561),
.B1(n_1579),
.B2(n_1583),
.Y(n_1677)
);

OAI22x1_ASAP7_75t_L g1678 ( 
.A1(n_1675),
.A2(n_1583),
.B1(n_1562),
.B2(n_1564),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1677),
.A2(n_1579),
.B1(n_1526),
.B2(n_1553),
.Y(n_1679)
);

CKINVDCx20_ASAP7_75t_R g1680 ( 
.A(n_1678),
.Y(n_1680)
);

CKINVDCx20_ASAP7_75t_R g1681 ( 
.A(n_1680),
.Y(n_1681)
);

NAND3xp33_ASAP7_75t_L g1682 ( 
.A(n_1681),
.B(n_1679),
.C(n_1568),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1682),
.B(n_1321),
.Y(n_1683)
);

OAI211xp5_ASAP7_75t_L g1684 ( 
.A1(n_1683),
.A2(n_1564),
.B(n_1578),
.C(n_1576),
.Y(n_1684)
);

AOI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1684),
.A2(n_1568),
.B1(n_1578),
.B2(n_1576),
.Y(n_1685)
);

AOI211xp5_ASAP7_75t_L g1686 ( 
.A1(n_1685),
.A2(n_1351),
.B(n_1572),
.C(n_1569),
.Y(n_1686)
);


endmodule