module fake_jpeg_28838_n_139 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_139);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_39),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_12),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_11),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_64),
.Y(n_78)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_65),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_53),
.Y(n_69)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_65),
.A2(n_46),
.B1(n_55),
.B2(n_48),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_75),
.B1(n_1),
.B2(n_2),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_72),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_62),
.B(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_71),
.B(n_77),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_46),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_54),
.B1(n_49),
.B2(n_45),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_74),
.A2(n_76),
.B1(n_3),
.B2(n_4),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_65),
.A2(n_53),
.B1(n_52),
.B2(n_42),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_44),
.B1(n_47),
.B2(n_19),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_0),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_86),
.Y(n_94)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_82),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_1),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_2),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_89),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_90),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_3),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_75),
.B(n_21),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_73),
.A2(n_22),
.B1(n_36),
.B2(n_35),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_92),
.A2(n_17),
.B1(n_32),
.B2(n_30),
.Y(n_99)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_13),
.Y(n_102)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_18),
.C(n_41),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_96),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_91),
.B(n_4),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_73),
.B1(n_6),
.B2(n_7),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_26),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_5),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_108),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_82),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_90),
.C(n_93),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_5),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_110),
.B(n_112),
.Y(n_125)
);

OA21x2_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_83),
.B(n_92),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_113),
.B(n_119),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_6),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_98),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_115),
.A2(n_112),
.B1(n_110),
.B2(n_118),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_95),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_121),
.B(n_101),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_14),
.C(n_23),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_106),
.A2(n_9),
.B(n_10),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_123),
.B(n_127),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_130),
.Y(n_132)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_122),
.C(n_120),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_131),
.A2(n_126),
.B1(n_106),
.B2(n_101),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_132),
.B(n_107),
.Y(n_134)
);

NOR2xp67_ASAP7_75t_SL g135 ( 
.A(n_134),
.B(n_111),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_116),
.Y(n_136)
);

NOR3xp33_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_10),
.C(n_25),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_29),
.B(n_34),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_100),
.Y(n_139)
);


endmodule