module fake_jpeg_22904_n_253 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_253);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_253;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_24),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_38),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_37),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_1),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_43),
.Y(n_51)
);

INVx2_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_26),
.B(n_1),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_42),
.Y(n_60)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_50),
.Y(n_72)
);

OR2x4_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_20),
.Y(n_49)
);

NAND3xp33_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_61),
.C(n_51),
.Y(n_86)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_67),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_46),
.B(n_29),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_53),
.B(n_23),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_21),
.B1(n_17),
.B2(n_18),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_56),
.A2(n_64),
.B1(n_22),
.B2(n_31),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_35),
.B1(n_17),
.B2(n_21),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_59),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_60),
.B(n_26),
.Y(n_77)
);

CKINVDCx12_ASAP7_75t_R g62 ( 
.A(n_36),
.Y(n_62)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_17),
.B1(n_30),
.B2(n_35),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_28),
.Y(n_66)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

CKINVDCx12_ASAP7_75t_R g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_18),
.B1(n_20),
.B2(n_31),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_71),
.A2(n_88),
.B1(n_69),
.B2(n_31),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_51),
.C(n_56),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_74),
.B(n_27),
.C(n_3),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_77),
.B(n_83),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_45),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_87),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_31),
.B1(n_22),
.B2(n_44),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_82),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_30),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_84),
.B(n_90),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_86),
.A2(n_102),
.B1(n_34),
.B2(n_32),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_61),
.B(n_23),
.Y(n_87)
);

OA22x2_ASAP7_75t_SL g88 ( 
.A1(n_48),
.A2(n_31),
.B1(n_22),
.B2(n_45),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_24),
.Y(n_89)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_93),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_24),
.Y(n_92)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_57),
.B(n_33),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_97),
.B(n_34),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_19),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_100),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_57),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_45),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_24),
.Y(n_123)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_24),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_75),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_104),
.B(n_117),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_129),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_96),
.A2(n_65),
.B1(n_29),
.B2(n_32),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_106),
.A2(n_108),
.B1(n_112),
.B2(n_115),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_96),
.A2(n_65),
.B1(n_33),
.B2(n_25),
.Y(n_108)
);

MAJx2_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_35),
.C(n_19),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_126),
.C(n_87),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_L g112 ( 
.A1(n_88),
.A2(n_59),
.B1(n_30),
.B2(n_35),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_113),
.B(n_97),
.Y(n_148)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_28),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_83),
.B(n_78),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_71),
.Y(n_139)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_79),
.B(n_27),
.Y(n_127)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_128),
.A2(n_78),
.B(n_90),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_140),
.B(n_143),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_116),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_136),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_113),
.B(n_77),
.Y(n_136)
);

AND2x6_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_74),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_SL g175 ( 
.A(n_137),
.B(n_119),
.C(n_73),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_150),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_102),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_141),
.A2(n_145),
.B(n_114),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_82),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_151),
.C(n_129),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_101),
.Y(n_143)
);

XNOR2x2_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_83),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_110),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_148),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_72),
.Y(n_147)
);

BUFx24_ASAP7_75t_SL g159 ( 
.A(n_147),
.Y(n_159)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_152),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_76),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_114),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_109),
.B(n_79),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_155),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_76),
.Y(n_155)
);

CKINVDCx12_ASAP7_75t_R g156 ( 
.A(n_124),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_165),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_144),
.A2(n_117),
.B1(n_112),
.B2(n_106),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_158),
.B(n_178),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_164),
.B(n_160),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_145),
.A2(n_122),
.B(n_105),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_177),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_174),
.C(n_150),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_107),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_170),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_134),
.A2(n_122),
.B1(n_118),
.B2(n_108),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_171),
.A2(n_141),
.B(n_147),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_85),
.B1(n_93),
.B2(n_91),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_172),
.A2(n_179),
.B1(n_98),
.B2(n_133),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_118),
.C(n_84),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_180),
.Y(n_183)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_135),
.A2(n_85),
.B1(n_103),
.B2(n_94),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_190),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_143),
.Y(n_185)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_186),
.B(n_195),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_196),
.C(n_169),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_189),
.A2(n_192),
.B1(n_193),
.B2(n_198),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_143),
.Y(n_190)
);

MAJx2_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_197),
.C(n_176),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_180),
.A2(n_134),
.B1(n_140),
.B2(n_137),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_151),
.C(n_139),
.Y(n_196)
);

AOI322xp5_ASAP7_75t_L g197 ( 
.A1(n_164),
.A2(n_140),
.A3(n_119),
.B1(n_138),
.B2(n_73),
.C1(n_16),
.C2(n_15),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_L g198 ( 
.A1(n_167),
.A2(n_73),
.B1(n_3),
.B2(n_4),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_163),
.B(n_16),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_199),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_183),
.A2(n_178),
.B1(n_160),
.B2(n_179),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_200),
.A2(n_209),
.B1(n_181),
.B2(n_192),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_183),
.A2(n_162),
.B(n_175),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_201),
.A2(n_206),
.B(n_210),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_207),
.C(n_212),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_205),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_188),
.A2(n_157),
.B(n_174),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_173),
.C(n_168),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_193),
.A2(n_171),
.B1(n_159),
.B2(n_176),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_15),
.C(n_4),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_14),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_189),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_202),
.A2(n_181),
.B1(n_190),
.B2(n_185),
.Y(n_216)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_216),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_221),
.Y(n_230)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_208),
.B(n_182),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_184),
.C(n_182),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_225),
.C(n_214),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_203),
.A2(n_195),
.B1(n_194),
.B2(n_197),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_223),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_203),
.B(n_199),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_224),
.A2(n_206),
.B(n_212),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_2),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_6),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_226),
.B(n_7),
.Y(n_227)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_227),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_L g228 ( 
.A1(n_220),
.A2(n_200),
.B1(n_211),
.B2(n_201),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_228),
.A2(n_217),
.B1(n_223),
.B2(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_233),
.B(n_225),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_218),
.A2(n_210),
.B(n_209),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_235),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_238),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_216),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_229),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_243),
.A2(n_246),
.B(n_238),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_231),
.Y(n_244)
);

AOI221xp5_ASAP7_75t_L g249 ( 
.A1(n_244),
.A2(n_245),
.B1(n_246),
.B2(n_8),
.C(n_9),
.Y(n_249)
);

AOI31xp67_ASAP7_75t_SL g245 ( 
.A1(n_237),
.A2(n_228),
.A3(n_235),
.B(n_222),
.Y(n_245)
);

A2O1A1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_234),
.B(n_233),
.C(n_215),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_247),
.A2(n_249),
.B1(n_7),
.B2(n_9),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_242),
.A2(n_241),
.B(n_215),
.Y(n_248)
);

AOI322xp5_ASAP7_75t_L g251 ( 
.A1(n_248),
.A2(n_11),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C1(n_236),
.C2(n_242),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_250),
.B(n_251),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_11),
.Y(n_253)
);


endmodule