module fake_aes_5772_n_39 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_39);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_17;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NAND2xp5_ASAP7_75t_L g15 ( .A(n_12), .B(n_8), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_5), .Y(n_16) );
AND2x4_ASAP7_75t_L g17 ( .A(n_3), .B(n_4), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_14), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_1), .B(n_2), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_0), .B(n_5), .Y(n_20) );
CKINVDCx20_ASAP7_75t_R g21 ( .A(n_4), .Y(n_21) );
AOI22xp33_ASAP7_75t_L g22 ( .A1(n_17), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_22) );
BUFx4f_ASAP7_75t_SL g23 ( .A(n_21), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_18), .B(n_3), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
OAI21xp5_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_18), .B(n_15), .Y(n_26) );
INVxp67_ASAP7_75t_SL g27 ( .A(n_25), .Y(n_27) );
OR2x2_ASAP7_75t_L g28 ( .A(n_27), .B(n_25), .Y(n_28) );
AND2x4_ASAP7_75t_L g29 ( .A(n_27), .B(n_21), .Y(n_29) );
OAI22xp5_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_26), .B1(n_22), .B2(n_17), .Y(n_30) );
AOI22xp5_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_23), .B1(n_16), .B2(n_17), .Y(n_31) );
AOI211xp5_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_19), .B(n_16), .C(n_20), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
NOR2x1_ASAP7_75t_L g34 ( .A(n_33), .B(n_6), .Y(n_34) );
AND2x2_ASAP7_75t_L g35 ( .A(n_32), .B(n_7), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_34), .Y(n_36) );
INVx2_ASAP7_75t_L g37 ( .A(n_35), .Y(n_37) );
AOI22xp5_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_38) );
OA22x2_ASAP7_75t_L g39 ( .A1(n_38), .A2(n_37), .B1(n_36), .B2(n_13), .Y(n_39) );
endmodule