module real_aes_6253_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_746;
wire n_153;
wire n_532;
wire n_316;
wire n_284;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_753;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_0), .B(n_109), .C(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g123 ( .A(n_0), .Y(n_123) );
INVx1_ASAP7_75t_L g499 ( .A(n_1), .Y(n_499) );
INVx1_ASAP7_75t_L g213 ( .A(n_2), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g757 ( .A1(n_3), .A2(n_80), .B1(n_758), .B2(n_759), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_3), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_4), .A2(n_39), .B1(n_169), .B2(n_515), .Y(n_525) );
AOI21xp33_ASAP7_75t_L g193 ( .A1(n_5), .A2(n_150), .B(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_6), .B(n_143), .Y(n_490) );
AND2x6_ASAP7_75t_L g155 ( .A(n_7), .B(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_8), .A2(n_252), .B(n_253), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_9), .B(n_107), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_9), .B(n_40), .Y(n_124) );
INVx1_ASAP7_75t_L g200 ( .A(n_10), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_11), .B(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g148 ( .A(n_12), .Y(n_148) );
INVx1_ASAP7_75t_L g494 ( .A(n_13), .Y(n_494) );
INVx1_ASAP7_75t_L g258 ( .A(n_14), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_15), .B(n_181), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_16), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_17), .B(n_144), .Y(n_471) );
AO32x2_ASAP7_75t_L g523 ( .A1(n_18), .A2(n_143), .A3(n_178), .B1(n_477), .B2(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_19), .B(n_169), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_20), .B(n_164), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_21), .B(n_144), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_22), .A2(n_52), .B1(n_169), .B2(n_515), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_23), .B(n_150), .Y(n_224) );
AOI22xp33_ASAP7_75t_SL g521 ( .A1(n_24), .A2(n_77), .B1(n_169), .B2(n_181), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_25), .B(n_169), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_26), .B(n_172), .Y(n_171) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_27), .A2(n_256), .B(n_257), .C(n_259), .Y(n_255) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_28), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_29), .B(n_202), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_30), .B(n_198), .Y(n_215) );
AOI222xp33_ASAP7_75t_SL g126 ( .A1(n_31), .A2(n_127), .B1(n_133), .B2(n_741), .C1(n_742), .C2(n_747), .Y(n_126) );
OAI22xp5_ASAP7_75t_L g128 ( .A1(n_32), .A2(n_43), .B1(n_129), .B2(n_130), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_32), .Y(n_129) );
INVx1_ASAP7_75t_L g187 ( .A(n_33), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_34), .B(n_202), .Y(n_538) );
INVx2_ASAP7_75t_L g153 ( .A(n_35), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_36), .B(n_169), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_37), .B(n_202), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_38), .A2(n_155), .B(n_159), .C(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g107 ( .A(n_40), .Y(n_107) );
INVx1_ASAP7_75t_L g185 ( .A(n_41), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_42), .B(n_198), .Y(n_268) );
CKINVDCx14_ASAP7_75t_R g130 ( .A(n_43), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_44), .B(n_169), .Y(n_484) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_45), .A2(n_128), .B1(n_131), .B2(n_132), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_45), .Y(n_132) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_46), .A2(n_88), .B1(n_231), .B2(n_515), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_47), .B(n_169), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_48), .B(n_169), .Y(n_495) );
CKINVDCx16_ASAP7_75t_R g188 ( .A(n_49), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_50), .B(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_51), .B(n_150), .Y(n_246) );
AOI22xp33_ASAP7_75t_SL g476 ( .A1(n_53), .A2(n_62), .B1(n_169), .B2(n_181), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_54), .A2(n_159), .B1(n_181), .B2(n_183), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_55), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_56), .B(n_169), .Y(n_509) );
CKINVDCx16_ASAP7_75t_R g210 ( .A(n_57), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_58), .B(n_169), .Y(n_558) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_59), .A2(n_168), .B(n_197), .C(n_199), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_60), .Y(n_272) );
INVx1_ASAP7_75t_L g195 ( .A(n_61), .Y(n_195) );
INVx1_ASAP7_75t_L g156 ( .A(n_63), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_64), .B(n_169), .Y(n_500) );
INVx1_ASAP7_75t_L g147 ( .A(n_65), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_66), .Y(n_117) );
AO32x2_ASAP7_75t_L g518 ( .A1(n_67), .A2(n_143), .A3(n_238), .B1(n_477), .B2(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g557 ( .A(n_68), .Y(n_557) );
INVx1_ASAP7_75t_L g533 ( .A(n_69), .Y(n_533) );
A2O1A1Ixp33_ASAP7_75t_SL g163 ( .A1(n_70), .A2(n_164), .B(n_165), .C(n_168), .Y(n_163) );
INVxp67_ASAP7_75t_L g166 ( .A(n_71), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_72), .B(n_181), .Y(n_534) );
INVx1_ASAP7_75t_L g112 ( .A(n_73), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_74), .Y(n_191) );
INVx1_ASAP7_75t_L g265 ( .A(n_75), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_76), .A2(n_104), .B1(n_113), .B2(n_763), .Y(n_103) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_78), .A2(n_155), .B(n_159), .C(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_79), .B(n_515), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_80), .Y(n_758) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_81), .B(n_181), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_82), .B(n_214), .Y(n_227) );
INVx2_ASAP7_75t_L g145 ( .A(n_83), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_84), .B(n_164), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_85), .B(n_181), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_86), .A2(n_155), .B(n_159), .C(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g109 ( .A(n_87), .Y(n_109) );
OR2x2_ASAP7_75t_L g120 ( .A(n_87), .B(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g462 ( .A(n_87), .B(n_122), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_89), .A2(n_102), .B1(n_181), .B2(n_182), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_90), .B(n_202), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g218 ( .A(n_91), .Y(n_218) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_92), .A2(n_155), .B(n_159), .C(n_241), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g248 ( .A(n_93), .Y(n_248) );
INVx1_ASAP7_75t_L g162 ( .A(n_94), .Y(n_162) );
CKINVDCx16_ASAP7_75t_R g254 ( .A(n_95), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_96), .B(n_214), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_97), .B(n_181), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_98), .B(n_143), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_99), .B(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_100), .A2(n_150), .B(n_157), .Y(n_149) );
OAI22xp5_ASAP7_75t_SL g755 ( .A1(n_101), .A2(n_756), .B1(n_757), .B2(n_760), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_101), .Y(n_760) );
INVx1_ASAP7_75t_L g763 ( .A(n_104), .Y(n_763) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
OR2x2_ASAP7_75t_L g463 ( .A(n_109), .B(n_122), .Y(n_463) );
NOR2x2_ASAP7_75t_L g749 ( .A(n_109), .B(n_121), .Y(n_749) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AOI22x1_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_126), .B1(n_750), .B2(n_752), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_118), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g751 ( .A(n_116), .Y(n_751) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g752 ( .A1(n_118), .A2(n_753), .B(n_761), .Y(n_752) );
NOR2xp33_ASAP7_75t_SL g118 ( .A(n_119), .B(n_125), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g762 ( .A(n_120), .Y(n_762) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_124), .Y(n_122) );
CKINVDCx14_ASAP7_75t_R g741 ( .A(n_127), .Y(n_741) );
INVx1_ASAP7_75t_L g131 ( .A(n_128), .Y(n_131) );
OAI22x1_ASAP7_75t_SL g133 ( .A1(n_134), .A2(n_460), .B1(n_463), .B2(n_464), .Y(n_133) );
OAI22xp5_ASAP7_75t_L g753 ( .A1(n_134), .A2(n_135), .B1(n_754), .B2(n_755), .Y(n_753) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_135), .A2(n_743), .B1(n_744), .B2(n_746), .Y(n_742) );
AND2x2_ASAP7_75t_SL g135 ( .A(n_136), .B(n_397), .Y(n_135) );
NOR4xp25_ASAP7_75t_L g136 ( .A(n_137), .B(n_327), .C(n_358), .D(n_377), .Y(n_136) );
NAND4xp25_ASAP7_75t_L g137 ( .A(n_138), .B(n_285), .C(n_300), .D(n_318), .Y(n_137) );
AOI222xp33_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_220), .B1(n_261), .B2(n_273), .C1(n_278), .C2(n_280), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_203), .Y(n_139) );
INVx1_ASAP7_75t_L g341 ( .A(n_140), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_174), .Y(n_140) );
AND2x2_ASAP7_75t_L g204 ( .A(n_141), .B(n_192), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_141), .B(n_207), .Y(n_370) );
INVx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
OR2x2_ASAP7_75t_L g277 ( .A(n_142), .B(n_176), .Y(n_277) );
AND2x2_ASAP7_75t_L g286 ( .A(n_142), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g312 ( .A(n_142), .Y(n_312) );
AND2x2_ASAP7_75t_L g333 ( .A(n_142), .B(n_176), .Y(n_333) );
BUFx2_ASAP7_75t_L g356 ( .A(n_142), .Y(n_356) );
AND2x2_ASAP7_75t_L g380 ( .A(n_142), .B(n_177), .Y(n_380) );
AND2x2_ASAP7_75t_L g444 ( .A(n_142), .B(n_192), .Y(n_444) );
OA21x2_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_149), .B(n_171), .Y(n_142) );
INVx4_ASAP7_75t_L g173 ( .A(n_143), .Y(n_173) );
OA21x2_ASAP7_75t_L g481 ( .A1(n_143), .A2(n_482), .B(n_490), .Y(n_481) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g178 ( .A(n_144), .Y(n_178) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
AND2x2_ASAP7_75t_SL g202 ( .A(n_145), .B(n_146), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
BUFx2_ASAP7_75t_L g252 ( .A(n_150), .Y(n_252) );
AND2x4_ASAP7_75t_L g150 ( .A(n_151), .B(n_155), .Y(n_150) );
NAND2x1p5_ASAP7_75t_L g189 ( .A(n_151), .B(n_155), .Y(n_189) );
AND2x2_ASAP7_75t_L g151 ( .A(n_152), .B(n_154), .Y(n_151) );
INVx1_ASAP7_75t_L g489 ( .A(n_152), .Y(n_489) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g160 ( .A(n_153), .Y(n_160) );
INVx1_ASAP7_75t_L g182 ( .A(n_153), .Y(n_182) );
INVx1_ASAP7_75t_L g161 ( .A(n_154), .Y(n_161) );
INVx1_ASAP7_75t_L g164 ( .A(n_154), .Y(n_164) );
INVx3_ASAP7_75t_L g167 ( .A(n_154), .Y(n_167) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_154), .Y(n_184) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_154), .Y(n_198) );
INVx4_ASAP7_75t_SL g170 ( .A(n_155), .Y(n_170) );
BUFx3_ASAP7_75t_L g477 ( .A(n_155), .Y(n_477) );
OAI21xp5_ASAP7_75t_L g482 ( .A1(n_155), .A2(n_483), .B(n_486), .Y(n_482) );
OAI21xp5_ASAP7_75t_L g492 ( .A1(n_155), .A2(n_493), .B(n_497), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_155), .A2(n_508), .B(n_512), .Y(n_507) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_155), .A2(n_532), .B(n_535), .Y(n_531) );
O2A1O1Ixp33_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_162), .B(n_163), .C(n_170), .Y(n_157) );
O2A1O1Ixp33_ASAP7_75t_L g194 ( .A1(n_158), .A2(n_170), .B(n_195), .C(n_196), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g253 ( .A1(n_158), .A2(n_170), .B(n_254), .C(n_255), .Y(n_253) );
INVx5_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x6_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_160), .Y(n_169) );
BUFx3_ASAP7_75t_L g231 ( .A(n_160), .Y(n_231) );
INVx1_ASAP7_75t_L g515 ( .A(n_160), .Y(n_515) );
INVx1_ASAP7_75t_L g511 ( .A(n_164), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_167), .B(n_200), .Y(n_199) );
INVx5_ASAP7_75t_L g214 ( .A(n_167), .Y(n_214) );
OAI22xp5_ASAP7_75t_SL g519 ( .A1(n_167), .A2(n_198), .B1(n_520), .B2(n_521), .Y(n_519) );
O2A1O1Ixp5_ASAP7_75t_SL g532 ( .A1(n_168), .A2(n_214), .B(n_533), .C(n_534), .Y(n_532) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_169), .Y(n_245) );
OAI22xp33_ASAP7_75t_L g179 ( .A1(n_170), .A2(n_180), .B1(n_188), .B2(n_189), .Y(n_179) );
OA21x2_ASAP7_75t_L g192 ( .A1(n_172), .A2(n_193), .B(n_201), .Y(n_192) );
INVx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_SL g233 ( .A(n_173), .B(n_234), .Y(n_233) );
NAND3xp33_ASAP7_75t_L g472 ( .A(n_173), .B(n_473), .C(n_477), .Y(n_472) );
AO21x1_ASAP7_75t_L g565 ( .A1(n_173), .A2(n_473), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g345 ( .A(n_174), .B(n_276), .Y(n_345) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_175), .B(n_370), .Y(n_369) );
OR2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_192), .Y(n_175) );
OR2x2_ASAP7_75t_L g305 ( .A(n_176), .B(n_208), .Y(n_305) );
AND2x2_ASAP7_75t_L g317 ( .A(n_176), .B(n_276), .Y(n_317) );
BUFx2_ASAP7_75t_L g449 ( .A(n_176), .Y(n_449) );
INVx3_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
OR2x2_ASAP7_75t_L g206 ( .A(n_177), .B(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g299 ( .A(n_177), .B(n_208), .Y(n_299) );
AND2x2_ASAP7_75t_L g352 ( .A(n_177), .B(n_192), .Y(n_352) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_177), .Y(n_388) );
AO21x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_190), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_178), .B(n_191), .Y(n_190) );
AO21x2_ASAP7_75t_L g208 ( .A1(n_178), .A2(n_209), .B(n_217), .Y(n_208) );
INVx2_ASAP7_75t_L g232 ( .A(n_178), .Y(n_232) );
INVx2_ASAP7_75t_L g216 ( .A(n_181), .Y(n_216) );
INVx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
OAI22xp5_ASAP7_75t_SL g183 ( .A1(n_184), .A2(n_185), .B1(n_186), .B2(n_187), .Y(n_183) );
INVx2_ASAP7_75t_L g186 ( .A(n_184), .Y(n_186) );
INVx4_ASAP7_75t_L g256 ( .A(n_184), .Y(n_256) );
OAI21xp5_ASAP7_75t_L g209 ( .A1(n_189), .A2(n_210), .B(n_211), .Y(n_209) );
OAI21xp5_ASAP7_75t_L g264 ( .A1(n_189), .A2(n_265), .B(n_266), .Y(n_264) );
AND2x2_ASAP7_75t_L g275 ( .A(n_192), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_SL g287 ( .A(n_192), .Y(n_287) );
INVx2_ASAP7_75t_L g298 ( .A(n_192), .Y(n_298) );
BUFx2_ASAP7_75t_L g322 ( .A(n_192), .Y(n_322) );
AND2x2_ASAP7_75t_SL g379 ( .A(n_192), .B(n_380), .Y(n_379) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_197), .A2(n_513), .B(n_514), .Y(n_512) );
O2A1O1Ixp5_ASAP7_75t_L g556 ( .A1(n_197), .A2(n_498), .B(n_557), .C(n_558), .Y(n_556) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx4_ASAP7_75t_L g244 ( .A(n_198), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_198), .A2(n_474), .B1(n_475), .B2(n_476), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_198), .A2(n_475), .B1(n_525), .B2(n_526), .Y(n_524) );
INVx1_ASAP7_75t_L g219 ( .A(n_202), .Y(n_219) );
INVx2_ASAP7_75t_L g238 ( .A(n_202), .Y(n_238) );
OA21x2_ASAP7_75t_L g250 ( .A1(n_202), .A2(n_251), .B(n_260), .Y(n_250) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_202), .A2(n_507), .B(n_516), .Y(n_506) );
OA21x2_ASAP7_75t_L g530 ( .A1(n_202), .A2(n_531), .B(n_538), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
AOI332xp33_ASAP7_75t_L g300 ( .A1(n_204), .A2(n_301), .A3(n_305), .B1(n_306), .B2(n_310), .B3(n_313), .C1(n_314), .C2(n_316), .Y(n_300) );
NAND2x1_ASAP7_75t_L g385 ( .A(n_204), .B(n_276), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_204), .B(n_290), .Y(n_436) );
A2O1A1Ixp33_ASAP7_75t_SL g318 ( .A1(n_205), .A2(n_319), .B(n_322), .C(n_323), .Y(n_318) );
AND2x2_ASAP7_75t_L g457 ( .A(n_205), .B(n_298), .Y(n_457) );
INVx3_ASAP7_75t_SL g205 ( .A(n_206), .Y(n_205) );
OR2x2_ASAP7_75t_L g354 ( .A(n_206), .B(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g359 ( .A(n_206), .B(n_356), .Y(n_359) );
INVx1_ASAP7_75t_L g290 ( .A(n_207), .Y(n_290) );
AND2x2_ASAP7_75t_L g393 ( .A(n_207), .B(n_352), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_207), .B(n_333), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_207), .B(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_207), .B(n_311), .Y(n_419) );
INVx3_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx3_ASAP7_75t_L g276 ( .A(n_208), .Y(n_276) );
O2A1O1Ixp33_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_215), .C(n_216), .Y(n_212) );
INVx2_ASAP7_75t_L g475 ( .A(n_214), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_214), .A2(n_484), .B(n_485), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_214), .A2(n_554), .B(n_555), .Y(n_553) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_216), .A2(n_494), .B(n_495), .C(n_496), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_218), .B(n_219), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_219), .B(n_248), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_219), .B(n_272), .Y(n_271) );
OAI31xp33_ASAP7_75t_L g458 ( .A1(n_220), .A2(n_379), .A3(n_386), .B(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_235), .Y(n_220) );
AND2x2_ASAP7_75t_L g261 ( .A(n_221), .B(n_262), .Y(n_261) );
NAND2x1_ASAP7_75t_SL g281 ( .A(n_221), .B(n_282), .Y(n_281) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_221), .Y(n_368) );
AND2x2_ASAP7_75t_L g373 ( .A(n_221), .B(n_284), .Y(n_373) );
INVx3_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
A2O1A1Ixp33_ASAP7_75t_L g285 ( .A1(n_222), .A2(n_286), .B(n_288), .C(n_291), .Y(n_285) );
OR2x2_ASAP7_75t_L g302 ( .A(n_222), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g315 ( .A(n_222), .Y(n_315) );
AND2x2_ASAP7_75t_L g321 ( .A(n_222), .B(n_263), .Y(n_321) );
INVx2_ASAP7_75t_L g339 ( .A(n_222), .Y(n_339) );
AND2x2_ASAP7_75t_L g350 ( .A(n_222), .B(n_304), .Y(n_350) );
AND2x2_ASAP7_75t_L g382 ( .A(n_222), .B(n_340), .Y(n_382) );
AND2x2_ASAP7_75t_L g386 ( .A(n_222), .B(n_309), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_222), .B(n_235), .Y(n_391) );
AND2x2_ASAP7_75t_L g425 ( .A(n_222), .B(n_426), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_222), .B(n_328), .Y(n_459) );
OR2x6_ASAP7_75t_L g222 ( .A(n_223), .B(n_233), .Y(n_222) );
AOI21xp5_ASAP7_75t_SL g223 ( .A1(n_224), .A2(n_225), .B(n_232), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_229), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_229), .A2(n_268), .B(n_269), .Y(n_267) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g259 ( .A(n_231), .Y(n_259) );
INVx1_ASAP7_75t_L g270 ( .A(n_232), .Y(n_270) );
OA21x2_ASAP7_75t_L g491 ( .A1(n_232), .A2(n_492), .B(n_501), .Y(n_491) );
OA21x2_ASAP7_75t_L g551 ( .A1(n_232), .A2(n_552), .B(n_559), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_235), .B(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g367 ( .A(n_235), .Y(n_367) );
AND2x2_ASAP7_75t_L g429 ( .A(n_235), .B(n_350), .Y(n_429) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_249), .Y(n_235) );
OR2x2_ASAP7_75t_L g283 ( .A(n_236), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g293 ( .A(n_236), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_236), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g401 ( .A(n_236), .Y(n_401) );
AND2x2_ASAP7_75t_L g418 ( .A(n_236), .B(n_263), .Y(n_418) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g309 ( .A(n_237), .B(n_249), .Y(n_309) );
AND2x2_ASAP7_75t_L g338 ( .A(n_237), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g349 ( .A(n_237), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_237), .B(n_304), .Y(n_440) );
AO21x2_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B(n_247), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_240), .B(n_246), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B(n_245), .Y(n_241) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g262 ( .A(n_250), .B(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g284 ( .A(n_250), .Y(n_284) );
AND2x2_ASAP7_75t_L g340 ( .A(n_250), .B(n_304), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_256), .B(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g496 ( .A(n_256), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_256), .A2(n_536), .B(n_537), .Y(n_535) );
INVx1_ASAP7_75t_L g442 ( .A(n_261), .Y(n_442) );
INVx1_ASAP7_75t_L g446 ( .A(n_262), .Y(n_446) );
INVx2_ASAP7_75t_L g304 ( .A(n_263), .Y(n_304) );
AO21x2_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_270), .B(n_271), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_274), .B(n_277), .Y(n_273) );
INVx1_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_275), .B(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_275), .B(n_380), .Y(n_438) );
OR2x2_ASAP7_75t_L g279 ( .A(n_276), .B(n_277), .Y(n_279) );
INVx1_ASAP7_75t_SL g331 ( .A(n_276), .Y(n_331) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AOI221xp5_ASAP7_75t_L g334 ( .A1(n_282), .A2(n_335), .B1(n_337), .B2(n_341), .C(n_342), .Y(n_334) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g362 ( .A(n_283), .B(n_326), .Y(n_362) );
INVx2_ASAP7_75t_L g294 ( .A(n_284), .Y(n_294) );
INVx1_ASAP7_75t_L g320 ( .A(n_284), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_284), .B(n_304), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_284), .B(n_307), .Y(n_414) );
INVx1_ASAP7_75t_L g422 ( .A(n_284), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_286), .B(n_290), .Y(n_336) );
AND2x4_ASAP7_75t_L g311 ( .A(n_287), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g424 ( .A(n_290), .B(n_380), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_292), .B(n_295), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_293), .B(n_325), .Y(n_324) );
INVxp67_ASAP7_75t_L g432 ( .A(n_294), .Y(n_432) );
INVxp67_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g332 ( .A(n_298), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g404 ( .A(n_298), .B(n_380), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_298), .B(n_317), .Y(n_410) );
AOI322xp5_ASAP7_75t_L g364 ( .A1(n_299), .A2(n_333), .A3(n_340), .B1(n_365), .B2(n_368), .C1(n_369), .C2(n_371), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_299), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g430 ( .A(n_302), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g376 ( .A(n_303), .Y(n_376) );
INVx2_ASAP7_75t_L g307 ( .A(n_304), .Y(n_307) );
INVx1_ASAP7_75t_L g366 ( .A(n_304), .Y(n_366) );
CKINVDCx16_ASAP7_75t_R g313 ( .A(n_305), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
AND2x2_ASAP7_75t_L g402 ( .A(n_307), .B(n_315), .Y(n_402) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g314 ( .A(n_309), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g357 ( .A(n_309), .B(n_350), .Y(n_357) );
AND2x2_ASAP7_75t_L g361 ( .A(n_309), .B(n_321), .Y(n_361) );
OAI21xp33_ASAP7_75t_SL g371 ( .A1(n_310), .A2(n_372), .B(n_374), .Y(n_371) );
OAI22xp33_ASAP7_75t_L g441 ( .A1(n_310), .A2(n_442), .B1(n_443), .B2(n_445), .Y(n_441) );
INVx3_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g316 ( .A(n_311), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_311), .B(n_331), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_313), .B(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx1_ASAP7_75t_L g453 ( .A(n_320), .Y(n_453) );
INVx4_ASAP7_75t_L g326 ( .A(n_321), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_321), .B(n_348), .Y(n_396) );
INVx1_ASAP7_75t_SL g408 ( .A(n_322), .Y(n_408) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NOR2xp67_ASAP7_75t_L g421 ( .A(n_326), .B(n_422), .Y(n_421) );
OAI211xp5_ASAP7_75t_SL g327 ( .A1(n_328), .A2(n_329), .B(n_334), .C(n_351), .Y(n_327) );
OAI221xp5_ASAP7_75t_SL g447 ( .A1(n_329), .A2(n_367), .B1(n_446), .B2(n_448), .C(n_450), .Y(n_447) );
INVx1_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_331), .B(n_444), .Y(n_443) );
OAI31xp33_ASAP7_75t_L g423 ( .A1(n_332), .A2(n_409), .A3(n_424), .B(n_425), .Y(n_423) );
INVx1_ASAP7_75t_L g363 ( .A(n_333), .Y(n_363) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_340), .Y(n_337) );
INVx1_ASAP7_75t_L g413 ( .A(n_338), .Y(n_413) );
AND2x2_ASAP7_75t_L g426 ( .A(n_340), .B(n_349), .Y(n_426) );
AOI21xp33_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_344), .B(n_346), .Y(n_342) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
INVxp67_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_350), .B(n_453), .Y(n_452) );
OAI21xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_353), .B(n_357), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OAI221xp5_ASAP7_75t_SL g358 ( .A1(n_359), .A2(n_360), .B1(n_362), .B2(n_363), .C(n_364), .Y(n_358) );
A2O1A1Ixp33_ASAP7_75t_L g427 ( .A1(n_359), .A2(n_428), .B(n_430), .C(n_433), .Y(n_427) );
CKINVDCx16_ASAP7_75t_R g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_362), .B(n_412), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx1_ASAP7_75t_L g389 ( .A(n_370), .Y(n_389) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g375 ( .A(n_373), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g417 ( .A(n_373), .B(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI211xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_381), .B(n_383), .C(n_392), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OAI221xp5_ASAP7_75t_L g454 ( .A1(n_381), .A2(n_391), .B1(n_455), .B2(n_456), .C(n_458), .Y(n_454) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_386), .B1(n_387), .B2(n_390), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OAI21xp5_ASAP7_75t_SL g392 ( .A1(n_393), .A2(n_394), .B(n_395), .Y(n_392) );
INVx1_ASAP7_75t_SL g455 ( .A(n_394), .Y(n_455) );
INVxp67_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NOR4xp25_ASAP7_75t_L g397 ( .A(n_398), .B(n_427), .C(n_447), .D(n_454), .Y(n_397) );
OAI211xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_403), .B(n_405), .C(n_423), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_402), .Y(n_399) );
INVxp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
O2A1O1Ixp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_409), .B(n_411), .C(n_415), .Y(n_405) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g434 ( .A(n_412), .Y(n_434) );
OR2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
OR2x2_ASAP7_75t_L g445 ( .A(n_413), .B(n_446), .Y(n_445) );
OAI21xp33_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_419), .B(n_420), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AOI221xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B1(n_437), .B2(n_439), .C(n_441), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVxp67_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_444), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g743 ( .A(n_461), .Y(n_743) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g745 ( .A(n_463), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_464), .Y(n_746) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_SL g465 ( .A(n_466), .B(n_675), .Y(n_465) );
NOR5xp2_ASAP7_75t_L g466 ( .A(n_467), .B(n_588), .C(n_634), .D(n_647), .E(n_659), .Y(n_466) );
OAI211xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_502), .B(n_542), .C(n_569), .Y(n_467) );
INVx1_ASAP7_75t_SL g670 ( .A(n_468), .Y(n_670) );
OR2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_478), .Y(n_468) );
AND2x2_ASAP7_75t_L g594 ( .A(n_469), .B(n_479), .Y(n_594) );
AND2x2_ASAP7_75t_L g622 ( .A(n_469), .B(n_568), .Y(n_622) );
AND2x2_ASAP7_75t_L g630 ( .A(n_469), .B(n_573), .Y(n_630) );
INVx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g560 ( .A(n_470), .B(n_480), .Y(n_560) );
INVx2_ASAP7_75t_L g572 ( .A(n_470), .Y(n_572) );
AND2x2_ASAP7_75t_L g697 ( .A(n_470), .B(n_639), .Y(n_697) );
OR2x2_ASAP7_75t_L g699 ( .A(n_470), .B(n_700), .Y(n_699) );
AND2x4_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
INVx1_ASAP7_75t_L g566 ( .A(n_471), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_475), .A2(n_487), .B(n_488), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_L g497 ( .A1(n_475), .A2(n_498), .B(n_499), .C(n_500), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g552 ( .A1(n_477), .A2(n_553), .B(n_556), .Y(n_552) );
INVx2_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g610 ( .A(n_479), .B(n_582), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_479), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g724 ( .A(n_479), .B(n_564), .Y(n_724) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_491), .Y(n_479) );
AND2x2_ASAP7_75t_L g567 ( .A(n_480), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g614 ( .A(n_480), .Y(n_614) );
AND2x2_ASAP7_75t_L g639 ( .A(n_480), .B(n_551), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_480), .B(n_672), .Y(n_709) );
INVx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g573 ( .A(n_481), .B(n_551), .Y(n_573) );
AND2x2_ASAP7_75t_L g587 ( .A(n_481), .B(n_550), .Y(n_587) );
AND2x2_ASAP7_75t_L g604 ( .A(n_481), .B(n_491), .Y(n_604) );
AND2x2_ASAP7_75t_L g661 ( .A(n_481), .B(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_481), .B(n_568), .Y(n_674) );
AND2x2_ASAP7_75t_L g726 ( .A(n_481), .B(n_651), .Y(n_726) );
INVx2_ASAP7_75t_L g498 ( .A(n_489), .Y(n_498) );
AND2x2_ASAP7_75t_L g549 ( .A(n_491), .B(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g568 ( .A(n_491), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_491), .B(n_551), .Y(n_645) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_527), .B(n_539), .Y(n_502) );
INVx1_ASAP7_75t_SL g658 ( .A(n_503), .Y(n_658) );
AND2x4_ASAP7_75t_L g503 ( .A(n_504), .B(n_517), .Y(n_503) );
BUFx3_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_SL g546 ( .A(n_505), .B(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g541 ( .A(n_506), .Y(n_541) );
INVx1_ASAP7_75t_L g578 ( .A(n_506), .Y(n_578) );
AND2x2_ASAP7_75t_L g599 ( .A(n_506), .B(n_522), .Y(n_599) );
AND2x2_ASAP7_75t_L g633 ( .A(n_506), .B(n_523), .Y(n_633) );
OR2x2_ASAP7_75t_L g652 ( .A(n_506), .B(n_529), .Y(n_652) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_506), .Y(n_666) );
AND2x2_ASAP7_75t_L g679 ( .A(n_506), .B(n_680), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_510), .B(n_511), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_517), .A2(n_601), .B1(n_602), .B2(n_611), .Y(n_600) );
AND2x2_ASAP7_75t_L g684 ( .A(n_517), .B(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_522), .Y(n_517) );
INVx1_ASAP7_75t_L g545 ( .A(n_518), .Y(n_545) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_518), .Y(n_582) );
INVx1_ASAP7_75t_L g593 ( .A(n_518), .Y(n_593) );
AND2x2_ASAP7_75t_L g608 ( .A(n_518), .B(n_523), .Y(n_608) );
OR2x2_ASAP7_75t_L g562 ( .A(n_522), .B(n_547), .Y(n_562) );
AND2x2_ASAP7_75t_L g592 ( .A(n_522), .B(n_593), .Y(n_592) );
NOR2xp67_ASAP7_75t_L g680 ( .A(n_522), .B(n_681), .Y(n_680) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g540 ( .A(n_523), .B(n_541), .Y(n_540) );
BUFx2_ASAP7_75t_L g649 ( .A(n_523), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_527), .B(n_665), .Y(n_664) );
BUFx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g627 ( .A(n_528), .B(n_593), .Y(n_627) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g539 ( .A(n_529), .B(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g598 ( .A(n_529), .Y(n_598) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g547 ( .A(n_530), .Y(n_547) );
OR2x2_ASAP7_75t_L g577 ( .A(n_530), .B(n_578), .Y(n_577) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_530), .Y(n_632) );
AOI32xp33_ASAP7_75t_L g669 ( .A1(n_539), .A2(n_599), .A3(n_670), .B1(n_671), .B2(n_673), .Y(n_669) );
AND2x2_ASAP7_75t_L g595 ( .A(n_540), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_540), .B(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_540), .B(n_627), .Y(n_713) );
INVx1_ASAP7_75t_L g718 ( .A(n_540), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_548), .B1(n_561), .B2(n_563), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_546), .Y(n_543) );
AND2x2_ASAP7_75t_L g648 ( .A(n_544), .B(n_649), .Y(n_648) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_545), .B(n_547), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_546), .A2(n_570), .B1(n_574), .B2(n_584), .Y(n_569) );
AND2x2_ASAP7_75t_L g591 ( .A(n_546), .B(n_592), .Y(n_591) );
A2O1A1Ixp33_ASAP7_75t_L g642 ( .A1(n_546), .A2(n_560), .B(n_608), .C(n_643), .Y(n_642) );
OAI332xp33_ASAP7_75t_L g647 ( .A1(n_546), .A2(n_648), .A3(n_650), .B1(n_652), .B2(n_653), .B3(n_655), .C1(n_656), .C2(n_658), .Y(n_647) );
INVx2_ASAP7_75t_L g688 ( .A(n_546), .Y(n_688) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_547), .Y(n_606) );
INVx1_ASAP7_75t_L g681 ( .A(n_547), .Y(n_681) );
AND2x2_ASAP7_75t_L g735 ( .A(n_547), .B(n_599), .Y(n_735) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_560), .Y(n_548) );
AND2x2_ASAP7_75t_L g615 ( .A(n_550), .B(n_565), .Y(n_615) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g564 ( .A(n_551), .B(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g663 ( .A(n_551), .B(n_565), .Y(n_663) );
INVx1_ASAP7_75t_L g672 ( .A(n_551), .Y(n_672) );
INVx1_ASAP7_75t_L g646 ( .A(n_560), .Y(n_646) );
INVxp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g730 ( .A(n_562), .B(n_582), .Y(n_730) );
INVx1_ASAP7_75t_SL g641 ( .A(n_563), .Y(n_641) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_567), .Y(n_563) );
AND2x2_ASAP7_75t_L g668 ( .A(n_564), .B(n_626), .Y(n_668) );
INVx1_ASAP7_75t_L g687 ( .A(n_564), .Y(n_687) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_564), .B(n_654), .Y(n_689) );
INVx1_ASAP7_75t_L g586 ( .A(n_565), .Y(n_586) );
AND2x2_ASAP7_75t_L g590 ( .A(n_567), .B(n_571), .Y(n_590) );
AND2x2_ASAP7_75t_L g657 ( .A(n_567), .B(n_615), .Y(n_657) );
INVx2_ASAP7_75t_L g700 ( .A(n_567), .Y(n_700) );
INVx2_ASAP7_75t_L g583 ( .A(n_568), .Y(n_583) );
AND2x2_ASAP7_75t_L g585 ( .A(n_568), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
INVx1_ASAP7_75t_L g601 ( .A(n_571), .Y(n_601) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_572), .B(n_645), .Y(n_651) );
OR2x2_ASAP7_75t_L g715 ( .A(n_572), .B(n_674), .Y(n_715) );
INVx1_ASAP7_75t_L g739 ( .A(n_572), .Y(n_739) );
INVx1_ASAP7_75t_L g695 ( .A(n_573), .Y(n_695) );
AND2x2_ASAP7_75t_L g740 ( .A(n_573), .B(n_583), .Y(n_740) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_579), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_577), .A2(n_603), .B1(n_605), .B2(n_609), .Y(n_602) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OAI322xp33_ASAP7_75t_SL g686 ( .A1(n_580), .A2(n_687), .A3(n_688), .B1(n_689), .B2(n_690), .C1(n_693), .C2(n_695), .Y(n_686) );
OR2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
AND2x2_ASAP7_75t_L g683 ( .A(n_581), .B(n_599), .Y(n_683) );
OR2x2_ASAP7_75t_L g717 ( .A(n_581), .B(n_718), .Y(n_717) );
OR2x2_ASAP7_75t_L g720 ( .A(n_581), .B(n_652), .Y(n_720) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g665 ( .A(n_582), .B(n_666), .Y(n_665) );
OR2x2_ASAP7_75t_L g721 ( .A(n_582), .B(n_652), .Y(n_721) );
INVx3_ASAP7_75t_L g654 ( .A(n_583), .Y(n_654) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_587), .Y(n_584) );
INVx1_ASAP7_75t_L g710 ( .A(n_585), .Y(n_710) );
AOI222xp33_ASAP7_75t_L g589 ( .A1(n_587), .A2(n_590), .B1(n_591), .B2(n_594), .C1(n_595), .C2(n_597), .Y(n_589) );
INVx1_ASAP7_75t_L g620 ( .A(n_587), .Y(n_620) );
NAND3xp33_ASAP7_75t_SL g588 ( .A(n_589), .B(n_600), .C(n_617), .Y(n_588) );
AND2x2_ASAP7_75t_L g705 ( .A(n_592), .B(n_606), .Y(n_705) );
BUFx2_ASAP7_75t_L g596 ( .A(n_593), .Y(n_596) );
INVx1_ASAP7_75t_L g637 ( .A(n_593), .Y(n_637) );
AOI221xp5_ASAP7_75t_L g682 ( .A1(n_594), .A2(n_630), .B1(n_683), .B2(n_684), .C(n_686), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_596), .B(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_599), .Y(n_623) );
AND2x2_ASAP7_75t_L g636 ( .A(n_599), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_604), .B(n_615), .Y(n_616) );
OR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
OAI21xp33_ASAP7_75t_L g611 ( .A1(n_606), .A2(n_612), .B(n_616), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_606), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g703 ( .A(n_608), .B(n_685), .Y(n_703) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
INVx1_ASAP7_75t_L g626 ( .A(n_614), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_615), .B(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g732 ( .A(n_615), .Y(n_732) );
AOI221xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_623), .B1(n_624), .B2(n_627), .C(n_628), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g707 ( .A(n_619), .B(n_708), .Y(n_707) );
OR2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g728 ( .A(n_627), .B(n_633), .Y(n_728) );
INVxp67_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
OAI31xp33_ASAP7_75t_SL g696 ( .A1(n_631), .A2(n_670), .A3(n_697), .B(n_698), .Y(n_696) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx1_ASAP7_75t_L g685 ( .A(n_632), .Y(n_685) );
NAND2xp5_ASAP7_75t_SL g736 ( .A(n_633), .B(n_637), .Y(n_736) );
OAI221xp5_ASAP7_75t_SL g634 ( .A1(n_635), .A2(n_638), .B1(n_640), .B2(n_641), .C(n_642), .Y(n_634) );
INVx1_ASAP7_75t_L g640 ( .A(n_636), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_639), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
INVx1_ASAP7_75t_L g655 ( .A(n_648), .Y(n_655) );
INVx2_ASAP7_75t_L g691 ( .A(n_649), .Y(n_691) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OR2x2_ASAP7_75t_L g677 ( .A(n_654), .B(n_663), .Y(n_677) );
A2O1A1Ixp33_ASAP7_75t_L g727 ( .A1(n_654), .A2(n_671), .B(n_728), .C(n_729), .Y(n_727) );
OAI221xp5_ASAP7_75t_SL g659 ( .A1(n_655), .A2(n_660), .B1(n_664), .B2(n_667), .C(n_669), .Y(n_659) );
INVx1_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
A2O1A1Ixp33_ASAP7_75t_L g722 ( .A1(n_658), .A2(n_723), .B(n_725), .C(n_727), .Y(n_722) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AOI221xp5_ASAP7_75t_L g711 ( .A1(n_661), .A2(n_712), .B1(n_714), .B2(n_716), .C(n_719), .Y(n_711) );
INVx1_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
NOR4xp25_ASAP7_75t_L g675 ( .A(n_676), .B(n_701), .C(n_722), .D(n_733), .Y(n_675) );
OAI211xp5_ASAP7_75t_SL g676 ( .A1(n_677), .A2(n_678), .B(n_682), .C(n_696), .Y(n_676) );
INVx1_ASAP7_75t_SL g731 ( .A(n_683), .Y(n_731) );
OR2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
INVx1_ASAP7_75t_SL g694 ( .A(n_692), .Y(n_694) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_699), .A2(n_708), .B1(n_720), .B2(n_721), .Y(n_719) );
A2O1A1Ixp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_704), .B(n_706), .C(n_711), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AOI31xp33_ASAP7_75t_L g733 ( .A1(n_704), .A2(n_734), .A3(n_736), .B(n_737), .Y(n_733) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVxp67_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OR2x2_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_731), .B(n_732), .Y(n_729) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_740), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_755), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
endmodule