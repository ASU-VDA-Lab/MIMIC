module fake_netlist_6_1052_n_123 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_6, n_15, n_3, n_14, n_0, n_4, n_22, n_13, n_11, n_17, n_12, n_20, n_7, n_2, n_5, n_19, n_123);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_13;
input n_11;
input n_17;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;

output n_123;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_121;
wire n_23;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_109;
wire n_122;
wire n_45;
wire n_34;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_110;
wire n_61;
wire n_112;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_94;
wire n_97;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_60;
wire n_35;
wire n_115;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_19),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVxp67_ASAP7_75t_SL g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVxp67_ASAP7_75t_SL g36 ( 
.A(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_23),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_36),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_25),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_28),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_44),
.Y(n_63)
);

BUFx4_ASAP7_75t_SL g64 ( 
.A(n_54),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_46),
.Y(n_65)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_60),
.B(n_32),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_51),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

AOI21x1_ASAP7_75t_SL g71 ( 
.A1(n_67),
.A2(n_59),
.B(n_53),
.Y(n_71)
);

CKINVDCx12_ASAP7_75t_R g72 ( 
.A(n_65),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

AND2x4_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_30),
.Y(n_74)
);

AND2x4_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_65),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_74),
.A2(n_63),
.B(n_66),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_78),
.A2(n_73),
.B(n_75),
.C(n_74),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_75),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_83),
.A2(n_77),
.B1(n_73),
.B2(n_75),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_84),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_75),
.Y(n_90)
);

AND2x4_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_80),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_73),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_57),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_73),
.B1(n_35),
.B2(n_90),
.Y(n_95)
);

AND2x4_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_89),
.Y(n_96)
);

INVxp67_ASAP7_75t_SL g97 ( 
.A(n_94),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_89),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_92),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_92),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_45),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_87),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_41),
.Y(n_104)
);

NAND3x1_ASAP7_75t_SL g105 ( 
.A(n_102),
.B(n_64),
.C(n_95),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_103),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_43),
.Y(n_108)
);

NAND3x1_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_41),
.C(n_4),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

AOI22x1_ASAP7_75t_L g111 ( 
.A1(n_105),
.A2(n_62),
.B1(n_55),
.B2(n_58),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_52),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_5),
.Y(n_113)
);

OR5x1_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_7),
.C(n_71),
.D(n_13),
.E(n_14),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_112),
.A2(n_7),
.B1(n_52),
.B2(n_58),
.Y(n_115)
);

XNOR2x1_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_10),
.Y(n_116)
);

AND3x4_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_74),
.C(n_71),
.Y(n_117)
);

NAND4xp75_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_15),
.C(n_16),
.D(n_17),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_114),
.A2(n_74),
.B1(n_22),
.B2(n_20),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_116),
.B1(n_76),
.B2(n_56),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_118),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_122),
.A2(n_120),
.B1(n_117),
.B2(n_76),
.Y(n_123)
);


endmodule