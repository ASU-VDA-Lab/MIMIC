module real_aes_8473_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_755;
wire n_153;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_449;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_502;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g238 ( .A1(n_0), .A2(n_239), .B(n_240), .C(n_244), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_1), .B(n_180), .Y(n_245) );
INVx1_ASAP7_75t_L g110 ( .A(n_2), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_3), .B(n_152), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_4), .A2(n_138), .B(n_143), .C(n_505), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_5), .A2(n_133), .B(n_543), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_6), .A2(n_133), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_7), .B(n_180), .Y(n_549) );
AO21x2_ASAP7_75t_L g183 ( .A1(n_8), .A2(n_168), .B(n_184), .Y(n_183) );
AND2x6_ASAP7_75t_L g138 ( .A(n_9), .B(n_139), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_10), .A2(n_138), .B(n_143), .C(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g487 ( .A(n_11), .Y(n_487) );
INVx1_ASAP7_75t_L g107 ( .A(n_12), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_12), .B(n_42), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_13), .B(n_243), .Y(n_507) );
INVx1_ASAP7_75t_L g162 ( .A(n_14), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_15), .B(n_152), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_16), .A2(n_153), .B(n_495), .C(n_497), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_17), .B(n_180), .Y(n_498) );
AOI222xp33_ASAP7_75t_L g468 ( .A1(n_18), .A2(n_469), .B1(n_746), .B2(n_752), .C1(n_755), .C2(n_756), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_19), .B(n_217), .Y(n_586) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_20), .A2(n_143), .B(n_194), .C(n_213), .Y(n_212) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_21), .A2(n_192), .B(n_242), .C(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_22), .B(n_243), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_23), .B(n_243), .Y(n_527) );
CKINVDCx16_ASAP7_75t_R g534 ( .A(n_24), .Y(n_534) );
INVx1_ASAP7_75t_L g526 ( .A(n_25), .Y(n_526) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_26), .A2(n_143), .B(n_187), .C(n_194), .Y(n_186) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_27), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_28), .Y(n_503) );
INVx1_ASAP7_75t_L g583 ( .A(n_29), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_30), .A2(n_133), .B(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g136 ( .A(n_31), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_32), .A2(n_141), .B(n_156), .C(n_202), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_33), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_34), .A2(n_242), .B(n_546), .C(n_548), .Y(n_545) );
INVxp67_ASAP7_75t_L g584 ( .A(n_35), .Y(n_584) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_36), .A2(n_47), .B1(n_124), .B2(n_125), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_36), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_37), .B(n_189), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_38), .A2(n_143), .B(n_194), .C(n_525), .Y(n_524) );
CKINVDCx14_ASAP7_75t_R g544 ( .A(n_39), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_40), .A2(n_46), .B1(n_750), .B2(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_40), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_41), .A2(n_104), .B1(n_115), .B2(n_762), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_42), .B(n_107), .Y(n_106) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_43), .A2(n_244), .B(n_485), .C(n_486), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_44), .B(n_211), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g258 ( .A(n_45), .Y(n_258) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_46), .Y(n_750) );
INVx1_ASAP7_75t_L g125 ( .A(n_47), .Y(n_125) );
OAI321xp33_ASAP7_75t_L g121 ( .A1(n_48), .A2(n_122), .A3(n_456), .B1(n_462), .B2(n_463), .C(n_465), .Y(n_121) );
INVx1_ASAP7_75t_L g462 ( .A(n_48), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_49), .B(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_50), .B(n_133), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_51), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g580 ( .A(n_52), .Y(n_580) );
A2O1A1Ixp33_ASAP7_75t_L g140 ( .A1(n_53), .A2(n_141), .B(n_146), .C(n_156), .Y(n_140) );
INVx1_ASAP7_75t_L g241 ( .A(n_54), .Y(n_241) );
INVx1_ASAP7_75t_L g147 ( .A(n_55), .Y(n_147) );
INVx1_ASAP7_75t_L g515 ( .A(n_56), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_57), .B(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_58), .B(n_133), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_59), .Y(n_220) );
CKINVDCx14_ASAP7_75t_R g483 ( .A(n_60), .Y(n_483) );
INVx1_ASAP7_75t_L g139 ( .A(n_61), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_62), .B(n_133), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_63), .B(n_180), .Y(n_179) );
A2O1A1Ixp33_ASAP7_75t_L g173 ( .A1(n_64), .A2(n_174), .B(n_176), .C(n_178), .Y(n_173) );
INVx1_ASAP7_75t_L g161 ( .A(n_65), .Y(n_161) );
INVx1_ASAP7_75t_SL g547 ( .A(n_66), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_67), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_68), .B(n_152), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_69), .B(n_180), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_70), .B(n_153), .Y(n_255) );
INVx1_ASAP7_75t_L g537 ( .A(n_71), .Y(n_537) );
CKINVDCx16_ASAP7_75t_R g237 ( .A(n_72), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_73), .B(n_149), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_74), .A2(n_143), .B(n_156), .C(n_226), .Y(n_225) );
CKINVDCx16_ASAP7_75t_R g172 ( .A(n_75), .Y(n_172) );
INVx1_ASAP7_75t_L g114 ( .A(n_76), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_77), .A2(n_133), .B(n_482), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_78), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_79), .A2(n_133), .B(n_492), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_80), .A2(n_211), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g493 ( .A(n_81), .Y(n_493) );
CKINVDCx16_ASAP7_75t_R g523 ( .A(n_82), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_83), .B(n_148), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_84), .A2(n_747), .B1(n_748), .B2(n_749), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_84), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g206 ( .A(n_85), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_86), .A2(n_133), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g496 ( .A(n_87), .Y(n_496) );
INVx2_ASAP7_75t_L g159 ( .A(n_88), .Y(n_159) );
INVx1_ASAP7_75t_L g506 ( .A(n_89), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_90), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_91), .B(n_243), .Y(n_256) );
INVx2_ASAP7_75t_L g111 ( .A(n_92), .Y(n_111) );
OR2x2_ASAP7_75t_L g458 ( .A(n_92), .B(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g745 ( .A(n_92), .B(n_460), .Y(n_745) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_93), .A2(n_143), .B(n_156), .C(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_94), .B(n_133), .Y(n_200) );
INVx1_ASAP7_75t_L g203 ( .A(n_95), .Y(n_203) );
INVxp67_ASAP7_75t_L g177 ( .A(n_96), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_97), .B(n_168), .Y(n_488) );
INVx2_ASAP7_75t_L g518 ( .A(n_98), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_99), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g227 ( .A(n_100), .Y(n_227) );
INVx1_ASAP7_75t_L g251 ( .A(n_101), .Y(n_251) );
AND2x2_ASAP7_75t_L g163 ( .A(n_102), .B(n_158), .Y(n_163) );
INVx2_ASAP7_75t_L g762 ( .A(n_104), .Y(n_762) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_108), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx14_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_110), .B(n_111), .C(n_112), .Y(n_109) );
AND2x2_ASAP7_75t_L g460 ( .A(n_110), .B(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g474 ( .A(n_111), .B(n_460), .Y(n_474) );
NOR2x2_ASAP7_75t_L g754 ( .A(n_111), .B(n_459), .Y(n_754) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_467), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx3_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g761 ( .A(n_119), .Y(n_761) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_122), .B(n_464), .Y(n_463) );
XOR2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_126), .Y(n_122) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_126), .A2(n_471), .B1(n_475), .B2(n_742), .Y(n_470) );
INVx4_ASAP7_75t_L g759 ( .A(n_126), .Y(n_759) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OR5x1_ASAP7_75t_L g127 ( .A(n_128), .B(n_329), .C(n_407), .D(n_431), .E(n_448), .Y(n_127) );
OAI211xp5_ASAP7_75t_SL g128 ( .A1(n_129), .A2(n_195), .B(n_246), .C(n_306), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_164), .Y(n_129) );
AND2x2_ASAP7_75t_L g260 ( .A(n_130), .B(n_166), .Y(n_260) );
INVx5_ASAP7_75t_SL g288 ( .A(n_130), .Y(n_288) );
AND2x2_ASAP7_75t_L g324 ( .A(n_130), .B(n_309), .Y(n_324) );
OR2x2_ASAP7_75t_L g363 ( .A(n_130), .B(n_165), .Y(n_363) );
OR2x2_ASAP7_75t_L g394 ( .A(n_130), .B(n_285), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_130), .B(n_298), .Y(n_430) );
AND2x2_ASAP7_75t_L g442 ( .A(n_130), .B(n_285), .Y(n_442) );
OR2x6_ASAP7_75t_L g130 ( .A(n_131), .B(n_163), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_140), .B(n_158), .Y(n_131) );
BUFx2_ASAP7_75t_L g211 ( .A(n_133), .Y(n_211) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_138), .Y(n_133) );
NAND2x1p5_ASAP7_75t_L g252 ( .A(n_134), .B(n_138), .Y(n_252) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
INVx1_ASAP7_75t_L g178 ( .A(n_135), .Y(n_178) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g144 ( .A(n_136), .Y(n_144) );
INVx1_ASAP7_75t_L g193 ( .A(n_136), .Y(n_193) );
INVx1_ASAP7_75t_L g145 ( .A(n_137), .Y(n_145) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_137), .Y(n_150) );
INVx3_ASAP7_75t_L g153 ( .A(n_137), .Y(n_153) );
INVx1_ASAP7_75t_L g189 ( .A(n_137), .Y(n_189) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_137), .Y(n_243) );
INVx4_ASAP7_75t_SL g157 ( .A(n_138), .Y(n_157) );
BUFx3_ASAP7_75t_L g194 ( .A(n_138), .Y(n_194) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
O2A1O1Ixp33_ASAP7_75t_L g171 ( .A1(n_142), .A2(n_157), .B(n_172), .C(n_173), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_SL g236 ( .A1(n_142), .A2(n_157), .B(n_237), .C(n_238), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_SL g482 ( .A1(n_142), .A2(n_157), .B(n_483), .C(n_484), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_SL g492 ( .A1(n_142), .A2(n_157), .B(n_493), .C(n_494), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_SL g514 ( .A1(n_142), .A2(n_157), .B(n_515), .C(n_516), .Y(n_514) );
O2A1O1Ixp33_ASAP7_75t_L g543 ( .A1(n_142), .A2(n_157), .B(n_544), .C(n_545), .Y(n_543) );
O2A1O1Ixp33_ASAP7_75t_SL g579 ( .A1(n_142), .A2(n_157), .B(n_580), .C(n_581), .Y(n_579) );
INVx5_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
BUFx3_ASAP7_75t_L g155 ( .A(n_144), .Y(n_155) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_144), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_151), .C(n_154), .Y(n_146) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_148), .A2(n_154), .B(n_203), .C(n_204), .Y(n_202) );
O2A1O1Ixp5_ASAP7_75t_L g505 ( .A1(n_148), .A2(n_506), .B(n_507), .C(n_508), .Y(n_505) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_148), .A2(n_508), .B(n_537), .C(n_538), .Y(n_536) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx4_ASAP7_75t_L g175 ( .A(n_150), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_152), .B(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g239 ( .A(n_152), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_L g525 ( .A1(n_152), .A2(n_216), .B(n_526), .C(n_527), .Y(n_525) );
OAI22xp33_ASAP7_75t_L g582 ( .A1(n_152), .A2(n_175), .B1(n_583), .B2(n_584), .Y(n_582) );
INVx5_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_153), .B(n_487), .Y(n_486) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g244 ( .A(n_155), .Y(n_244) );
INVx1_ASAP7_75t_L g497 ( .A(n_155), .Y(n_497) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_158), .A2(n_200), .B(n_201), .Y(n_199) );
INVx2_ASAP7_75t_L g218 ( .A(n_158), .Y(n_218) );
INVx1_ASAP7_75t_L g221 ( .A(n_158), .Y(n_221) );
OA21x2_ASAP7_75t_L g480 ( .A1(n_158), .A2(n_481), .B(n_488), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_L g522 ( .A1(n_158), .A2(n_252), .B(n_523), .C(n_524), .Y(n_522) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_159), .B(n_160), .Y(n_158) );
AND2x2_ASAP7_75t_L g169 ( .A(n_159), .B(n_160), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
AND2x2_ASAP7_75t_L g441 ( .A(n_164), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
OR2x2_ASAP7_75t_L g304 ( .A(n_165), .B(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_182), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_166), .B(n_285), .Y(n_284) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_166), .Y(n_297) );
INVx3_ASAP7_75t_L g312 ( .A(n_166), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_166), .B(n_182), .Y(n_336) );
OR2x2_ASAP7_75t_L g345 ( .A(n_166), .B(n_288), .Y(n_345) );
AND2x2_ASAP7_75t_L g349 ( .A(n_166), .B(n_309), .Y(n_349) );
AND2x2_ASAP7_75t_L g355 ( .A(n_166), .B(n_356), .Y(n_355) );
INVxp67_ASAP7_75t_L g392 ( .A(n_166), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_166), .B(n_249), .Y(n_406) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_170), .B(n_179), .Y(n_166) );
OA21x2_ASAP7_75t_L g490 ( .A1(n_167), .A2(n_491), .B(n_498), .Y(n_490) );
OA21x2_ASAP7_75t_L g512 ( .A1(n_167), .A2(n_513), .B(n_519), .Y(n_512) );
OA21x2_ASAP7_75t_L g541 ( .A1(n_167), .A2(n_542), .B(n_549), .Y(n_541) );
HB1xp67_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx4_ASAP7_75t_L g181 ( .A(n_168), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_168), .A2(n_185), .B(n_186), .Y(n_184) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g259 ( .A(n_169), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_174), .A2(n_227), .B(n_228), .C(n_229), .Y(n_226) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_175), .B(n_496), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_175), .B(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g216 ( .A(n_178), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_178), .B(n_582), .Y(n_581) );
OA21x2_ASAP7_75t_L g234 ( .A1(n_180), .A2(n_235), .B(n_245), .Y(n_234) );
INVx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_181), .B(n_206), .Y(n_205) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_181), .A2(n_224), .B(n_232), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_181), .B(n_233), .Y(n_232) );
AO21x2_ASAP7_75t_L g249 ( .A1(n_181), .A2(n_250), .B(n_257), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_181), .B(n_510), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_181), .B(n_529), .Y(n_528) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_181), .A2(n_533), .B(n_539), .Y(n_532) );
OR2x2_ASAP7_75t_L g298 ( .A(n_182), .B(n_249), .Y(n_298) );
AND2x2_ASAP7_75t_L g309 ( .A(n_182), .B(n_285), .Y(n_309) );
AND2x2_ASAP7_75t_L g321 ( .A(n_182), .B(n_312), .Y(n_321) );
NAND2xp5_ASAP7_75t_SL g344 ( .A(n_182), .B(n_249), .Y(n_344) );
INVx1_ASAP7_75t_SL g356 ( .A(n_182), .Y(n_356) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g248 ( .A(n_183), .B(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_183), .B(n_288), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_190), .B(n_191), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_191), .A2(n_255), .B(n_256), .Y(n_254) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx3_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_207), .Y(n_196) );
AND2x2_ASAP7_75t_L g269 ( .A(n_197), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_197), .B(n_222), .Y(n_273) );
AND2x2_ASAP7_75t_L g276 ( .A(n_197), .B(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_197), .B(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g301 ( .A(n_197), .B(n_292), .Y(n_301) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_197), .Y(n_320) );
AND2x2_ASAP7_75t_L g341 ( .A(n_197), .B(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g351 ( .A(n_197), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g397 ( .A(n_197), .B(n_280), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_197), .B(n_303), .Y(n_424) );
INVx5_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
BUFx2_ASAP7_75t_L g294 ( .A(n_198), .Y(n_294) );
AND2x2_ASAP7_75t_L g360 ( .A(n_198), .B(n_292), .Y(n_360) );
AND2x2_ASAP7_75t_L g444 ( .A(n_198), .B(n_312), .Y(n_444) );
OR2x6_ASAP7_75t_L g198 ( .A(n_199), .B(n_205), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_207), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g433 ( .A(n_207), .Y(n_433) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_222), .Y(n_207) );
AND2x2_ASAP7_75t_L g263 ( .A(n_208), .B(n_264), .Y(n_263) );
AND2x4_ASAP7_75t_L g272 ( .A(n_208), .B(n_270), .Y(n_272) );
INVx5_ASAP7_75t_L g280 ( .A(n_208), .Y(n_280) );
AND2x2_ASAP7_75t_L g303 ( .A(n_208), .B(n_234), .Y(n_303) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_208), .Y(n_340) );
OR2x6_ASAP7_75t_L g208 ( .A(n_209), .B(n_219), .Y(n_208) );
AOI21xp5_ASAP7_75t_SL g209 ( .A1(n_210), .A2(n_212), .B(n_217), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_216), .Y(n_213) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_218), .B(n_540), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_221), .A2(n_502), .B(n_509), .Y(n_501) );
INVx1_ASAP7_75t_L g381 ( .A(n_222), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_222), .B(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g414 ( .A(n_222), .B(n_280), .Y(n_414) );
A2O1A1Ixp33_ASAP7_75t_L g443 ( .A1(n_222), .A2(n_337), .B(n_444), .C(n_445), .Y(n_443) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_234), .Y(n_222) );
BUFx2_ASAP7_75t_L g264 ( .A(n_223), .Y(n_264) );
INVx2_ASAP7_75t_L g268 ( .A(n_223), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_231), .Y(n_224) );
HB1xp67_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx3_ASAP7_75t_L g548 ( .A(n_230), .Y(n_548) );
INVx2_ASAP7_75t_L g270 ( .A(n_234), .Y(n_270) );
AND2x2_ASAP7_75t_L g277 ( .A(n_234), .B(n_268), .Y(n_277) );
AND2x2_ASAP7_75t_L g368 ( .A(n_234), .B(n_280), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_242), .B(n_547), .Y(n_546) );
INVx4_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g485 ( .A(n_243), .Y(n_485) );
INVx2_ASAP7_75t_L g508 ( .A(n_244), .Y(n_508) );
AOI211x1_ASAP7_75t_SL g246 ( .A1(n_247), .A2(n_261), .B(n_274), .C(n_299), .Y(n_246) );
INVx1_ASAP7_75t_L g365 ( .A(n_247), .Y(n_365) );
AND2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_260), .Y(n_247) );
INVx5_ASAP7_75t_SL g285 ( .A(n_249), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_249), .B(n_355), .Y(n_354) );
AOI311xp33_ASAP7_75t_L g373 ( .A1(n_249), .A2(n_374), .A3(n_376), .B(n_377), .C(n_383), .Y(n_373) );
A2O1A1Ixp33_ASAP7_75t_L g408 ( .A1(n_249), .A2(n_321), .B(n_409), .C(n_412), .Y(n_408) );
OAI21xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_252), .B(n_253), .Y(n_250) );
OAI21xp5_ASAP7_75t_L g502 ( .A1(n_252), .A2(n_503), .B(n_504), .Y(n_502) );
OAI21xp5_ASAP7_75t_L g533 ( .A1(n_252), .A2(n_534), .B(n_535), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx2_ASAP7_75t_L g576 ( .A(n_259), .Y(n_576) );
INVxp67_ASAP7_75t_L g328 ( .A(n_260), .Y(n_328) );
NAND4xp25_ASAP7_75t_SL g261 ( .A(n_262), .B(n_265), .C(n_271), .D(n_273), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_262), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g319 ( .A(n_263), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_269), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_266), .B(n_272), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_266), .B(n_279), .Y(n_399) );
BUFx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_267), .B(n_280), .Y(n_417) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g292 ( .A(n_268), .Y(n_292) );
INVxp67_ASAP7_75t_L g327 ( .A(n_269), .Y(n_327) );
AND2x4_ASAP7_75t_L g279 ( .A(n_270), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g353 ( .A(n_270), .B(n_292), .Y(n_353) );
INVx1_ASAP7_75t_L g380 ( .A(n_270), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_270), .B(n_367), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_271), .B(n_341), .Y(n_361) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_272), .B(n_294), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_272), .B(n_341), .Y(n_440) );
INVx1_ASAP7_75t_L g451 ( .A(n_273), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_278), .B(n_281), .C(n_289), .Y(n_274) );
INVx1_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g293 ( .A(n_277), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g331 ( .A(n_277), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g313 ( .A(n_278), .Y(n_313) );
AND2x2_ASAP7_75t_L g290 ( .A(n_279), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_279), .B(n_341), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_279), .B(n_360), .Y(n_384) );
OR2x2_ASAP7_75t_L g300 ( .A(n_280), .B(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g332 ( .A(n_280), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_280), .B(n_292), .Y(n_347) );
AND2x2_ASAP7_75t_L g404 ( .A(n_280), .B(n_360), .Y(n_404) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_280), .Y(n_411) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AOI221xp5_ASAP7_75t_L g415 ( .A1(n_282), .A2(n_294), .B1(n_416), .B2(n_418), .C(n_421), .Y(n_415) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_286), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g305 ( .A(n_285), .B(n_288), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_285), .B(n_355), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_285), .B(n_312), .Y(n_420) );
INVx1_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g405 ( .A(n_287), .B(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g419 ( .A(n_287), .B(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_288), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g316 ( .A(n_288), .B(n_309), .Y(n_316) );
AND2x2_ASAP7_75t_L g386 ( .A(n_288), .B(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_288), .B(n_335), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_288), .B(n_436), .Y(n_435) );
OAI21xp5_ASAP7_75t_SL g289 ( .A1(n_290), .A2(n_293), .B(n_295), .Y(n_289) );
INVx2_ASAP7_75t_L g322 ( .A(n_290), .Y(n_322) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g342 ( .A(n_292), .Y(n_342) );
OR2x2_ASAP7_75t_L g346 ( .A(n_294), .B(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g449 ( .A(n_294), .B(n_417), .Y(n_449) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AOI21xp33_ASAP7_75t_SL g299 ( .A1(n_300), .A2(n_302), .B(n_304), .Y(n_299) );
INVx1_ASAP7_75t_L g453 ( .A(n_300), .Y(n_453) );
INVx2_ASAP7_75t_SL g367 ( .A(n_301), .Y(n_367) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_304), .A2(n_385), .B(n_449), .C(n_450), .Y(n_448) );
OAI322xp33_ASAP7_75t_SL g317 ( .A1(n_305), .A2(n_318), .A3(n_321), .B1(n_322), .B2(n_323), .C1(n_325), .C2(n_328), .Y(n_317) );
INVx2_ASAP7_75t_L g337 ( .A(n_305), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_313), .B1(n_314), .B2(n_316), .C(n_317), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OAI22xp33_ASAP7_75t_SL g383 ( .A1(n_308), .A2(n_384), .B1(n_385), .B2(n_388), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_309), .B(n_312), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_309), .B(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g382 ( .A(n_311), .B(n_344), .Y(n_382) );
INVx1_ASAP7_75t_L g372 ( .A(n_312), .Y(n_372) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g425 ( .A1(n_316), .A2(n_426), .B(n_428), .Y(n_425) );
AOI21xp33_ASAP7_75t_L g350 ( .A1(n_318), .A2(n_351), .B(n_354), .Y(n_350) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NOR2xp67_ASAP7_75t_SL g379 ( .A(n_320), .B(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_320), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g436 ( .A(n_321), .Y(n_436) );
INVx1_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND4xp25_ASAP7_75t_L g329 ( .A(n_330), .B(n_357), .C(n_373), .D(n_389), .Y(n_329) );
AOI211xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_333), .B(n_338), .C(n_350), .Y(n_330) );
INVx1_ASAP7_75t_L g422 ( .A(n_331), .Y(n_422) );
AND2x2_ASAP7_75t_L g370 ( .A(n_332), .B(n_353), .Y(n_370) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_337), .B(n_372), .Y(n_371) );
OAI22xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_343), .B1(n_346), .B2(n_348), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_340), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g388 ( .A(n_341), .Y(n_388) );
O2A1O1Ixp33_ASAP7_75t_L g402 ( .A1(n_341), .A2(n_380), .B(n_403), .C(n_405), .Y(n_402) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_L g387 ( .A(n_344), .Y(n_387) );
INVx1_ASAP7_75t_L g447 ( .A(n_345), .Y(n_447) );
NAND2xp33_ASAP7_75t_SL g437 ( .A(n_346), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g376 ( .A(n_355), .Y(n_376) );
O2A1O1Ixp33_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_361), .B(n_362), .C(n_364), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_366), .B1(n_369), .B2(n_371), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_367), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_372), .B(n_393), .Y(n_455) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AOI21xp33_ASAP7_75t_SL g377 ( .A1(n_378), .A2(n_381), .B(n_382), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_395), .B1(n_398), .B2(n_400), .C(n_402), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVxp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_405), .A2(n_422), .B1(n_423), .B2(n_424), .Y(n_421) );
NAND3xp33_ASAP7_75t_SL g407 ( .A(n_408), .B(n_415), .C(n_425), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
CKINVDCx16_ASAP7_75t_R g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVxp67_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OAI211xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_433), .B(n_434), .C(n_443), .Y(n_431) );
INVx1_ASAP7_75t_L g452 ( .A(n_432), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_437), .B1(n_439), .B2(n_441), .Y(n_434) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_452), .B1(n_453), .B2(n_454), .Y(n_450) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_L g464 ( .A(n_458), .Y(n_464) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g466 ( .A(n_464), .Y(n_466) );
NAND3xp33_ASAP7_75t_L g467 ( .A(n_465), .B(n_468), .C(n_760), .Y(n_467) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AOI22x1_ASAP7_75t_SL g757 ( .A1(n_471), .A2(n_742), .B1(n_758), .B2(n_759), .Y(n_757) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g758 ( .A(n_475), .Y(n_758) );
OR2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_672), .Y(n_475) );
NAND5xp2_ASAP7_75t_L g476 ( .A(n_477), .B(n_587), .C(n_619), .D(n_636), .E(n_659), .Y(n_476) );
AOI221xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_520), .B1(n_550), .B2(n_554), .C(n_558), .Y(n_477) );
INVx1_ASAP7_75t_L g699 ( .A(n_478), .Y(n_699) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_499), .Y(n_478) );
AND3x2_ASAP7_75t_L g674 ( .A(n_479), .B(n_501), .C(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_489), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_480), .B(n_556), .Y(n_555) );
BUFx3_ASAP7_75t_L g565 ( .A(n_480), .Y(n_565) );
AND2x2_ASAP7_75t_L g569 ( .A(n_480), .B(n_511), .Y(n_569) );
INVx2_ASAP7_75t_L g596 ( .A(n_480), .Y(n_596) );
OR2x2_ASAP7_75t_L g607 ( .A(n_480), .B(n_512), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_480), .B(n_500), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_480), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g686 ( .A(n_480), .B(n_512), .Y(n_686) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_489), .Y(n_568) );
AND2x2_ASAP7_75t_L g627 ( .A(n_489), .B(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_489), .B(n_500), .Y(n_646) );
INVx1_ASAP7_75t_SL g489 ( .A(n_490), .Y(n_489) );
OR2x2_ASAP7_75t_L g557 ( .A(n_490), .B(n_500), .Y(n_557) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_490), .Y(n_564) );
AND2x2_ASAP7_75t_L g613 ( .A(n_490), .B(n_512), .Y(n_613) );
NAND3xp33_ASAP7_75t_L g638 ( .A(n_490), .B(n_499), .C(n_596), .Y(n_638) );
AND2x2_ASAP7_75t_L g703 ( .A(n_490), .B(n_501), .Y(n_703) );
AND2x2_ASAP7_75t_L g737 ( .A(n_490), .B(n_500), .Y(n_737) );
INVxp67_ASAP7_75t_L g566 ( .A(n_499), .Y(n_566) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_511), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_500), .B(n_596), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_500), .B(n_627), .Y(n_635) );
AND2x2_ASAP7_75t_L g685 ( .A(n_500), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g713 ( .A(n_500), .Y(n_713) );
INVx4_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g620 ( .A(n_501), .B(n_613), .Y(n_620) );
BUFx3_ASAP7_75t_L g652 ( .A(n_501), .Y(n_652) );
INVx2_ASAP7_75t_L g628 ( .A(n_511), .Y(n_628) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_512), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_520), .A2(n_688), .B1(n_690), .B2(n_691), .Y(n_687) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_530), .Y(n_520) );
AND2x2_ASAP7_75t_L g550 ( .A(n_521), .B(n_551), .Y(n_550) );
INVx3_ASAP7_75t_SL g561 ( .A(n_521), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_521), .B(n_591), .Y(n_623) );
OR2x2_ASAP7_75t_L g642 ( .A(n_521), .B(n_531), .Y(n_642) );
AND2x2_ASAP7_75t_L g647 ( .A(n_521), .B(n_599), .Y(n_647) );
AND2x2_ASAP7_75t_L g650 ( .A(n_521), .B(n_592), .Y(n_650) );
AND2x2_ASAP7_75t_L g662 ( .A(n_521), .B(n_541), .Y(n_662) );
AND2x2_ASAP7_75t_L g678 ( .A(n_521), .B(n_532), .Y(n_678) );
AND2x4_ASAP7_75t_L g681 ( .A(n_521), .B(n_552), .Y(n_681) );
OR2x2_ASAP7_75t_L g698 ( .A(n_521), .B(n_634), .Y(n_698) );
OR2x2_ASAP7_75t_L g729 ( .A(n_521), .B(n_574), .Y(n_729) );
NAND2xp5_ASAP7_75t_SL g731 ( .A(n_521), .B(n_657), .Y(n_731) );
OR2x6_ASAP7_75t_L g521 ( .A(n_522), .B(n_528), .Y(n_521) );
AND2x2_ASAP7_75t_L g605 ( .A(n_530), .B(n_572), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_530), .B(n_592), .Y(n_724) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_541), .Y(n_530) );
AND2x2_ASAP7_75t_L g560 ( .A(n_531), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g591 ( .A(n_531), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g599 ( .A(n_531), .B(n_574), .Y(n_599) );
AND2x2_ASAP7_75t_L g617 ( .A(n_531), .B(n_552), .Y(n_617) );
OR2x2_ASAP7_75t_L g634 ( .A(n_531), .B(n_592), .Y(n_634) );
INVx2_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
BUFx2_ASAP7_75t_L g553 ( .A(n_532), .Y(n_553) );
AND2x2_ASAP7_75t_L g657 ( .A(n_532), .B(n_541), .Y(n_657) );
INVx2_ASAP7_75t_L g552 ( .A(n_541), .Y(n_552) );
INVx1_ASAP7_75t_L g669 ( .A(n_541), .Y(n_669) );
AND2x2_ASAP7_75t_L g719 ( .A(n_541), .B(n_561), .Y(n_719) );
AND2x2_ASAP7_75t_L g571 ( .A(n_551), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g603 ( .A(n_551), .B(n_561), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_551), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
AND2x2_ASAP7_75t_L g590 ( .A(n_552), .B(n_561), .Y(n_590) );
OR2x2_ASAP7_75t_L g706 ( .A(n_553), .B(n_680), .Y(n_706) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_556), .B(n_686), .Y(n_692) );
INVx2_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
OAI32xp33_ASAP7_75t_L g648 ( .A1(n_557), .A2(n_649), .A3(n_651), .B1(n_653), .B2(n_654), .Y(n_648) );
OR2x2_ASAP7_75t_L g665 ( .A(n_557), .B(n_607), .Y(n_665) );
OAI21xp33_ASAP7_75t_SL g690 ( .A1(n_557), .A2(n_567), .B(n_595), .Y(n_690) );
OAI22xp33_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_562), .B1(n_567), .B2(n_570), .Y(n_558) );
INVxp33_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_560), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_561), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g616 ( .A(n_561), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g716 ( .A(n_561), .B(n_657), .Y(n_716) );
OR2x2_ASAP7_75t_L g740 ( .A(n_561), .B(n_634), .Y(n_740) );
AOI21xp33_ASAP7_75t_L g723 ( .A1(n_562), .A2(n_622), .B(n_724), .Y(n_723) );
OR2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_566), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
INVx1_ASAP7_75t_L g600 ( .A(n_564), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_564), .B(n_569), .Y(n_618) );
AND2x2_ASAP7_75t_L g640 ( .A(n_565), .B(n_613), .Y(n_640) );
INVx1_ASAP7_75t_L g653 ( .A(n_565), .Y(n_653) );
OR2x2_ASAP7_75t_L g658 ( .A(n_565), .B(n_592), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_568), .B(n_607), .Y(n_606) );
OAI22xp33_ASAP7_75t_L g588 ( .A1(n_569), .A2(n_589), .B1(n_594), .B2(n_598), .Y(n_588) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_572), .A2(n_631), .B1(n_638), .B2(n_639), .Y(n_637) );
AND2x2_ASAP7_75t_L g715 ( .A(n_572), .B(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_574), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g734 ( .A(n_574), .B(n_617), .Y(n_734) );
AO21x2_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_577), .B(n_585), .Y(n_574) );
INVx1_ASAP7_75t_L g593 ( .A(n_575), .Y(n_593) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OA21x2_ASAP7_75t_L g592 ( .A1(n_578), .A2(n_586), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AOI221xp5_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_600), .B1(n_601), .B2(n_606), .C(n_608), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_590), .B(n_592), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_590), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g609 ( .A(n_591), .Y(n_609) );
O2A1O1Ixp33_ASAP7_75t_L g696 ( .A1(n_591), .A2(n_697), .B(n_698), .C(n_699), .Y(n_696) );
AND2x2_ASAP7_75t_L g701 ( .A(n_591), .B(n_681), .Y(n_701) );
O2A1O1Ixp33_ASAP7_75t_SL g739 ( .A1(n_591), .A2(n_680), .B(n_740), .C(n_741), .Y(n_739) );
BUFx3_ASAP7_75t_L g631 ( .A(n_592), .Y(n_631) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_595), .B(n_652), .Y(n_695) );
AOI211xp5_ASAP7_75t_L g714 ( .A1(n_595), .A2(n_715), .B(n_717), .C(n_723), .Y(n_714) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
INVxp67_ASAP7_75t_L g675 ( .A(n_597), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_599), .B(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_602), .B(n_604), .Y(n_601) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
AOI211xp5_ASAP7_75t_L g619 ( .A1(n_603), .A2(n_620), .B(n_621), .C(n_629), .Y(n_619) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g704 ( .A(n_607), .Y(n_704) );
OR2x2_ASAP7_75t_L g721 ( .A(n_607), .B(n_651), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B1(n_615), .B2(n_618), .Y(n_608) );
OAI22xp33_ASAP7_75t_L g621 ( .A1(n_610), .A2(n_622), .B1(n_623), .B2(n_624), .Y(n_621) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
OR2x2_ASAP7_75t_L g708 ( .A(n_612), .B(n_652), .Y(n_708) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g663 ( .A(n_613), .B(n_653), .Y(n_663) );
INVx1_ASAP7_75t_L g671 ( .A(n_614), .Y(n_671) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_617), .B(n_631), .Y(n_679) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_627), .B(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g736 ( .A(n_628), .Y(n_736) );
AOI21xp33_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_632), .B(n_635), .Y(n_629) );
INVx1_ASAP7_75t_L g666 ( .A(n_630), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_631), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_631), .B(n_662), .Y(n_661) );
NAND2x1p5_ASAP7_75t_L g682 ( .A(n_631), .B(n_657), .Y(n_682) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_631), .B(n_678), .Y(n_689) );
OAI211xp5_ASAP7_75t_L g693 ( .A1(n_631), .A2(n_641), .B(n_681), .C(n_694), .Y(n_693) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
AOI221xp5_ASAP7_75t_SL g636 ( .A1(n_637), .A2(n_641), .B1(n_643), .B2(n_647), .C(n_648), .Y(n_636) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVxp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_645), .B(n_653), .Y(n_727) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
O2A1O1Ixp33_ASAP7_75t_L g738 ( .A1(n_647), .A2(n_662), .B(n_664), .C(n_739), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_650), .B(n_657), .Y(n_722) );
NAND2xp5_ASAP7_75t_SL g741 ( .A(n_651), .B(n_704), .Y(n_741) );
CKINVDCx16_ASAP7_75t_R g651 ( .A(n_652), .Y(n_651) );
INVxp33_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_656), .B(n_658), .Y(n_655) );
AOI21xp33_ASAP7_75t_SL g667 ( .A1(n_656), .A2(n_668), .B(n_670), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_656), .B(n_729), .Y(n_728) );
INVx2_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_657), .B(n_711), .Y(n_710) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_663), .B1(n_664), .B2(n_666), .C(n_667), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_663), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g697 ( .A(n_669), .Y(n_697) );
NAND5xp2_ASAP7_75t_L g672 ( .A(n_673), .B(n_700), .C(n_714), .D(n_725), .E(n_738), .Y(n_672) );
AOI211xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_676), .B(n_683), .C(n_696), .Y(n_673) );
INVx2_ASAP7_75t_SL g720 ( .A(n_674), .Y(n_720) );
NAND4xp25_ASAP7_75t_SL g676 ( .A(n_677), .B(n_679), .C(n_680), .D(n_682), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx3_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OAI211xp5_ASAP7_75t_SL g683 ( .A1(n_682), .A2(n_684), .B(n_687), .C(n_693), .Y(n_683) );
CKINVDCx20_ASAP7_75t_R g684 ( .A(n_685), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g725 ( .A1(n_685), .A2(n_726), .B1(n_728), .B2(n_730), .C(n_732), .Y(n_725) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AOI221xp5_ASAP7_75t_SL g700 ( .A1(n_701), .A2(n_702), .B1(n_705), .B2(n_707), .C(n_709), .Y(n_700) );
AND2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_708), .A2(n_731), .B1(n_733), .B2(n_735), .Y(n_732) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_720), .B1(n_721), .B2(n_722), .Y(n_717) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_746), .Y(n_755) );
CKINVDCx16_ASAP7_75t_R g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
endmodule