module fake_jpeg_31304_n_372 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_372);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_372;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_32),
.B(n_17),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_51),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

CKINVDCx6p67_ASAP7_75t_R g117 ( 
.A(n_47),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_14),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_32),
.B(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_28),
.Y(n_77)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_15),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_63),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_20),
.B(n_0),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_34),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_64),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_71),
.Y(n_85)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_18),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_73),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_81),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_21),
.C(n_42),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_80),
.B(n_92),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_38),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_43),
.B1(n_42),
.B2(n_34),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_82),
.A2(n_88),
.B1(n_106),
.B2(n_113),
.Y(n_142)
);

NAND2xp33_ASAP7_75t_SL g84 ( 
.A(n_59),
.B(n_43),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_84),
.Y(n_154)
);

NAND2xp33_ASAP7_75t_SL g86 ( 
.A(n_56),
.B(n_43),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g145 ( 
.A1(n_86),
.A2(n_69),
.B1(n_52),
.B2(n_39),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_64),
.A2(n_43),
.B1(n_42),
.B2(n_21),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_L g89 ( 
.A1(n_58),
.A2(n_41),
.B(n_29),
.Y(n_89)
);

OAI32xp33_ASAP7_75t_L g134 ( 
.A1(n_89),
.A2(n_70),
.A3(n_47),
.B1(n_39),
.B2(n_18),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_21),
.B1(n_31),
.B2(n_29),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_90),
.A2(n_96),
.B1(n_110),
.B2(n_120),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_63),
.A2(n_41),
.B(n_29),
.C(n_27),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_20),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_119),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_54),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_94),
.A2(n_61),
.B1(n_50),
.B2(n_53),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_45),
.A2(n_33),
.B1(n_38),
.B2(n_20),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_46),
.B(n_38),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_98),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_55),
.B(n_41),
.C(n_27),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_101),
.B(n_30),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_33),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_103),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_56),
.A2(n_40),
.B1(n_22),
.B2(n_36),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_47),
.B(n_36),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_108),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_45),
.A2(n_36),
.B1(n_28),
.B2(n_24),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_52),
.A2(n_40),
.B1(n_22),
.B2(n_28),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_48),
.B(n_39),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_73),
.A2(n_24),
.B1(n_22),
.B2(n_40),
.Y(n_120)
);

BUFx2_ASAP7_75t_SL g122 ( 
.A(n_117),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_123),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_94),
.A2(n_73),
.B1(n_72),
.B2(n_71),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_126),
.A2(n_137),
.B1(n_144),
.B2(n_146),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_127),
.B(n_85),
.C(n_114),
.Y(n_171)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_128),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_90),
.A2(n_61),
.B1(n_71),
.B2(n_48),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_129),
.A2(n_138),
.B1(n_139),
.B2(n_100),
.Y(n_195)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_132),
.Y(n_165)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_77),
.B(n_72),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_133),
.B(n_140),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_134),
.B(n_117),
.Y(n_172)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_135),
.B(n_145),
.Y(n_187)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_136),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_89),
.A2(n_50),
.B1(n_53),
.B2(n_57),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_84),
.A2(n_57),
.B1(n_62),
.B2(n_65),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_65),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_95),
.A2(n_62),
.B1(n_24),
.B2(n_70),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_74),
.A2(n_70),
.B1(n_47),
.B2(n_69),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_101),
.B(n_39),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_147),
.B(n_39),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_117),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_159),
.Y(n_169)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_87),
.Y(n_150)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_153),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g155 ( 
.A1(n_86),
.A2(n_39),
.B1(n_66),
.B2(n_44),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_155),
.A2(n_83),
.B1(n_109),
.B2(n_118),
.Y(n_180)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_87),
.Y(n_156)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_111),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_157),
.B(n_158),
.Y(n_192)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_111),
.Y(n_158)
);

OAI32xp33_ASAP7_75t_L g159 ( 
.A1(n_76),
.A2(n_68),
.A3(n_39),
.B1(n_15),
.B2(n_14),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_97),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_74),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_161),
.Y(n_164)
);

NOR3xp33_ASAP7_75t_SL g163 ( 
.A(n_121),
.B(n_79),
.C(n_125),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_163),
.B(n_167),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_154),
.A2(n_85),
.B1(n_92),
.B2(n_114),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_166),
.B(n_145),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_157),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_131),
.A2(n_119),
.B1(n_80),
.B2(n_114),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_168),
.A2(n_172),
.B1(n_177),
.B2(n_180),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_178),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_158),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_173),
.B(n_179),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

BUFx8_ASAP7_75t_L g216 ( 
.A(n_176),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_131),
.A2(n_83),
.B1(n_109),
.B2(n_85),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_124),
.B(n_79),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_125),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_184),
.B(n_190),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_124),
.B(n_97),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_185),
.B(n_196),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_133),
.A2(n_142),
.B1(n_137),
.B2(n_140),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_188),
.A2(n_191),
.B1(n_141),
.B2(n_129),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_127),
.B(n_102),
.C(n_99),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_134),
.A2(n_107),
.B1(n_104),
.B2(n_118),
.Y(n_191)
);

BUFx24_ASAP7_75t_SL g193 ( 
.A(n_149),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_121),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_195),
.A2(n_197),
.B1(n_148),
.B2(n_143),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_102),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_143),
.A2(n_104),
.B1(n_107),
.B2(n_116),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_199),
.B(n_213),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_201),
.A2(n_224),
.B1(n_165),
.B2(n_174),
.Y(n_240)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_175),
.Y(n_202)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_204),
.A2(n_205),
.B1(n_231),
.B2(n_233),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_188),
.A2(n_191),
.B1(n_187),
.B2(n_169),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_175),
.Y(n_208)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_208),
.Y(n_237)
);

AOI32xp33_ASAP7_75t_L g209 ( 
.A1(n_178),
.A2(n_184),
.A3(n_172),
.B1(n_163),
.B2(n_187),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_209),
.A2(n_212),
.B(n_228),
.Y(n_243)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_198),
.Y(n_210)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_210),
.Y(n_241)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_189),
.Y(n_211)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_211),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_128),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_218),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_194),
.B(n_149),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_215),
.B(n_219),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_192),
.Y(n_217)
);

NAND3xp33_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_222),
.C(n_223),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_168),
.B(n_123),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_220),
.B(n_183),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_167),
.B(n_152),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_221),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_173),
.B(n_141),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_183),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_195),
.A2(n_159),
.B1(n_145),
.B2(n_155),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_171),
.B(n_132),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_165),
.C(n_162),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_198),
.B(n_130),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_226),
.B(n_227),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_135),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_166),
.A2(n_145),
.B(n_155),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_183),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_230),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_177),
.A2(n_180),
.B1(n_170),
.B2(n_197),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_189),
.Y(n_232)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_232),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_170),
.A2(n_155),
.B1(n_116),
.B2(n_150),
.Y(n_233)
);

AOI221xp5_ASAP7_75t_L g234 ( 
.A1(n_209),
.A2(n_213),
.B1(n_220),
.B2(n_203),
.C(n_228),
.Y(n_234)
);

AOI221xp5_ASAP7_75t_L g281 ( 
.A1(n_234),
.A2(n_18),
.B1(n_1),
.B2(n_2),
.C(n_3),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_212),
.A2(n_165),
.B(n_174),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_236),
.A2(n_246),
.B(n_249),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_240),
.A2(n_262),
.B1(n_233),
.B2(n_230),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_260),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_212),
.A2(n_205),
.B(n_218),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_200),
.A2(n_181),
.B(n_162),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_217),
.A2(n_181),
.B1(n_182),
.B2(n_99),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_250),
.A2(n_255),
.B(n_0),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_206),
.A2(n_182),
.B(n_136),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_252),
.A2(n_232),
.B(n_112),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_204),
.A2(n_161),
.B1(n_100),
.B2(n_156),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_253),
.A2(n_75),
.B1(n_216),
.B2(n_30),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_261),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_200),
.A2(n_151),
.B(n_186),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_202),
.Y(n_258)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_258),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_215),
.B(n_12),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_259),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_214),
.B(n_186),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_231),
.A2(n_176),
.B1(n_164),
.B2(n_112),
.Y(n_262)
);

NAND3xp33_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_210),
.C(n_208),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_263),
.B(n_276),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_238),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_271),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_266),
.A2(n_278),
.B1(n_253),
.B2(n_248),
.Y(n_287)
);

OAI322xp33_ASAP7_75t_L g267 ( 
.A1(n_242),
.A2(n_207),
.A3(n_229),
.B1(n_225),
.B2(n_223),
.C1(n_216),
.C2(n_153),
.Y(n_267)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_267),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_260),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_268),
.B(n_272),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_229),
.Y(n_269)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_235),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_211),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_279),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_273),
.B(n_282),
.Y(n_294)
);

AOI322xp5_ASAP7_75t_L g274 ( 
.A1(n_243),
.A2(n_207),
.A3(n_153),
.B1(n_216),
.B2(n_75),
.C1(n_164),
.C2(n_12),
.Y(n_274)
);

AOI322xp5_ASAP7_75t_L g288 ( 
.A1(n_274),
.A2(n_281),
.A3(n_282),
.B1(n_265),
.B2(n_276),
.C1(n_273),
.C2(n_252),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_275),
.A2(n_283),
.B1(n_250),
.B2(n_245),
.Y(n_293)
);

A2O1A1O1Ixp25_ASAP7_75t_L g276 ( 
.A1(n_246),
.A2(n_216),
.B(n_15),
.C(n_13),
.D(n_18),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_240),
.A2(n_75),
.B1(n_30),
.B2(n_18),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_242),
.B(n_0),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_235),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_280),
.B(n_284),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_243),
.A2(n_18),
.B(n_1),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_246),
.A2(n_3),
.B(n_4),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_287),
.A2(n_288),
.B1(n_301),
.B2(n_302),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_244),
.C(n_249),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_292),
.C(n_295),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_244),
.C(n_249),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_293),
.B(n_296),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_234),
.C(n_236),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_285),
.B(n_259),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_258),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_266),
.A2(n_248),
.B1(n_255),
.B2(n_245),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_278),
.A2(n_255),
.B1(n_236),
.B2(n_250),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_267),
.B(n_261),
.C(n_257),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_304),
.C(n_306),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_257),
.C(n_247),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_247),
.C(n_262),
.Y(n_306)
);

NOR3xp33_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_291),
.C(n_295),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g334 ( 
.A(n_307),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_296),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_301),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_277),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_309),
.B(n_322),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_299),
.B(n_277),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_310),
.A2(n_318),
.B1(n_287),
.B2(n_256),
.Y(n_326)
);

OAI322xp33_ASAP7_75t_L g313 ( 
.A1(n_300),
.A2(n_279),
.A3(n_268),
.B1(n_284),
.B2(n_276),
.C1(n_274),
.C2(n_283),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_313),
.B(n_319),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_294),
.A2(n_271),
.B(n_264),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_315),
.A2(n_320),
.B(n_312),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_292),
.B(n_280),
.C(n_264),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_323),
.C(n_251),
.Y(n_330)
);

NOR3xp33_ASAP7_75t_SL g319 ( 
.A(n_305),
.B(n_241),
.C(n_237),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_302),
.A2(n_275),
.B(n_241),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_298),
.B(n_304),
.Y(n_321)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_321),
.Y(n_327)
);

XNOR2x1_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_237),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_303),
.B(n_256),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_324),
.B(n_325),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_326),
.B(n_329),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_310),
.A2(n_251),
.B1(n_4),
.B2(n_6),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_330),
.B(n_314),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_312),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_331),
.B(n_337),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_311),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_315),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_317),
.B(n_7),
.C(n_8),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_316),
.C(n_323),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_308),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_335),
.A2(n_320),
.B1(n_311),
.B2(n_319),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_321),
.B(n_9),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_338),
.B(n_339),
.Y(n_351)
);

OAI221xp5_ASAP7_75t_L g340 ( 
.A1(n_334),
.A2(n_313),
.B1(n_309),
.B2(n_314),
.C(n_316),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_340),
.A2(n_11),
.B(n_342),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_341),
.B(n_342),
.Y(n_355)
);

NAND4xp25_ASAP7_75t_L g345 ( 
.A(n_336),
.B(n_322),
.C(n_10),
.D(n_11),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_345),
.B(n_347),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_327),
.B(n_9),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_328),
.B(n_10),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_348),
.B(n_332),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_343),
.A2(n_324),
.B(n_327),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_349),
.B(n_350),
.Y(n_358)
);

NOR2x1_ASAP7_75t_L g350 ( 
.A(n_338),
.B(n_335),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_353),
.B(n_348),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_344),
.A2(n_330),
.B(n_333),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_354),
.B(n_356),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_341),
.A2(n_11),
.B1(n_328),
.B2(n_339),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_357),
.B(n_346),
.Y(n_361)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_352),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_359),
.B(n_360),
.Y(n_365)
);

AOI21x1_ASAP7_75t_L g366 ( 
.A1(n_361),
.A2(n_364),
.B(n_358),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_351),
.B(n_11),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_363),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_349),
.B(n_350),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_366),
.B(n_368),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_362),
.B(n_355),
.C(n_354),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_365),
.B(n_355),
.C(n_359),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_369),
.A2(n_367),
.B(n_356),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_371),
.B(n_370),
.Y(n_372)
);


endmodule