module fake_jpeg_4255_n_257 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_152;
wire n_182;
wire n_19;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_SL g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_40),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_1),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g39 ( 
.A1(n_20),
.A2(n_2),
.B(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_19),
.B1(n_21),
.B2(n_16),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_42),
.A2(n_44),
.B1(n_46),
.B2(n_50),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_19),
.B1(n_21),
.B2(n_16),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_48),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_21),
.B1(n_16),
.B2(n_30),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_16),
.Y(n_49)
);

OAI21xp33_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_22),
.B(n_29),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_17),
.B1(n_25),
.B2(n_24),
.Y(n_50)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_17),
.B1(n_25),
.B2(n_24),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_58),
.Y(n_94)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_59),
.B(n_60),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_55),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_62),
.B(n_65),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_20),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_74),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_23),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_SL g66 ( 
.A1(n_49),
.A2(n_40),
.B(n_28),
.C(n_27),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_66),
.A2(n_26),
.B1(n_35),
.B2(n_5),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_67),
.Y(n_110)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_42),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_47),
.B(n_23),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_32),
.B(n_31),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_20),
.B(n_15),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_44),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_45),
.B(n_29),
.Y(n_75)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_52),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_80),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_54),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_85),
.B1(n_87),
.B2(n_28),
.Y(n_92)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_54),
.B(n_32),
.Y(n_83)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_41),
.B(n_31),
.Y(n_84)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_53),
.A2(n_28),
.B1(n_27),
.B2(n_26),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_53),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_3),
.Y(n_112)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_88),
.A2(n_96),
.B1(n_104),
.B2(n_66),
.Y(n_122)
);

AND2x6_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_35),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_89),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_92),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_64),
.A2(n_60),
.B1(n_58),
.B2(n_74),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_27),
.B1(n_26),
.B2(n_20),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_98),
.B(n_81),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_35),
.C(n_15),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_82),
.C(n_79),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_64),
.A2(n_14),
.B1(n_4),
.B2(n_5),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_105),
.Y(n_128)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_116),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_119),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_118),
.B(n_120),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_97),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_123),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_122),
.A2(n_126),
.B1(n_134),
.B2(n_140),
.Y(n_156)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_108),
.B(n_69),
.Y(n_124)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_137),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_66),
.B1(n_62),
.B2(n_65),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_90),
.A2(n_65),
.B(n_66),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_127),
.A2(n_118),
.B(n_120),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_128),
.B(n_132),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_80),
.Y(n_129)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_59),
.Y(n_130)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_68),
.Y(n_131)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_113),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_94),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_135),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_90),
.A2(n_66),
.B1(n_56),
.B2(n_61),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_108),
.B(n_57),
.Y(n_136)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_110),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_114),
.A2(n_91),
.B(n_89),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_144),
.A2(n_149),
.B(n_152),
.Y(n_173)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_146),
.B(n_151),
.Y(n_176)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_114),
.A2(n_110),
.B(n_88),
.Y(n_152)
);

BUFx4f_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

INVx13_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_139),
.A2(n_107),
.B(n_104),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_154),
.A2(n_157),
.B1(n_166),
.B2(n_167),
.Y(n_185)
);

XNOR2x1_ASAP7_75t_SL g182 ( 
.A(n_155),
.B(n_102),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_135),
.A2(n_96),
.B1(n_99),
.B2(n_103),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_158),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_117),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_160),
.B(n_106),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_119),
.A2(n_99),
.B(n_103),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_133),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_138),
.A2(n_100),
.B1(n_77),
.B2(n_87),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_121),
.A2(n_105),
.B(n_112),
.Y(n_167)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

A2O1A1O1Ixp25_ASAP7_75t_L g170 ( 
.A1(n_144),
.A2(n_127),
.B(n_152),
.C(n_162),
.D(n_125),
.Y(n_170)
);

OAI322xp33_ASAP7_75t_L g199 ( 
.A1(n_170),
.A2(n_182),
.A3(n_156),
.B1(n_142),
.B2(n_159),
.C1(n_161),
.C2(n_164),
.Y(n_199)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_177),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_123),
.Y(n_172)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_140),
.Y(n_174)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_105),
.Y(n_175)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_132),
.Y(n_178)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_151),
.A2(n_112),
.B1(n_93),
.B2(n_115),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_188),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_102),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_187),
.Y(n_201)
);

HB1xp67_ASAP7_75t_SL g183 ( 
.A(n_154),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_183),
.A2(n_186),
.B1(n_73),
.B2(n_153),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_184),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_146),
.A2(n_73),
.B1(n_78),
.B2(n_106),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_167),
.B(n_150),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_162),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_200),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_178),
.A2(n_156),
.B1(n_149),
.B2(n_166),
.Y(n_197)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

OAI322xp33_ASAP7_75t_L g216 ( 
.A1(n_199),
.A2(n_179),
.A3(n_14),
.B1(n_169),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_173),
.B(n_163),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_160),
.Y(n_202)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_202),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_203),
.A2(n_191),
.B1(n_171),
.B2(n_198),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_180),
.A2(n_182),
.B1(n_168),
.B2(n_176),
.Y(n_204)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_204),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_185),
.A2(n_153),
.B1(n_6),
.B2(n_7),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_205),
.Y(n_210)
);

OAI21x1_ASAP7_75t_L g206 ( 
.A1(n_197),
.A2(n_185),
.B(n_187),
.Y(n_206)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_170),
.C(n_174),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_201),
.C(n_190),
.Y(n_226)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_211),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_198),
.A2(n_188),
.B1(n_177),
.B2(n_186),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_213),
.A2(n_218),
.B1(n_189),
.B2(n_195),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_175),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_217),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_216),
.B(n_4),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_169),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_192),
.A2(n_181),
.B(n_6),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_181),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_204),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_223),
.B(n_226),
.C(n_228),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_229),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_213),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_227),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_208),
.A2(n_190),
.B1(n_201),
.B2(n_196),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_196),
.C(n_193),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_7),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_230),
.B(n_207),
.C(n_219),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_220),
.A2(n_208),
.B1(n_211),
.B2(n_212),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_234),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_237),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_222),
.A2(n_210),
.B1(n_226),
.B2(n_221),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_227),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_235),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_217),
.Y(n_237)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_240),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_209),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_241),
.A2(n_242),
.B(n_243),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_218),
.Y(n_242)
);

AOI21x1_ASAP7_75t_L g243 ( 
.A1(n_233),
.A2(n_223),
.B(n_224),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_214),
.Y(n_245)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_245),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_232),
.C(n_230),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_247),
.A2(n_249),
.B(n_13),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_7),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_251),
.A2(n_248),
.B(n_246),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_249),
.B(n_8),
.Y(n_252)
);

AOI322xp5_ASAP7_75t_L g254 ( 
.A1(n_252),
.A2(n_9),
.A3(n_10),
.B1(n_12),
.B2(n_13),
.C1(n_251),
.C2(n_229),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_253),
.B(n_254),
.C(n_250),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_9),
.Y(n_256)
);

BUFx24_ASAP7_75t_SL g257 ( 
.A(n_256),
.Y(n_257)
);


endmodule